magic
tech sky130A
magscale 1 2
timestamp 1640987651
<< xpolycontact >>
rect -2520 4130 -2380 4610
rect -2520 -6950 -2380 -6470
rect -2130 4130 -1990 4610
rect -2130 -6950 -1990 -6470
rect -1740 4130 -1600 4610
rect 16380 4130 16520 4610
rect -330 -380 150 -98
rect 7150 -380 7630 -98
rect 14630 -380 15110 -98
rect -1350 -4552 -870 -4270
rect -588 -4552 -110 -4270
rect 14890 -4552 15368 -4270
rect 15650 -4552 16130 -4270
rect -1740 -6950 -1600 -6470
rect 16380 -6950 16520 -6470
rect 16770 4130 16910 4610
rect 16770 -6950 16910 -6470
rect 17160 4130 17300 4610
rect 17160 -6950 17300 -6470
rect -270 -9900 210 -9618
rect 7210 -9900 7690 -9618
rect 14690 -9900 15170 -9618
<< xpolyres >>
rect -2520 -6470 -2380 4130
rect -2130 -6470 -1990 4130
rect -1740 -6470 -1600 4130
rect 150 -380 7150 -98
rect 7630 -380 14630 -98
rect -870 -4552 -588 -4270
rect 15368 -4552 15650 -4270
rect 16380 -6470 16520 4130
rect 16770 -6470 16910 4130
rect 17160 -6470 17300 4130
rect 210 -9900 7210 -9618
rect 7690 -9900 14690 -9618
<< viali >>
rect -2480 4550 -2420 4590
rect -2480 4470 -2420 4510
rect -2480 4390 -2420 4430
rect -2480 4310 -2420 4350
rect -2480 4230 -2420 4270
rect -2480 4150 -2420 4190
rect -2090 4550 -2030 4590
rect -2090 4470 -2030 4510
rect -2090 4390 -2030 4430
rect -2090 4310 -2030 4350
rect -2090 4230 -2030 4270
rect -2090 4150 -2030 4190
rect -1700 4550 -1640 4590
rect -1700 4470 -1640 4510
rect -1700 4390 -1640 4430
rect -1700 4310 -1640 4350
rect -1700 4230 -1640 4270
rect -1700 4150 -1640 4190
rect 16420 4550 16480 4590
rect 16420 4470 16480 4510
rect 16420 4390 16480 4430
rect 16420 4310 16480 4350
rect 16420 4230 16480 4270
rect 16420 4150 16480 4190
rect 16810 4550 16870 4590
rect 16810 4470 16870 4510
rect 16810 4390 16870 4430
rect 16810 4310 16870 4350
rect 16810 4230 16870 4270
rect 16810 4150 16870 4190
rect 17200 4550 17260 4590
rect 17200 4470 17260 4510
rect 17200 4390 17260 4430
rect 17200 4310 17260 4350
rect 17200 4230 17260 4270
rect 17200 4150 17260 4190
rect -310 -180 -270 -140
rect -230 -180 -190 -140
rect -150 -180 -110 -140
rect -70 -180 -30 -140
rect 10 -180 50 -140
rect 90 -180 130 -140
rect -310 -260 -270 -220
rect -230 -260 -190 -220
rect -150 -260 -110 -220
rect -70 -260 -30 -220
rect 10 -260 50 -220
rect 90 -260 130 -220
rect -310 -340 -270 -300
rect -230 -340 -190 -300
rect -150 -340 -110 -300
rect -70 -340 -30 -300
rect 10 -340 50 -300
rect 90 -340 130 -300
rect 7170 -180 7210 -140
rect 7250 -180 7290 -140
rect 7330 -180 7370 -140
rect 7410 -180 7450 -140
rect 7490 -180 7530 -140
rect 7570 -180 7610 -140
rect 7170 -260 7210 -220
rect 7250 -260 7290 -220
rect 7330 -260 7370 -220
rect 7410 -260 7450 -220
rect 7490 -260 7530 -220
rect 7570 -260 7610 -220
rect 7170 -340 7210 -300
rect 7250 -340 7290 -300
rect 7330 -340 7370 -300
rect 7410 -340 7450 -300
rect 7490 -340 7530 -300
rect 7570 -340 7610 -300
rect 14650 -180 14690 -140
rect 14730 -180 14770 -140
rect 14810 -180 14850 -140
rect 14890 -180 14930 -140
rect 14970 -180 15010 -140
rect 15050 -180 15090 -140
rect 14650 -260 14690 -220
rect 14730 -260 14770 -220
rect 14810 -260 14850 -220
rect 14890 -260 14930 -220
rect 14970 -260 15010 -220
rect 15050 -260 15090 -220
rect 14650 -340 14690 -300
rect 14730 -340 14770 -300
rect 14810 -340 14850 -300
rect 14890 -340 14930 -300
rect 14970 -340 15010 -300
rect 15050 -340 15090 -300
rect -1330 -4352 -1290 -4312
rect -1250 -4352 -1210 -4312
rect -1170 -4352 -1130 -4312
rect -1090 -4352 -1050 -4312
rect -1010 -4352 -970 -4312
rect -930 -4352 -890 -4312
rect -1330 -4432 -1290 -4392
rect -1250 -4432 -1210 -4392
rect -1170 -4432 -1130 -4392
rect -1090 -4432 -1050 -4392
rect -1010 -4432 -970 -4392
rect -930 -4432 -890 -4392
rect -1330 -4512 -1290 -4472
rect -1250 -4512 -1210 -4472
rect -1170 -4512 -1130 -4472
rect -1090 -4512 -1050 -4472
rect -1010 -4512 -970 -4472
rect -930 -4512 -890 -4472
rect -570 -4352 -530 -4312
rect -490 -4352 -450 -4312
rect -410 -4352 -370 -4312
rect -330 -4352 -290 -4312
rect -250 -4352 -210 -4312
rect -170 -4352 -130 -4312
rect -570 -4432 -530 -4392
rect -490 -4432 -450 -4392
rect -410 -4432 -370 -4392
rect -330 -4432 -290 -4392
rect -250 -4432 -210 -4392
rect -170 -4432 -130 -4392
rect -570 -4512 -530 -4472
rect -490 -4512 -450 -4472
rect -410 -4512 -370 -4472
rect -330 -4512 -290 -4472
rect -250 -4512 -210 -4472
rect -170 -4512 -130 -4472
rect 14910 -4352 14950 -4312
rect 14990 -4352 15030 -4312
rect 15070 -4352 15110 -4312
rect 15150 -4352 15190 -4312
rect 15230 -4352 15270 -4312
rect 15310 -4352 15350 -4312
rect 14910 -4432 14950 -4392
rect 14990 -4432 15030 -4392
rect 15070 -4432 15110 -4392
rect 15150 -4432 15190 -4392
rect 15230 -4432 15270 -4392
rect 15310 -4432 15350 -4392
rect 14910 -4512 14950 -4472
rect 14990 -4512 15030 -4472
rect 15070 -4512 15110 -4472
rect 15150 -4512 15190 -4472
rect 15230 -4512 15270 -4472
rect 15310 -4512 15350 -4472
rect 15670 -4352 15710 -4312
rect 15750 -4352 15790 -4312
rect 15830 -4352 15870 -4312
rect 15910 -4352 15950 -4312
rect 15990 -4352 16030 -4312
rect 16070 -4352 16110 -4312
rect 15670 -4432 15710 -4392
rect 15750 -4432 15790 -4392
rect 15830 -4432 15870 -4392
rect 15910 -4432 15950 -4392
rect 15990 -4432 16030 -4392
rect 16070 -4432 16110 -4392
rect 15670 -4512 15710 -4472
rect 15750 -4512 15790 -4472
rect 15830 -4512 15870 -4472
rect 15910 -4512 15950 -4472
rect 15990 -4512 16030 -4472
rect 16070 -4512 16110 -4472
rect -2480 -6530 -2420 -6490
rect -2480 -6610 -2420 -6570
rect -2480 -6690 -2420 -6650
rect -2480 -6770 -2420 -6730
rect -2480 -6850 -2420 -6810
rect -2480 -6930 -2420 -6890
rect -2090 -6530 -2030 -6490
rect -2090 -6610 -2030 -6570
rect -2090 -6690 -2030 -6650
rect -2090 -6770 -2030 -6730
rect -2090 -6850 -2030 -6810
rect -2090 -6930 -2030 -6890
rect -1700 -6530 -1640 -6490
rect -1700 -6610 -1640 -6570
rect -1700 -6690 -1640 -6650
rect -1700 -6770 -1640 -6730
rect -1700 -6850 -1640 -6810
rect -1700 -6930 -1640 -6890
rect 16420 -6530 16480 -6490
rect 16420 -6610 16480 -6570
rect 16420 -6690 16480 -6650
rect 16420 -6770 16480 -6730
rect 16420 -6850 16480 -6810
rect 16420 -6930 16480 -6890
rect 16810 -6530 16870 -6490
rect 16810 -6610 16870 -6570
rect 16810 -6690 16870 -6650
rect 16810 -6770 16870 -6730
rect 16810 -6850 16870 -6810
rect 16810 -6930 16870 -6890
rect 17200 -6530 17260 -6490
rect 17200 -6610 17260 -6570
rect 17200 -6690 17260 -6650
rect 17200 -6770 17260 -6730
rect 17200 -6850 17260 -6810
rect 17200 -6930 17260 -6890
rect -250 -9700 -210 -9660
rect -170 -9700 -130 -9660
rect -90 -9700 -50 -9660
rect -10 -9700 30 -9660
rect 70 -9700 110 -9660
rect 150 -9700 190 -9660
rect -250 -9780 -210 -9740
rect -170 -9780 -130 -9740
rect -90 -9780 -50 -9740
rect -10 -9780 30 -9740
rect 70 -9780 110 -9740
rect 150 -9780 190 -9740
rect -250 -9860 -210 -9820
rect -170 -9860 -130 -9820
rect -90 -9860 -50 -9820
rect -10 -9860 30 -9820
rect 70 -9860 110 -9820
rect 150 -9860 190 -9820
rect 7230 -9700 7270 -9660
rect 7310 -9700 7350 -9660
rect 7390 -9700 7430 -9660
rect 7470 -9700 7510 -9660
rect 7550 -9700 7590 -9660
rect 7630 -9700 7670 -9660
rect 7230 -9780 7270 -9740
rect 7310 -9780 7350 -9740
rect 7390 -9780 7430 -9740
rect 7470 -9780 7510 -9740
rect 7550 -9780 7590 -9740
rect 7630 -9780 7670 -9740
rect 7230 -9860 7270 -9820
rect 7310 -9860 7350 -9820
rect 7390 -9860 7430 -9820
rect 7470 -9860 7510 -9820
rect 7550 -9860 7590 -9820
rect 7630 -9860 7670 -9820
rect 14710 -9700 14750 -9660
rect 14790 -9700 14830 -9660
rect 14870 -9700 14910 -9660
rect 14950 -9700 14990 -9660
rect 15030 -9700 15070 -9660
rect 15110 -9700 15150 -9660
rect 14710 -9780 14750 -9740
rect 14790 -9780 14830 -9740
rect 14870 -9780 14910 -9740
rect 14950 -9780 14990 -9740
rect 15030 -9780 15070 -9740
rect 15110 -9780 15150 -9740
rect 14710 -9860 14750 -9820
rect 14790 -9860 14830 -9820
rect 14870 -9860 14910 -9820
rect 14950 -9860 14990 -9820
rect 15030 -9860 15070 -9820
rect 15110 -9860 15150 -9820
<< metal1 >>
rect 23460 7210 23940 7230
rect 23460 7140 23490 7210
rect 23560 7140 23600 7210
rect 23670 7140 23710 7210
rect 23780 7140 23820 7210
rect 23890 7140 23940 7210
rect 23460 7100 23940 7140
rect 23460 7030 23490 7100
rect 23560 7030 23600 7100
rect 23670 7030 23710 7100
rect 23780 7030 23820 7100
rect 23890 7030 23940 7100
rect 23460 6920 23940 7030
rect 25860 7210 26340 7230
rect 25860 7140 25890 7210
rect 25960 7140 26000 7210
rect 26070 7140 26110 7210
rect 26180 7140 26220 7210
rect 26290 7140 26340 7210
rect 25860 7100 26340 7140
rect 25860 7030 25890 7100
rect 25960 7030 26000 7100
rect 26070 7030 26110 7100
rect 26180 7030 26220 7100
rect 26290 7030 26340 7100
rect 25860 6950 26340 7030
rect 11760 6880 13360 6900
rect 1540 6850 3140 6870
rect 1540 6780 1570 6850
rect 1640 6780 1680 6850
rect 1750 6780 1790 6850
rect 1860 6780 1900 6850
rect 1970 6780 2010 6850
rect 2080 6780 2120 6850
rect 2190 6780 2230 6850
rect 2300 6780 2340 6850
rect 2410 6780 2450 6850
rect 2520 6780 2560 6850
rect 2630 6780 2670 6850
rect 2740 6780 2780 6850
rect 2850 6780 2890 6850
rect 2960 6780 3000 6850
rect 3070 6780 3140 6850
rect 1540 6740 3140 6780
rect 1540 6670 1570 6740
rect 1640 6670 1680 6740
rect 1750 6670 1790 6740
rect 1860 6670 1900 6740
rect 1970 6670 2010 6740
rect 2080 6670 2120 6740
rect 2190 6670 2230 6740
rect 2300 6670 2340 6740
rect 2410 6670 2450 6740
rect 2520 6670 2560 6740
rect 2630 6670 2670 6740
rect 2740 6670 2780 6740
rect 2850 6670 2890 6740
rect 2960 6670 3000 6740
rect 3070 6670 3140 6740
rect 1540 6520 3140 6670
rect 11760 6810 11790 6880
rect 11860 6810 11900 6880
rect 11970 6810 12010 6880
rect 12080 6810 12120 6880
rect 12190 6810 12230 6880
rect 12300 6810 12340 6880
rect 12410 6810 12450 6880
rect 12520 6810 12560 6880
rect 12630 6810 12670 6880
rect 12740 6810 12780 6880
rect 12850 6810 12890 6880
rect 12960 6810 13000 6880
rect 13070 6810 13110 6880
rect 13180 6810 13220 6880
rect 13290 6810 13360 6880
rect 11760 6770 13360 6810
rect 11760 6700 11790 6770
rect 11860 6700 11900 6770
rect 11970 6700 12010 6770
rect 12080 6700 12120 6770
rect 12190 6700 12230 6770
rect 12300 6700 12340 6770
rect 12410 6700 12450 6770
rect 12520 6700 12560 6770
rect 12630 6700 12670 6770
rect 12740 6700 12780 6770
rect 12850 6700 12890 6770
rect 12960 6700 13000 6770
rect 13070 6700 13110 6770
rect 13180 6700 13220 6770
rect 13290 6700 13360 6770
rect 11760 6550 13360 6700
rect 21800 5670 22120 5690
rect 21800 5600 21820 5670
rect 21890 5600 21930 5670
rect 22000 5600 22120 5670
rect 21800 5560 22120 5600
rect 21800 5490 21820 5560
rect 21890 5490 21930 5560
rect 22000 5490 22120 5560
rect 21800 5450 22120 5490
rect 7400 5390 7490 5410
rect 7400 5320 7410 5390
rect 7480 5320 7490 5390
rect 7400 5280 7490 5320
rect 7400 5210 7410 5280
rect 7480 5210 7490 5280
rect 7400 5170 7490 5210
rect 7400 5100 7410 5170
rect 7480 5100 7490 5170
rect 7400 5060 7490 5100
rect 7400 4990 7410 5060
rect 7480 4990 7490 5060
rect 7400 4950 7490 4990
rect 7400 4880 7410 4950
rect 7480 4880 7490 4950
rect 7400 4860 7490 4880
rect 21800 5380 21820 5450
rect 21890 5380 21930 5450
rect 22000 5380 22120 5450
rect 21800 5340 22120 5380
rect 21800 5270 21820 5340
rect 21890 5270 21930 5340
rect 22000 5270 22120 5340
rect 21800 5230 22120 5270
rect 21800 5160 21820 5230
rect 21890 5160 21930 5230
rect 22000 5160 22120 5230
rect 21800 5120 22120 5160
rect 21800 5050 21820 5120
rect 21890 5050 21930 5120
rect 22000 5050 22120 5120
rect 21800 5010 22120 5050
rect 21800 4940 21820 5010
rect 21890 4940 21930 5010
rect 22000 4940 22120 5010
rect 21800 4900 22120 4940
rect 21800 4830 21820 4900
rect 21890 4830 21930 4900
rect 22000 4830 22120 4900
rect 21800 4790 22120 4830
rect 21800 4720 21820 4790
rect 21890 4720 21930 4790
rect 22000 4720 22120 4790
rect 21800 4680 22120 4720
rect 21800 4610 21820 4680
rect 21890 4610 21930 4680
rect 22000 4610 22120 4680
rect -2520 4590 -2380 4610
rect -2520 4580 -2480 4590
rect -2520 4510 -2490 4580
rect -2520 4470 -2480 4510
rect -2520 4400 -2490 4470
rect -2520 4390 -2480 4400
rect -2420 4390 -2380 4590
rect -2520 4360 -2380 4390
rect -2520 4290 -2490 4360
rect -2420 4290 -2380 4360
rect -2520 4270 -2380 4290
rect -2520 4250 -2480 4270
rect -2520 4180 -2490 4250
rect -2520 4150 -2480 4180
rect -2420 4150 -2380 4270
rect -2520 4130 -2380 4150
rect -2130 4590 -1600 4610
rect -2130 4550 -2090 4590
rect -2030 4550 -1700 4590
rect -1640 4550 -1600 4590
rect -2130 4510 -1600 4550
rect -2130 4470 -2090 4510
rect -2030 4470 -1700 4510
rect -1640 4470 -1600 4510
rect -2130 4430 -1600 4470
rect -2130 4390 -2090 4430
rect -2030 4390 -1700 4430
rect -1640 4390 -1600 4430
rect -2130 4350 -1600 4390
rect -2130 4310 -2090 4350
rect -2030 4310 -1700 4350
rect -1640 4310 -1600 4350
rect -2130 4270 -1600 4310
rect -2130 4230 -2090 4270
rect -2030 4230 -1700 4270
rect -1640 4230 -1600 4270
rect -2130 4190 -1600 4230
rect -2130 4150 -2090 4190
rect -2030 4150 -1700 4190
rect -1640 4150 -1600 4190
rect -2130 4130 -1600 4150
rect 16380 4590 16910 4610
rect 16380 4550 16420 4590
rect 16480 4550 16810 4590
rect 16870 4550 16910 4590
rect 16380 4510 16910 4550
rect 16380 4470 16420 4510
rect 16480 4470 16810 4510
rect 16870 4470 16910 4510
rect 16380 4430 16910 4470
rect 16380 4390 16420 4430
rect 16480 4390 16810 4430
rect 16870 4390 16910 4430
rect 16380 4350 16910 4390
rect 16380 4310 16420 4350
rect 16480 4310 16810 4350
rect 16870 4310 16910 4350
rect 16380 4270 16910 4310
rect 16380 4230 16420 4270
rect 16480 4230 16810 4270
rect 16870 4230 16910 4270
rect 16380 4190 16910 4230
rect 16380 4150 16420 4190
rect 16480 4150 16810 4190
rect 16870 4150 16910 4190
rect 16380 4130 16910 4150
rect 17160 4590 17300 4610
rect 17160 4390 17200 4590
rect 17260 4580 17300 4590
rect 17270 4510 17300 4580
rect 17260 4470 17300 4510
rect 17270 4400 17300 4470
rect 17260 4390 17300 4400
rect 17160 4360 17300 4390
rect 17160 4290 17200 4360
rect 17270 4290 17300 4360
rect 17160 4270 17300 4290
rect 17160 4150 17200 4270
rect 17260 4250 17300 4270
rect 17270 4180 17300 4250
rect 17260 4150 17300 4180
rect 17160 4130 17300 4150
rect 21800 4570 22120 4610
rect 21800 4500 21820 4570
rect 21890 4500 21930 4570
rect 22000 4500 22120 4570
rect 21800 3990 22120 4500
rect 24700 3360 25030 3380
rect 24700 3290 24720 3360
rect 24790 3290 24830 3360
rect 24900 3290 24940 3360
rect 25010 3290 25030 3360
rect 24700 3250 25030 3290
rect 24700 3180 24720 3250
rect 24790 3180 24830 3250
rect 24900 3180 24940 3250
rect 25010 3180 25030 3250
rect 24700 3140 25030 3180
rect 24700 3070 24720 3140
rect 24790 3070 24830 3140
rect 24900 3070 24940 3140
rect 25010 3070 25030 3140
rect 24700 3050 25030 3070
rect 22420 2600 22900 2670
rect 22420 2530 22470 2600
rect 22540 2530 22580 2600
rect 22650 2530 22690 2600
rect 22760 2530 22800 2600
rect 22870 2530 22900 2600
rect 22420 2490 22900 2530
rect 22420 2420 22470 2490
rect 22540 2420 22580 2490
rect 22650 2420 22690 2490
rect 22760 2420 22800 2490
rect 22870 2420 22900 2490
rect 22420 2400 22900 2420
rect 26900 2600 27380 2660
rect 26900 2530 26950 2600
rect 27020 2530 27060 2600
rect 27130 2530 27170 2600
rect 27240 2530 27280 2600
rect 27350 2530 27380 2600
rect 26900 2490 27380 2530
rect 26900 2420 26950 2490
rect 27020 2420 27060 2490
rect 27130 2420 27170 2490
rect 27240 2420 27280 2490
rect 27350 2420 27380 2490
rect 26900 2400 27380 2420
rect 0 1160 310 1180
rect 0 1090 20 1160
rect 90 1090 130 1160
rect 200 1090 230 1160
rect 300 1090 310 1160
rect 0 1050 310 1090
rect 0 980 20 1050
rect 90 980 130 1050
rect 200 980 230 1050
rect 300 980 310 1050
rect 0 940 310 980
rect 0 870 20 940
rect 90 870 130 940
rect 200 870 230 940
rect 300 870 310 940
rect 0 850 310 870
rect 14590 1160 14900 1180
rect 14590 1090 14600 1160
rect 14670 1090 14700 1160
rect 14770 1090 14810 1160
rect 14880 1090 14900 1160
rect 14590 1050 14900 1090
rect 14590 980 14600 1050
rect 14670 980 14700 1050
rect 14770 980 14810 1050
rect 14880 980 14900 1050
rect 14590 940 14900 980
rect 14590 870 14600 940
rect 14670 870 14700 940
rect 14770 870 14810 940
rect 14880 870 14900 940
rect 14590 850 14900 870
rect 23460 920 23940 940
rect 23460 850 23490 920
rect 23560 850 23600 920
rect 23670 850 23710 920
rect 23780 850 23820 920
rect 23890 850 23940 920
rect 23460 810 23940 850
rect 23460 740 23490 810
rect 23560 740 23600 810
rect 23670 740 23710 810
rect 23780 740 23820 810
rect 23890 740 23940 810
rect 23460 640 23940 740
rect 25860 920 26340 940
rect 25860 850 25890 920
rect 25960 850 26000 920
rect 26070 850 26110 920
rect 26180 850 26220 920
rect 26290 850 26340 920
rect 25860 810 26340 850
rect 25860 740 25890 810
rect 25960 740 26000 810
rect 26070 740 26110 810
rect 26180 740 26220 810
rect 26290 740 26340 810
rect 25860 650 26340 740
rect -330 -140 150 -98
rect -330 -180 -310 -140
rect -110 -180 -80 -140
rect -10 -180 10 -140
rect 130 -180 150 -140
rect -330 -210 -300 -180
rect -230 -210 -190 -180
rect -120 -210 -80 -180
rect -10 -210 30 -180
rect 100 -210 150 -180
rect -330 -220 150 -210
rect -330 -260 -310 -220
rect -270 -260 -230 -220
rect -190 -260 -150 -220
rect -110 -260 -70 -220
rect -30 -260 10 -220
rect 50 -260 90 -220
rect 130 -260 150 -220
rect -330 -270 150 -260
rect -330 -300 -300 -270
rect -230 -300 -190 -270
rect -120 -300 -80 -270
rect -10 -300 30 -270
rect 100 -300 150 -270
rect -330 -340 -310 -300
rect -110 -340 -80 -300
rect -10 -340 10 -300
rect 130 -340 150 -300
rect -330 -380 150 -340
rect 1080 -790 2680 40
rect 7150 -120 7630 -98
rect 7150 -140 7180 -120
rect 7240 -140 7280 -120
rect 7340 -140 7440 -120
rect 7500 -140 7540 -120
rect 7600 -140 7630 -120
rect 7150 -180 7170 -140
rect 7240 -180 7250 -140
rect 7370 -180 7410 -140
rect 7530 -180 7540 -140
rect 7610 -180 7630 -140
rect 7150 -210 7630 -180
rect 7150 -220 7180 -210
rect 7240 -220 7280 -210
rect 7340 -220 7440 -210
rect 7500 -220 7540 -210
rect 7600 -220 7630 -210
rect 7150 -260 7170 -220
rect 7240 -260 7250 -220
rect 7370 -260 7410 -220
rect 7530 -260 7540 -220
rect 7610 -260 7630 -220
rect 7150 -270 7180 -260
rect 7240 -270 7280 -260
rect 7340 -270 7440 -260
rect 7500 -270 7540 -260
rect 7600 -270 7630 -260
rect 7150 -300 7630 -270
rect 7150 -340 7170 -300
rect 7240 -340 7250 -300
rect 7370 -340 7410 -300
rect 7530 -340 7540 -300
rect 7610 -340 7630 -300
rect 7150 -360 7180 -340
rect 7240 -360 7280 -340
rect 7340 -360 7440 -340
rect 7500 -360 7540 -340
rect 7600 -360 7630 -340
rect 7150 -380 7630 -360
rect 1080 -860 1150 -790
rect 1220 -860 1260 -790
rect 1330 -860 1370 -790
rect 1440 -860 1480 -790
rect 1550 -860 1590 -790
rect 1660 -860 1700 -790
rect 1770 -860 1810 -790
rect 1880 -860 1920 -790
rect 1990 -860 2030 -790
rect 2100 -860 2140 -790
rect 2210 -860 2250 -790
rect 2320 -860 2360 -790
rect 2430 -860 2470 -790
rect 2540 -860 2580 -790
rect 2650 -860 2680 -790
rect 1080 -900 2680 -860
rect 1080 -970 1150 -900
rect 1220 -970 1260 -900
rect 1330 -970 1370 -900
rect 1440 -970 1480 -900
rect 1550 -970 1590 -900
rect 1660 -970 1700 -900
rect 1770 -970 1810 -900
rect 1880 -970 1920 -900
rect 1990 -970 2030 -900
rect 2100 -970 2140 -900
rect 2210 -970 2250 -900
rect 2320 -970 2360 -900
rect 2430 -970 2470 -900
rect 2540 -970 2580 -900
rect 2650 -970 2680 -900
rect 1080 -990 2680 -970
rect 12220 -790 13820 40
rect 14630 -140 15110 -98
rect 14630 -180 14650 -140
rect 14850 -180 14880 -140
rect 14950 -180 14970 -140
rect 15090 -180 15110 -140
rect 14630 -210 14660 -180
rect 14730 -210 14770 -180
rect 14840 -210 14880 -180
rect 14950 -210 14990 -180
rect 15060 -210 15110 -180
rect 14630 -220 15110 -210
rect 14630 -260 14650 -220
rect 14690 -260 14730 -220
rect 14770 -260 14810 -220
rect 14850 -260 14890 -220
rect 14930 -260 14970 -220
rect 15010 -260 15050 -220
rect 15090 -260 15110 -220
rect 14630 -270 15110 -260
rect 14630 -300 14660 -270
rect 14730 -300 14770 -270
rect 14840 -300 14880 -270
rect 14950 -300 14990 -270
rect 15060 -300 15110 -270
rect 14630 -340 14650 -300
rect 14850 -340 14880 -300
rect 14950 -340 14970 -300
rect 15090 -340 15110 -300
rect 14630 -380 15110 -340
rect 12220 -860 12250 -790
rect 12320 -860 12360 -790
rect 12430 -860 12470 -790
rect 12540 -860 12580 -790
rect 12650 -860 12690 -790
rect 12760 -860 12800 -790
rect 12870 -860 12910 -790
rect 12980 -860 13020 -790
rect 13090 -860 13130 -790
rect 13200 -860 13240 -790
rect 13310 -860 13350 -790
rect 13420 -860 13460 -790
rect 13530 -860 13570 -790
rect 13640 -860 13680 -790
rect 13750 -860 13820 -790
rect 12220 -900 13820 -860
rect 12220 -970 12250 -900
rect 12320 -970 12360 -900
rect 12430 -970 12470 -900
rect 12540 -970 12580 -900
rect 12650 -970 12690 -900
rect 12760 -970 12800 -900
rect 12870 -970 12910 -900
rect 12980 -970 13020 -900
rect 13090 -970 13130 -900
rect 13200 -970 13240 -900
rect 13310 -970 13350 -900
rect 13420 -970 13460 -900
rect 13530 -970 13570 -900
rect 13640 -970 13680 -900
rect 13750 -970 13820 -900
rect 12220 -990 13820 -970
rect 21800 -850 22060 -820
rect 21800 -920 21820 -850
rect 21890 -920 21930 -850
rect 22000 -920 22060 -850
rect 21800 -960 22060 -920
rect 21800 -1030 21820 -960
rect 21890 -1030 21930 -960
rect 22000 -1030 22060 -960
rect 21800 -1070 22060 -1030
rect 21800 -1140 21820 -1070
rect 21890 -1140 21930 -1070
rect 22000 -1140 22060 -1070
rect 21800 -1180 22060 -1140
rect 21800 -1250 21820 -1180
rect 21890 -1250 21930 -1180
rect 22000 -1250 22060 -1180
rect 21800 -1290 22060 -1250
rect 21800 -1360 21820 -1290
rect 21890 -1360 21930 -1290
rect 22000 -1360 22060 -1290
rect 21800 -1400 22060 -1360
rect 21800 -1470 21820 -1400
rect 21890 -1470 21930 -1400
rect 22000 -1470 22060 -1400
rect 21800 -1510 22060 -1470
rect 21800 -1580 21820 -1510
rect 21890 -1580 21930 -1510
rect 22000 -1580 22060 -1510
rect 21800 -1620 22060 -1580
rect 21800 -1690 21820 -1620
rect 21890 -1690 21930 -1620
rect 22000 -1690 22060 -1620
rect 21800 -1730 22060 -1690
rect 21800 -1800 21820 -1730
rect 21890 -1800 21930 -1730
rect 22000 -1800 22060 -1730
rect 21800 -1840 22060 -1800
rect 21800 -1910 21820 -1840
rect 21890 -1910 21930 -1840
rect 22000 -1910 22060 -1840
rect 21800 -1950 22060 -1910
rect 21800 -2020 21820 -1950
rect 21890 -2020 21930 -1950
rect 22000 -2020 22060 -1950
rect 21800 -2040 22060 -2020
rect 1540 -2780 3140 -2760
rect 1540 -2850 1570 -2780
rect 1640 -2850 1680 -2780
rect 1750 -2850 1790 -2780
rect 1860 -2850 1900 -2780
rect 1970 -2850 2010 -2780
rect 2080 -2850 2120 -2780
rect 2190 -2850 2230 -2780
rect 2300 -2850 2340 -2780
rect 2410 -2850 2450 -2780
rect 2520 -2850 2560 -2780
rect 2630 -2850 2670 -2780
rect 2740 -2850 2780 -2780
rect 2850 -2850 2890 -2780
rect 2960 -2850 3000 -2780
rect 3070 -2850 3140 -2780
rect 1540 -2890 3140 -2850
rect 1540 -2960 1570 -2890
rect 1640 -2960 1680 -2890
rect 1750 -2960 1790 -2890
rect 1860 -2960 1900 -2890
rect 1970 -2960 2010 -2890
rect 2080 -2960 2120 -2890
rect 2190 -2960 2230 -2890
rect 2300 -2960 2340 -2890
rect 2410 -2960 2450 -2890
rect 2520 -2960 2560 -2890
rect 2630 -2960 2670 -2890
rect 2740 -2960 2780 -2890
rect 2850 -2960 2890 -2890
rect 2960 -2960 3000 -2890
rect 3070 -2960 3140 -2890
rect 1540 -3020 3140 -2960
rect 11760 -2780 13360 -2760
rect 11760 -2850 11790 -2780
rect 11860 -2850 11900 -2780
rect 11970 -2850 12010 -2780
rect 12080 -2850 12120 -2780
rect 12190 -2850 12230 -2780
rect 12300 -2850 12340 -2780
rect 12410 -2850 12450 -2780
rect 12520 -2850 12560 -2780
rect 12630 -2850 12670 -2780
rect 12740 -2850 12780 -2780
rect 12850 -2850 12890 -2780
rect 12960 -2850 13000 -2780
rect 13070 -2850 13110 -2780
rect 13180 -2850 13220 -2780
rect 13290 -2850 13360 -2780
rect 11760 -2890 13360 -2850
rect 11760 -2960 11790 -2890
rect 11860 -2960 11900 -2890
rect 11970 -2960 12010 -2890
rect 12080 -2960 12120 -2890
rect 12190 -2960 12230 -2890
rect 12300 -2960 12340 -2890
rect 12410 -2960 12450 -2890
rect 12520 -2960 12560 -2890
rect 12630 -2960 12670 -2890
rect 12740 -2960 12780 -2890
rect 12850 -2960 12890 -2890
rect 12960 -2960 13000 -2890
rect 13070 -2960 13110 -2890
rect 13180 -2960 13220 -2890
rect 13290 -2960 13360 -2890
rect 11760 -3020 13360 -2960
rect 24720 -3050 25050 -3030
rect 24720 -3120 24740 -3050
rect 24810 -3120 24850 -3050
rect 24920 -3120 24960 -3050
rect 25030 -3120 25050 -3050
rect 24720 -3160 25050 -3120
rect 24720 -3230 24740 -3160
rect 24810 -3230 24850 -3160
rect 24920 -3230 24960 -3160
rect 25030 -3230 25050 -3160
rect 24720 -3270 25050 -3230
rect 24720 -3340 24740 -3270
rect 24810 -3340 24850 -3270
rect 24920 -3340 24960 -3270
rect 25030 -3340 25050 -3270
rect 24720 -3360 25050 -3340
rect 22420 -3690 22900 -3630
rect 22420 -3760 22470 -3690
rect 22540 -3760 22580 -3690
rect 22650 -3760 22690 -3690
rect 22760 -3760 22800 -3690
rect 22870 -3760 22900 -3690
rect 22420 -3800 22900 -3760
rect 7290 -3880 7620 -3860
rect 7290 -3950 7310 -3880
rect 7380 -3950 7420 -3880
rect 7490 -3950 7530 -3880
rect 7600 -3950 7620 -3880
rect 22420 -3870 22470 -3800
rect 22540 -3870 22580 -3800
rect 22650 -3870 22690 -3800
rect 22760 -3870 22800 -3800
rect 22870 -3870 22900 -3800
rect 22420 -3890 22900 -3870
rect 26900 -3690 27380 -3630
rect 26900 -3760 26950 -3690
rect 27020 -3760 27060 -3690
rect 27130 -3760 27170 -3690
rect 27240 -3760 27280 -3690
rect 27350 -3760 27380 -3690
rect 26900 -3800 27380 -3760
rect 26900 -3870 26950 -3800
rect 27020 -3870 27060 -3800
rect 27130 -3870 27170 -3800
rect 27240 -3870 27280 -3800
rect 27350 -3870 27380 -3800
rect 26900 -3890 27380 -3870
rect 7290 -3990 7620 -3950
rect 7290 -4060 7310 -3990
rect 7380 -4060 7420 -3990
rect 7490 -4060 7530 -3990
rect 7600 -4060 7620 -3990
rect 7290 -4100 7620 -4060
rect 7290 -4170 7310 -4100
rect 7380 -4170 7420 -4100
rect 7490 -4170 7530 -4100
rect 7600 -4170 7620 -4100
rect 7290 -4190 7620 -4170
rect -1350 -4312 -870 -4270
rect -1350 -4432 -1330 -4312
rect -1290 -4350 -1250 -4312
rect -1210 -4350 -1170 -4312
rect -1130 -4350 -1090 -4312
rect -1050 -4350 -1010 -4312
rect -970 -4350 -930 -4312
rect -1260 -4352 -1250 -4350
rect -1130 -4352 -1110 -4350
rect -1040 -4352 -1010 -4350
rect -890 -4352 -870 -4312
rect -1260 -4392 -1220 -4352
rect -1150 -4392 -1110 -4352
rect -1040 -4392 -1000 -4352
rect -930 -4392 -870 -4352
rect -1260 -4420 -1250 -4392
rect -1130 -4420 -1110 -4392
rect -1040 -4420 -1010 -4392
rect -1290 -4432 -1250 -4420
rect -1210 -4432 -1170 -4420
rect -1130 -4432 -1090 -4420
rect -1050 -4432 -1010 -4420
rect -970 -4432 -930 -4420
rect -890 -4432 -870 -4392
rect -1350 -4460 -870 -4432
rect -1350 -4530 -1330 -4460
rect -1260 -4472 -1220 -4460
rect -1150 -4472 -1110 -4460
rect -1040 -4472 -1000 -4460
rect -930 -4472 -870 -4460
rect -1260 -4512 -1250 -4472
rect -1130 -4512 -1110 -4472
rect -1040 -4512 -1010 -4472
rect -890 -4512 -870 -4472
rect -1260 -4530 -1220 -4512
rect -1150 -4530 -1110 -4512
rect -1040 -4530 -1000 -4512
rect -930 -4530 -870 -4512
rect -1350 -4552 -870 -4530
rect -588 -4290 -110 -4270
rect -588 -4312 -560 -4290
rect -490 -4312 -450 -4290
rect -380 -4312 -340 -4290
rect -270 -4312 -230 -4290
rect -160 -4312 -110 -4290
rect -588 -4352 -570 -4312
rect -370 -4352 -340 -4312
rect -270 -4352 -250 -4312
rect -130 -4352 -110 -4312
rect -588 -4360 -560 -4352
rect -490 -4360 -450 -4352
rect -380 -4360 -340 -4352
rect -270 -4360 -230 -4352
rect -160 -4360 -110 -4352
rect -588 -4392 -110 -4360
rect -588 -4432 -570 -4392
rect -530 -4400 -490 -4392
rect -450 -4400 -410 -4392
rect -370 -4400 -330 -4392
rect -290 -4400 -250 -4392
rect -210 -4400 -170 -4392
rect -370 -4432 -340 -4400
rect -270 -4432 -250 -4400
rect -130 -4432 -110 -4392
rect -588 -4470 -560 -4432
rect -490 -4470 -450 -4432
rect -380 -4470 -340 -4432
rect -270 -4470 -230 -4432
rect -160 -4470 -110 -4432
rect -588 -4472 -110 -4470
rect -588 -4512 -570 -4472
rect -530 -4512 -490 -4472
rect -450 -4512 -410 -4472
rect -370 -4512 -330 -4472
rect -290 -4512 -250 -4472
rect -210 -4512 -170 -4472
rect -130 -4512 -110 -4472
rect -588 -4552 -110 -4512
rect 14890 -4290 15368 -4270
rect 14890 -4312 14940 -4290
rect 15010 -4312 15050 -4290
rect 15120 -4312 15160 -4290
rect 15230 -4312 15270 -4290
rect 15340 -4312 15368 -4290
rect 14890 -4352 14910 -4312
rect 15030 -4352 15050 -4312
rect 15120 -4352 15150 -4312
rect 15350 -4352 15368 -4312
rect 14890 -4360 14940 -4352
rect 15010 -4360 15050 -4352
rect 15120 -4360 15160 -4352
rect 15230 -4360 15270 -4352
rect 15340 -4360 15368 -4352
rect 14890 -4392 15368 -4360
rect 14890 -4432 14910 -4392
rect 14950 -4400 14990 -4392
rect 15030 -4400 15070 -4392
rect 15110 -4400 15150 -4392
rect 15190 -4400 15230 -4392
rect 15030 -4432 15050 -4400
rect 15120 -4432 15150 -4400
rect 15270 -4400 15310 -4392
rect 15350 -4432 15368 -4392
rect 14890 -4470 14940 -4432
rect 15010 -4470 15050 -4432
rect 15120 -4470 15160 -4432
rect 15230 -4470 15270 -4432
rect 15340 -4470 15368 -4432
rect 14890 -4472 15368 -4470
rect 14890 -4512 14910 -4472
rect 14950 -4512 14990 -4472
rect 15030 -4512 15070 -4472
rect 15110 -4512 15150 -4472
rect 15190 -4512 15230 -4472
rect 15270 -4512 15310 -4472
rect 15350 -4512 15368 -4472
rect 14890 -4552 15368 -4512
rect 15650 -4312 16130 -4270
rect 15650 -4352 15670 -4312
rect 15710 -4350 15750 -4312
rect 15790 -4350 15830 -4312
rect 15870 -4350 15910 -4312
rect 15950 -4350 15990 -4312
rect 16030 -4350 16070 -4312
rect 15790 -4352 15820 -4350
rect 15890 -4352 15910 -4350
rect 16030 -4352 16040 -4350
rect 15650 -4392 15710 -4352
rect 15780 -4392 15820 -4352
rect 15890 -4392 15930 -4352
rect 16000 -4392 16040 -4352
rect 15650 -4432 15670 -4392
rect 15790 -4420 15820 -4392
rect 15890 -4420 15910 -4392
rect 16030 -4420 16040 -4392
rect 15710 -4432 15750 -4420
rect 15790 -4432 15830 -4420
rect 15870 -4432 15910 -4420
rect 15950 -4432 15990 -4420
rect 16030 -4432 16070 -4420
rect 16110 -4432 16130 -4312
rect 15650 -4460 16130 -4432
rect 15650 -4472 15710 -4460
rect 15780 -4472 15820 -4460
rect 15890 -4472 15930 -4460
rect 16000 -4472 16040 -4460
rect 15650 -4512 15670 -4472
rect 15790 -4512 15820 -4472
rect 15890 -4512 15910 -4472
rect 16030 -4512 16040 -4472
rect 15650 -4530 15710 -4512
rect 15780 -4530 15820 -4512
rect 15890 -4530 15930 -4512
rect 16000 -4530 16040 -4512
rect 16110 -4530 16130 -4460
rect 15650 -4552 16130 -4530
rect 7570 -6460 7870 -6420
rect -2520 -6490 -1990 -6470
rect -2520 -6530 -2480 -6490
rect -2420 -6530 -2090 -6490
rect -2030 -6530 -1990 -6490
rect -2520 -6570 -1990 -6530
rect -2520 -6610 -2480 -6570
rect -2420 -6610 -2090 -6570
rect -2030 -6610 -1990 -6570
rect -2520 -6650 -1990 -6610
rect -2520 -6690 -2480 -6650
rect -2420 -6690 -2090 -6650
rect -2030 -6690 -1990 -6650
rect -2520 -6730 -1990 -6690
rect -2520 -6770 -2480 -6730
rect -2420 -6770 -2090 -6730
rect -2030 -6770 -1990 -6730
rect -2520 -6810 -1990 -6770
rect -2520 -6850 -2480 -6810
rect -2420 -6850 -2090 -6810
rect -2030 -6850 -1990 -6810
rect -2520 -6890 -1990 -6850
rect -2520 -6930 -2480 -6890
rect -2420 -6930 -2090 -6890
rect -2030 -6930 -1990 -6890
rect -2520 -6950 -1990 -6930
rect -1740 -6490 -1600 -6470
rect -1740 -6520 -1700 -6490
rect -1740 -6590 -1710 -6520
rect -1740 -6610 -1700 -6590
rect -1640 -6610 -1600 -6490
rect 7570 -6520 7590 -6460
rect 7650 -6520 7690 -6460
rect 7750 -6520 7790 -6460
rect 7850 -6520 7870 -6460
rect 7570 -6560 7870 -6520
rect -1740 -6630 -1600 -6610
rect 7570 -6620 7590 -6560
rect 7650 -6620 7690 -6560
rect 7750 -6620 7790 -6560
rect 7850 -6620 7870 -6560
rect -1740 -6700 -1710 -6630
rect -1640 -6700 -1600 -6630
rect 7570 -6660 7870 -6620
rect -1740 -6730 -1600 -6700
rect 7570 -6720 7590 -6660
rect 7650 -6720 7690 -6660
rect 7750 -6720 7790 -6660
rect 7850 -6720 7870 -6660
rect 16380 -6490 16520 -6470
rect 16380 -6610 16420 -6490
rect 16480 -6520 16520 -6490
rect 16490 -6590 16520 -6520
rect 16480 -6610 16520 -6590
rect 16380 -6630 16520 -6610
rect -1740 -6740 -1700 -6730
rect -1740 -6810 -1710 -6740
rect -1740 -6850 -1700 -6810
rect -1740 -6920 -1710 -6850
rect -1740 -6930 -1700 -6920
rect -1640 -6930 -1600 -6730
rect 7570 -6760 7870 -6720
rect 16380 -6700 16420 -6630
rect 16490 -6700 16520 -6630
rect 16380 -6730 16520 -6700
rect 7570 -6820 7590 -6760
rect 7650 -6820 7690 -6760
rect 7750 -6820 7790 -6760
rect 7850 -6820 7870 -6760
rect 7570 -6850 7870 -6820
rect 16380 -6930 16420 -6730
rect 16480 -6740 16520 -6730
rect 16490 -6810 16520 -6740
rect 16480 -6850 16520 -6810
rect 16490 -6920 16520 -6850
rect 16480 -6930 16520 -6920
rect -1740 -6950 -1600 -6930
rect 16380 -6950 16520 -6930
rect 16770 -6490 17300 -6470
rect 16770 -6530 16810 -6490
rect 16870 -6530 17200 -6490
rect 17260 -6530 17300 -6490
rect 16770 -6570 17300 -6530
rect 16770 -6610 16810 -6570
rect 16870 -6610 17200 -6570
rect 17260 -6610 17300 -6570
rect 16770 -6650 17300 -6610
rect 16770 -6690 16810 -6650
rect 16870 -6690 17200 -6650
rect 17260 -6690 17300 -6650
rect 16770 -6730 17300 -6690
rect 16770 -6770 16810 -6730
rect 16870 -6770 17200 -6730
rect 17260 -6770 17300 -6730
rect 16770 -6810 17300 -6770
rect 16770 -6850 16810 -6810
rect 16870 -6850 17200 -6810
rect 17260 -6850 17300 -6810
rect 16770 -6890 17300 -6850
rect 16770 -6930 16810 -6890
rect 16870 -6930 17200 -6890
rect 17260 -6930 17300 -6890
rect 16770 -6950 17300 -6930
rect 0 -8140 310 -8120
rect 0 -8210 20 -8140
rect 90 -8210 130 -8140
rect 200 -8210 230 -8140
rect 300 -8210 310 -8140
rect 0 -8250 310 -8210
rect 0 -8320 20 -8250
rect 90 -8320 130 -8250
rect 200 -8320 230 -8250
rect 300 -8320 310 -8250
rect 0 -8360 310 -8320
rect 0 -8430 20 -8360
rect 90 -8430 130 -8360
rect 200 -8430 230 -8360
rect 300 -8430 310 -8360
rect 0 -8450 310 -8430
rect 14590 -8230 14900 -8210
rect 14590 -8300 14600 -8230
rect 14670 -8300 14700 -8230
rect 14770 -8300 14810 -8230
rect 14880 -8300 14900 -8230
rect 14590 -8340 14900 -8300
rect 14590 -8410 14600 -8340
rect 14670 -8410 14700 -8340
rect 14770 -8410 14810 -8340
rect 14880 -8410 14900 -8340
rect 14590 -8450 14900 -8410
rect 14590 -8520 14600 -8450
rect 14670 -8520 14700 -8450
rect 14770 -8520 14810 -8450
rect 14880 -8520 14900 -8450
rect 14590 -8540 14900 -8520
rect 21610 -8360 22540 -8330
rect 21610 -8430 21630 -8360
rect 21700 -8430 21730 -8360
rect 21800 -8430 21830 -8360
rect 21900 -8430 22540 -8360
rect 21610 -8460 22540 -8430
rect 21610 -8530 21630 -8460
rect 21700 -8530 21730 -8460
rect 21800 -8530 21830 -8460
rect 21900 -8530 22540 -8460
rect 21610 -8560 22540 -8530
rect 21610 -8630 21630 -8560
rect 21700 -8630 21730 -8560
rect 21800 -8630 21830 -8560
rect 21900 -8630 22540 -8560
rect 21610 -8650 22540 -8630
rect 22630 -9010 22950 -8980
rect 22630 -9080 22650 -9010
rect 22720 -9080 22750 -9010
rect 22820 -9080 22850 -9010
rect 22920 -9080 22950 -9010
rect 22630 -9110 22950 -9080
rect 22630 -9180 22650 -9110
rect 22720 -9180 22750 -9110
rect 22820 -9180 22850 -9110
rect 22920 -9180 22950 -9110
rect 22630 -9210 22950 -9180
rect 22630 -9280 22650 -9210
rect 22720 -9280 22750 -9210
rect 22820 -9280 22850 -9210
rect 22920 -9280 22950 -9210
rect 22630 -9300 22950 -9280
rect -270 -9660 210 -9618
rect -270 -9700 -250 -9660
rect -50 -9700 -20 -9660
rect 50 -9700 70 -9660
rect 190 -9700 210 -9660
rect -270 -9730 -240 -9700
rect -170 -9730 -130 -9700
rect -60 -9730 -20 -9700
rect 50 -9730 90 -9700
rect 160 -9730 210 -9700
rect -270 -9740 210 -9730
rect -270 -9780 -250 -9740
rect -210 -9780 -170 -9740
rect -130 -9780 -90 -9740
rect -50 -9780 -10 -9740
rect 30 -9780 70 -9740
rect 110 -9780 150 -9740
rect 190 -9780 210 -9740
rect -270 -9790 210 -9780
rect -270 -9820 -240 -9790
rect -170 -9820 -130 -9790
rect -60 -9820 -20 -9790
rect 50 -9820 90 -9790
rect 160 -9820 210 -9790
rect -270 -9860 -250 -9820
rect -50 -9860 -20 -9820
rect 50 -9860 70 -9820
rect 190 -9860 210 -9820
rect -270 -9900 210 -9860
rect 1080 -10340 2680 -9500
rect 7210 -9640 7690 -9618
rect 7210 -9660 7240 -9640
rect 7300 -9660 7340 -9640
rect 7400 -9660 7500 -9640
rect 7560 -9660 7600 -9640
rect 7660 -9660 7690 -9640
rect 7210 -9700 7230 -9660
rect 7300 -9700 7310 -9660
rect 7430 -9700 7470 -9660
rect 7590 -9700 7600 -9660
rect 7670 -9700 7690 -9660
rect 7210 -9730 7690 -9700
rect 7210 -9740 7240 -9730
rect 7300 -9740 7340 -9730
rect 7400 -9740 7500 -9730
rect 7560 -9740 7600 -9730
rect 7660 -9740 7690 -9730
rect 7210 -9780 7230 -9740
rect 7300 -9780 7310 -9740
rect 7430 -9780 7470 -9740
rect 7590 -9780 7600 -9740
rect 7670 -9780 7690 -9740
rect 7210 -9790 7240 -9780
rect 7300 -9790 7340 -9780
rect 7400 -9790 7500 -9780
rect 7560 -9790 7600 -9780
rect 7660 -9790 7690 -9780
rect 7210 -9820 7690 -9790
rect 7210 -9860 7230 -9820
rect 7300 -9860 7310 -9820
rect 7430 -9860 7470 -9820
rect 7590 -9860 7600 -9820
rect 7670 -9860 7690 -9820
rect 7210 -9880 7240 -9860
rect 7300 -9880 7340 -9860
rect 7400 -9880 7500 -9860
rect 7560 -9880 7600 -9860
rect 7660 -9880 7690 -9860
rect 7210 -9900 7690 -9880
rect 1080 -10410 1150 -10340
rect 1220 -10410 1260 -10340
rect 1330 -10410 1370 -10340
rect 1440 -10410 1480 -10340
rect 1550 -10410 1590 -10340
rect 1660 -10410 1700 -10340
rect 1770 -10410 1810 -10340
rect 1880 -10410 1920 -10340
rect 1990 -10410 2030 -10340
rect 2100 -10410 2140 -10340
rect 2210 -10410 2250 -10340
rect 2320 -10410 2360 -10340
rect 2430 -10410 2470 -10340
rect 2540 -10410 2580 -10340
rect 2650 -10410 2680 -10340
rect 1080 -10450 2680 -10410
rect 1080 -10520 1150 -10450
rect 1220 -10520 1260 -10450
rect 1330 -10520 1370 -10450
rect 1440 -10520 1480 -10450
rect 1550 -10520 1590 -10450
rect 1660 -10520 1700 -10450
rect 1770 -10520 1810 -10450
rect 1880 -10520 1920 -10450
rect 1990 -10520 2030 -10450
rect 2100 -10520 2140 -10450
rect 2210 -10520 2250 -10450
rect 2320 -10520 2360 -10450
rect 2430 -10520 2470 -10450
rect 2540 -10520 2580 -10450
rect 2650 -10520 2680 -10450
rect 1080 -10540 2680 -10520
rect 12220 -10370 13820 -9520
rect 14690 -9660 15170 -9618
rect 14690 -9700 14710 -9660
rect 14910 -9700 14940 -9660
rect 15010 -9700 15030 -9660
rect 15150 -9700 15170 -9660
rect 14690 -9730 14720 -9700
rect 14790 -9730 14830 -9700
rect 14900 -9730 14940 -9700
rect 15010 -9730 15050 -9700
rect 15120 -9730 15170 -9700
rect 14690 -9740 15170 -9730
rect 14690 -9780 14710 -9740
rect 14750 -9780 14790 -9740
rect 14830 -9780 14870 -9740
rect 14910 -9780 14950 -9740
rect 14990 -9780 15030 -9740
rect 15070 -9780 15110 -9740
rect 15150 -9780 15170 -9740
rect 14690 -9790 15170 -9780
rect 14690 -9820 14720 -9790
rect 14790 -9820 14830 -9790
rect 14900 -9820 14940 -9790
rect 15010 -9820 15050 -9790
rect 15120 -9820 15170 -9790
rect 14690 -9860 14710 -9820
rect 14910 -9860 14940 -9820
rect 15010 -9860 15030 -9820
rect 15150 -9860 15170 -9820
rect 14690 -9900 15170 -9860
rect 12220 -10440 12290 -10370
rect 12360 -10440 12400 -10370
rect 12470 -10440 12510 -10370
rect 12580 -10440 12620 -10370
rect 12690 -10440 12730 -10370
rect 12800 -10440 12840 -10370
rect 12910 -10440 12950 -10370
rect 13020 -10440 13060 -10370
rect 13130 -10440 13170 -10370
rect 13240 -10440 13280 -10370
rect 13350 -10440 13390 -10370
rect 13460 -10440 13500 -10370
rect 13570 -10440 13610 -10370
rect 13680 -10440 13720 -10370
rect 13790 -10440 13820 -10370
rect 12220 -10480 13820 -10440
rect 12220 -10550 12290 -10480
rect 12360 -10550 12400 -10480
rect 12470 -10550 12510 -10480
rect 12580 -10550 12620 -10480
rect 12690 -10550 12730 -10480
rect 12800 -10550 12840 -10480
rect 12910 -10550 12950 -10480
rect 13020 -10550 13060 -10480
rect 13130 -10550 13170 -10480
rect 13240 -10550 13280 -10480
rect 13350 -10550 13390 -10480
rect 13460 -10550 13500 -10480
rect 13570 -10550 13610 -10480
rect 13680 -10550 13720 -10480
rect 13790 -10550 13820 -10480
rect 12220 -10570 13820 -10550
rect 1510 -12300 3110 -12280
rect 1510 -12370 1540 -12300
rect 1610 -12370 1650 -12300
rect 1720 -12370 1760 -12300
rect 1830 -12370 1870 -12300
rect 1940 -12370 1980 -12300
rect 2050 -12370 2090 -12300
rect 2160 -12370 2200 -12300
rect 2270 -12370 2310 -12300
rect 2380 -12370 2420 -12300
rect 2490 -12370 2530 -12300
rect 2600 -12370 2640 -12300
rect 2710 -12370 2750 -12300
rect 2820 -12370 2860 -12300
rect 2930 -12370 2970 -12300
rect 3040 -12370 3110 -12300
rect 1510 -12410 3110 -12370
rect 1510 -12480 1540 -12410
rect 1610 -12480 1650 -12410
rect 1720 -12480 1760 -12410
rect 1830 -12480 1870 -12410
rect 1940 -12480 1980 -12410
rect 2050 -12480 2090 -12410
rect 2160 -12480 2200 -12410
rect 2270 -12480 2310 -12410
rect 2380 -12480 2420 -12410
rect 2490 -12480 2530 -12410
rect 2600 -12480 2640 -12410
rect 2710 -12480 2750 -12410
rect 2820 -12480 2860 -12410
rect 2930 -12480 2970 -12410
rect 3040 -12480 3110 -12410
rect 1510 -12550 3110 -12480
rect 11790 -12300 13390 -12280
rect 11790 -12370 11820 -12300
rect 11890 -12370 11930 -12300
rect 12000 -12370 12040 -12300
rect 12110 -12370 12150 -12300
rect 12220 -12370 12260 -12300
rect 12330 -12370 12370 -12300
rect 12440 -12370 12480 -12300
rect 12550 -12370 12590 -12300
rect 12660 -12370 12700 -12300
rect 12770 -12370 12810 -12300
rect 12880 -12370 12920 -12300
rect 12990 -12370 13030 -12300
rect 13100 -12370 13140 -12300
rect 13210 -12370 13250 -12300
rect 13320 -12370 13390 -12300
rect 11790 -12410 13390 -12370
rect 11790 -12480 11820 -12410
rect 11890 -12480 11930 -12410
rect 12000 -12480 12040 -12410
rect 12110 -12480 12150 -12410
rect 12220 -12480 12260 -12410
rect 12330 -12480 12370 -12410
rect 12440 -12480 12480 -12410
rect 12550 -12480 12590 -12410
rect 12660 -12480 12700 -12410
rect 12770 -12480 12810 -12410
rect 12880 -12480 12920 -12410
rect 12990 -12480 13030 -12410
rect 13100 -12480 13140 -12410
rect 13210 -12480 13250 -12410
rect 13320 -12480 13390 -12410
rect 11790 -12550 13390 -12480
rect 21610 -14020 22820 -13990
rect 21610 -14090 21630 -14020
rect 21700 -14090 21730 -14020
rect 21800 -14090 21830 -14020
rect 21900 -14090 22820 -14020
rect 21610 -14120 22820 -14090
rect 21610 -14190 21630 -14120
rect 21700 -14190 21730 -14120
rect 21800 -14190 21830 -14120
rect 21900 -14190 22820 -14120
rect 21610 -14220 22820 -14190
rect 21610 -14290 21630 -14220
rect 21700 -14290 21730 -14220
rect 21800 -14290 21830 -14220
rect 21900 -14290 22820 -14220
rect 21610 -14310 22820 -14290
rect 22900 -14870 23220 -14840
rect 22900 -14940 22920 -14870
rect 22990 -14940 23020 -14870
rect 23090 -14940 23120 -14870
rect 23190 -14940 23220 -14870
rect 22900 -14970 23220 -14940
rect 22900 -15040 22920 -14970
rect 22990 -15040 23020 -14970
rect 23090 -15040 23120 -14970
rect 23190 -15040 23220 -14970
rect 22900 -15070 23220 -15040
rect 22900 -15140 22920 -15070
rect 22990 -15140 23020 -15070
rect 23090 -15140 23120 -15070
rect 23190 -15140 23220 -15070
rect 22900 -15160 23220 -15140
rect 6440 -17750 6750 -17730
rect 6440 -17820 6460 -17750
rect 6530 -17820 6560 -17750
rect 6630 -17820 6660 -17750
rect 6730 -17820 6750 -17750
rect 6440 -17860 6750 -17820
rect 6440 -17930 6460 -17860
rect 6530 -17930 6560 -17860
rect 6630 -17930 6660 -17860
rect 6730 -17930 6750 -17860
rect 6440 -17970 6750 -17930
rect 6440 -18040 6460 -17970
rect 6530 -18040 6560 -17970
rect 6630 -18040 6660 -17970
rect 6730 -18040 6750 -17970
rect 6440 -18080 6750 -18040
rect 6440 -18150 6460 -18080
rect 6530 -18150 6560 -18080
rect 6630 -18150 6660 -18080
rect 6730 -18150 6750 -18080
rect 6440 -18170 6750 -18150
rect 8150 -17750 8460 -17730
rect 8150 -17820 8170 -17750
rect 8240 -17820 8270 -17750
rect 8340 -17820 8370 -17750
rect 8440 -17820 8460 -17750
rect 8150 -17860 8460 -17820
rect 8150 -17930 8170 -17860
rect 8240 -17930 8270 -17860
rect 8340 -17930 8370 -17860
rect 8440 -17930 8460 -17860
rect 8150 -17970 8460 -17930
rect 8150 -18040 8170 -17970
rect 8240 -18040 8270 -17970
rect 8340 -18040 8370 -17970
rect 8440 -18040 8460 -17970
rect 8150 -18080 8460 -18040
rect 8150 -18150 8170 -18080
rect 8240 -18150 8270 -18080
rect 8340 -18150 8370 -18080
rect 8440 -18150 8460 -18080
rect 8150 -18170 8460 -18150
rect 21610 -20100 22620 -20070
rect 21610 -20170 21630 -20100
rect 21700 -20170 21730 -20100
rect 21800 -20170 21830 -20100
rect 21900 -20170 22620 -20100
rect 21610 -20200 22620 -20170
rect 21610 -20270 21630 -20200
rect 21700 -20270 21730 -20200
rect 21800 -20270 21830 -20200
rect 21900 -20270 22620 -20200
rect 21610 -20300 22620 -20270
rect 21610 -20370 21630 -20300
rect 21700 -20370 21730 -20300
rect 21800 -20370 21830 -20300
rect 21900 -20370 22620 -20300
rect 21610 -20390 22620 -20370
rect 22680 -20730 23000 -20700
rect 22680 -20800 22700 -20730
rect 22770 -20800 22800 -20730
rect 22870 -20800 22900 -20730
rect 22970 -20800 23000 -20730
rect 22680 -20830 23000 -20800
rect 22680 -20900 22700 -20830
rect 22770 -20900 22800 -20830
rect 22870 -20900 22900 -20830
rect 22970 -20900 23000 -20830
rect 22680 -20930 23000 -20900
rect 22680 -21000 22700 -20930
rect 22770 -21000 22800 -20930
rect 22870 -21000 22900 -20930
rect 22970 -21000 23000 -20930
rect 22680 -21020 23000 -21000
rect 1550 -22660 3150 -22590
rect 1550 -22730 1620 -22660
rect 1690 -22730 1730 -22660
rect 1800 -22730 1840 -22660
rect 1910 -22730 1950 -22660
rect 2020 -22730 2060 -22660
rect 2130 -22730 2170 -22660
rect 2240 -22730 2280 -22660
rect 2350 -22730 2390 -22660
rect 2460 -22730 2500 -22660
rect 2570 -22730 2610 -22660
rect 2680 -22730 2720 -22660
rect 2790 -22730 2830 -22660
rect 2900 -22730 2940 -22660
rect 3010 -22730 3050 -22660
rect 3120 -22730 3150 -22660
rect 1550 -22770 3150 -22730
rect 1550 -22840 1620 -22770
rect 1690 -22840 1730 -22770
rect 1800 -22840 1840 -22770
rect 1910 -22840 1950 -22770
rect 2020 -22840 2060 -22770
rect 2130 -22840 2170 -22770
rect 2240 -22840 2280 -22770
rect 2350 -22840 2390 -22770
rect 2460 -22840 2500 -22770
rect 2570 -22840 2610 -22770
rect 2680 -22840 2720 -22770
rect 2790 -22840 2830 -22770
rect 2900 -22840 2940 -22770
rect 3010 -22840 3050 -22770
rect 3120 -22840 3150 -22770
rect 1550 -22860 3150 -22840
rect 11750 -22660 13350 -22590
rect 11750 -22730 11820 -22660
rect 11890 -22730 11930 -22660
rect 12000 -22730 12040 -22660
rect 12110 -22730 12150 -22660
rect 12220 -22730 12260 -22660
rect 12330 -22730 12370 -22660
rect 12440 -22730 12480 -22660
rect 12550 -22730 12590 -22660
rect 12660 -22730 12700 -22660
rect 12770 -22730 12810 -22660
rect 12880 -22730 12920 -22660
rect 12990 -22730 13030 -22660
rect 13100 -22730 13140 -22660
rect 13210 -22730 13250 -22660
rect 13320 -22730 13350 -22660
rect 11750 -22770 13350 -22730
rect 11750 -22840 11820 -22770
rect 11890 -22840 11930 -22770
rect 12000 -22840 12040 -22770
rect 12110 -22840 12150 -22770
rect 12220 -22840 12260 -22770
rect 12330 -22840 12370 -22770
rect 12440 -22840 12480 -22770
rect 12550 -22840 12590 -22770
rect 12660 -22840 12700 -22770
rect 12770 -22840 12810 -22770
rect 12880 -22840 12920 -22770
rect 12990 -22840 13030 -22770
rect 13100 -22840 13140 -22770
rect 13210 -22840 13250 -22770
rect 13320 -22840 13350 -22770
rect 11750 -22860 13350 -22840
<< via1 >>
rect 23490 7140 23560 7210
rect 23600 7140 23670 7210
rect 23710 7140 23780 7210
rect 23820 7140 23890 7210
rect 23490 7030 23560 7100
rect 23600 7030 23670 7100
rect 23710 7030 23780 7100
rect 23820 7030 23890 7100
rect 25890 7140 25960 7210
rect 26000 7140 26070 7210
rect 26110 7140 26180 7210
rect 26220 7140 26290 7210
rect 25890 7030 25960 7100
rect 26000 7030 26070 7100
rect 26110 7030 26180 7100
rect 26220 7030 26290 7100
rect 1570 6780 1640 6850
rect 1680 6780 1750 6850
rect 1790 6780 1860 6850
rect 1900 6780 1970 6850
rect 2010 6780 2080 6850
rect 2120 6780 2190 6850
rect 2230 6780 2300 6850
rect 2340 6780 2410 6850
rect 2450 6780 2520 6850
rect 2560 6780 2630 6850
rect 2670 6780 2740 6850
rect 2780 6780 2850 6850
rect 2890 6780 2960 6850
rect 3000 6780 3070 6850
rect 1570 6670 1640 6740
rect 1680 6670 1750 6740
rect 1790 6670 1860 6740
rect 1900 6670 1970 6740
rect 2010 6670 2080 6740
rect 2120 6670 2190 6740
rect 2230 6670 2300 6740
rect 2340 6670 2410 6740
rect 2450 6670 2520 6740
rect 2560 6670 2630 6740
rect 2670 6670 2740 6740
rect 2780 6670 2850 6740
rect 2890 6670 2960 6740
rect 3000 6670 3070 6740
rect 11790 6810 11860 6880
rect 11900 6810 11970 6880
rect 12010 6810 12080 6880
rect 12120 6810 12190 6880
rect 12230 6810 12300 6880
rect 12340 6810 12410 6880
rect 12450 6810 12520 6880
rect 12560 6810 12630 6880
rect 12670 6810 12740 6880
rect 12780 6810 12850 6880
rect 12890 6810 12960 6880
rect 13000 6810 13070 6880
rect 13110 6810 13180 6880
rect 13220 6810 13290 6880
rect 11790 6700 11860 6770
rect 11900 6700 11970 6770
rect 12010 6700 12080 6770
rect 12120 6700 12190 6770
rect 12230 6700 12300 6770
rect 12340 6700 12410 6770
rect 12450 6700 12520 6770
rect 12560 6700 12630 6770
rect 12670 6700 12740 6770
rect 12780 6700 12850 6770
rect 12890 6700 12960 6770
rect 13000 6700 13070 6770
rect 13110 6700 13180 6770
rect 13220 6700 13290 6770
rect 7380 6230 7440 6290
rect 7480 6230 7540 6290
rect 22780 6210 22850 6280
rect 22890 6210 22960 6280
rect 23000 6210 23070 6280
rect 23110 6210 23180 6280
rect 7380 6080 7440 6190
rect 7480 6080 7540 6190
rect 22780 6100 22850 6170
rect 22890 6100 22960 6170
rect 23000 6100 23070 6170
rect 23110 6100 23180 6170
rect 7380 5980 7440 6040
rect 7480 5980 7540 6040
rect 22780 5990 22850 6060
rect 22890 5990 22960 6060
rect 23000 5990 23070 6060
rect 23110 5990 23180 6060
rect 21820 5600 21890 5670
rect 21930 5600 22000 5670
rect 21820 5490 21890 5560
rect 21930 5490 22000 5560
rect 7410 5320 7480 5390
rect 7410 5210 7480 5280
rect 7410 5100 7480 5170
rect 7410 4990 7480 5060
rect 7410 4880 7480 4950
rect 21820 5380 21890 5450
rect 21930 5380 22000 5450
rect 21820 5270 21890 5340
rect 21930 5270 22000 5340
rect 21820 5160 21890 5230
rect 21930 5160 22000 5230
rect 21820 5050 21890 5120
rect 21930 5050 22000 5120
rect 21820 4940 21890 5010
rect 21930 4940 22000 5010
rect 21820 4830 21890 4900
rect 21930 4830 22000 4900
rect 27710 4810 27770 4870
rect 27810 4810 27870 4870
rect 27910 4810 27970 4870
rect 21820 4720 21890 4790
rect 21930 4720 22000 4790
rect 27710 4710 27770 4770
rect 27810 4710 27870 4770
rect 27910 4710 27970 4770
rect 21820 4610 21890 4680
rect 21930 4610 22000 4680
rect 27710 4610 27770 4670
rect 27810 4610 27870 4670
rect 27910 4610 27970 4670
rect -2490 4550 -2480 4580
rect -2480 4550 -2420 4580
rect -2490 4510 -2420 4550
rect -2490 4430 -2420 4470
rect -2490 4400 -2480 4430
rect -2480 4400 -2420 4430
rect -2490 4350 -2420 4360
rect -2490 4310 -2480 4350
rect -2480 4310 -2420 4350
rect -2490 4290 -2420 4310
rect -2490 4230 -2480 4250
rect -2480 4230 -2420 4250
rect -2490 4190 -2420 4230
rect -2490 4180 -2480 4190
rect -2480 4180 -2420 4190
rect 17200 4550 17260 4580
rect 17260 4550 17270 4580
rect 17200 4510 17270 4550
rect 17200 4430 17270 4470
rect 17200 4400 17260 4430
rect 17260 4400 17270 4430
rect 17200 4350 17270 4360
rect 17200 4310 17260 4350
rect 17260 4310 17270 4350
rect 17200 4290 17270 4310
rect 17200 4230 17260 4250
rect 17260 4230 17270 4250
rect 17200 4190 17270 4230
rect 17200 4180 17260 4190
rect 17260 4180 17270 4190
rect 21820 4500 21890 4570
rect 21930 4500 22000 4570
rect 27710 4510 27770 4570
rect 27810 4510 27870 4570
rect 27910 4510 27970 4570
rect 27710 4410 27770 4470
rect 27810 4410 27870 4470
rect 27910 4410 27970 4470
rect 27710 4310 27770 4370
rect 27810 4310 27870 4370
rect 27910 4310 27970 4370
rect 27710 4210 27770 4270
rect 27810 4210 27870 4270
rect 27910 4210 27970 4270
rect 27710 4110 27770 4170
rect 27810 4110 27870 4170
rect 27910 4110 27970 4170
rect 27710 4010 27770 4070
rect 27810 4010 27870 4070
rect 27910 4010 27970 4070
rect 24720 3290 24790 3360
rect 24830 3290 24900 3360
rect 24940 3290 25010 3360
rect 7050 3220 7110 3280
rect 7150 3220 7210 3280
rect 7250 3220 7310 3280
rect 7590 3220 7650 3280
rect 7690 3220 7750 3280
rect 7790 3220 7850 3280
rect 24720 3180 24790 3250
rect 24830 3180 24900 3250
rect 24940 3180 25010 3250
rect 7050 3120 7110 3180
rect 7150 3120 7210 3180
rect 7250 3120 7310 3180
rect 7590 3120 7650 3180
rect 7690 3120 7750 3180
rect 7790 3120 7850 3180
rect 7050 3020 7110 3080
rect 7150 3020 7210 3080
rect 7250 3020 7310 3080
rect 7590 3020 7650 3080
rect 7690 3020 7750 3080
rect 7790 3020 7850 3080
rect 24720 3070 24790 3140
rect 24830 3070 24900 3140
rect 24940 3070 25010 3140
rect 4770 2830 4830 2890
rect 4870 2830 4930 2890
rect 4970 2830 5030 2890
rect 9870 2830 9930 2890
rect 9970 2830 10030 2890
rect 10070 2830 10130 2890
rect 4770 2730 4830 2790
rect 4870 2730 4930 2790
rect 4970 2730 5030 2790
rect 9870 2730 9930 2790
rect 9970 2730 10030 2790
rect 10070 2730 10130 2790
rect 4770 2630 4830 2690
rect 4870 2630 4930 2690
rect 4970 2630 5030 2690
rect 9870 2630 9930 2690
rect 9970 2630 10030 2690
rect 10070 2630 10130 2690
rect 22470 2530 22540 2600
rect 22580 2530 22650 2600
rect 22690 2530 22760 2600
rect 22800 2530 22870 2600
rect 22470 2420 22540 2490
rect 22580 2420 22650 2490
rect 22690 2420 22760 2490
rect 22800 2420 22870 2490
rect 26950 2530 27020 2600
rect 27060 2530 27130 2600
rect 27170 2530 27240 2600
rect 27280 2530 27350 2600
rect 26950 2420 27020 2490
rect 27060 2420 27130 2490
rect 27170 2420 27240 2490
rect 27280 2420 27350 2490
rect 20 1090 90 1160
rect 130 1090 200 1160
rect 230 1090 300 1160
rect 20 980 90 1050
rect 130 980 200 1050
rect 230 980 300 1050
rect 20 870 90 940
rect 130 870 200 940
rect 230 870 300 940
rect 14600 1090 14670 1160
rect 14700 1090 14770 1160
rect 14810 1090 14880 1160
rect 14600 980 14670 1050
rect 14700 980 14770 1050
rect 14810 980 14880 1050
rect 14600 870 14670 940
rect 14700 870 14770 940
rect 14810 870 14880 940
rect 23490 850 23560 920
rect 23600 850 23670 920
rect 23710 850 23780 920
rect 23820 850 23890 920
rect 23490 740 23560 810
rect 23600 740 23670 810
rect 23710 740 23780 810
rect 23820 740 23890 810
rect 25890 850 25960 920
rect 26000 850 26070 920
rect 26110 850 26180 920
rect 26220 850 26290 920
rect 25890 740 25960 810
rect 26000 740 26070 810
rect 26110 740 26180 810
rect 26220 740 26290 810
rect -300 -180 -270 -140
rect -270 -180 -230 -140
rect -190 -180 -150 -140
rect -150 -180 -120 -140
rect -80 -180 -70 -140
rect -70 -180 -30 -140
rect -30 -180 -10 -140
rect 30 -180 50 -140
rect 50 -180 90 -140
rect 90 -180 100 -140
rect -300 -210 -230 -180
rect -190 -210 -120 -180
rect -80 -210 -10 -180
rect 30 -210 100 -180
rect -300 -300 -230 -270
rect -190 -300 -120 -270
rect -80 -300 -10 -270
rect 30 -300 100 -270
rect -300 -340 -270 -300
rect -270 -340 -230 -300
rect -190 -340 -150 -300
rect -150 -340 -120 -300
rect -80 -340 -70 -300
rect -70 -340 -30 -300
rect -30 -340 -10 -300
rect 30 -340 50 -300
rect 50 -340 90 -300
rect 90 -340 100 -300
rect 7180 -140 7240 -120
rect 7280 -140 7340 -120
rect 7440 -140 7500 -120
rect 7540 -140 7600 -120
rect 7180 -180 7210 -140
rect 7210 -180 7240 -140
rect 7280 -180 7290 -140
rect 7290 -180 7330 -140
rect 7330 -180 7340 -140
rect 7440 -180 7450 -140
rect 7450 -180 7490 -140
rect 7490 -180 7500 -140
rect 7540 -180 7570 -140
rect 7570 -180 7600 -140
rect 7180 -220 7240 -210
rect 7280 -220 7340 -210
rect 7440 -220 7500 -210
rect 7540 -220 7600 -210
rect 7180 -260 7210 -220
rect 7210 -260 7240 -220
rect 7280 -260 7290 -220
rect 7290 -260 7330 -220
rect 7330 -260 7340 -220
rect 7440 -260 7450 -220
rect 7450 -260 7490 -220
rect 7490 -260 7500 -220
rect 7540 -260 7570 -220
rect 7570 -260 7600 -220
rect 7180 -270 7240 -260
rect 7280 -270 7340 -260
rect 7440 -270 7500 -260
rect 7540 -270 7600 -260
rect 7180 -340 7210 -300
rect 7210 -340 7240 -300
rect 7280 -340 7290 -300
rect 7290 -340 7330 -300
rect 7330 -340 7340 -300
rect 7440 -340 7450 -300
rect 7450 -340 7490 -300
rect 7490 -340 7500 -300
rect 7540 -340 7570 -300
rect 7570 -340 7600 -300
rect 7180 -360 7240 -340
rect 7280 -360 7340 -340
rect 7440 -360 7500 -340
rect 7540 -360 7600 -340
rect 1150 -860 1220 -790
rect 1260 -860 1330 -790
rect 1370 -860 1440 -790
rect 1480 -860 1550 -790
rect 1590 -860 1660 -790
rect 1700 -860 1770 -790
rect 1810 -860 1880 -790
rect 1920 -860 1990 -790
rect 2030 -860 2100 -790
rect 2140 -860 2210 -790
rect 2250 -860 2320 -790
rect 2360 -860 2430 -790
rect 2470 -860 2540 -790
rect 2580 -860 2650 -790
rect 1150 -970 1220 -900
rect 1260 -970 1330 -900
rect 1370 -970 1440 -900
rect 1480 -970 1550 -900
rect 1590 -970 1660 -900
rect 1700 -970 1770 -900
rect 1810 -970 1880 -900
rect 1920 -970 1990 -900
rect 2030 -970 2100 -900
rect 2140 -970 2210 -900
rect 2250 -970 2320 -900
rect 2360 -970 2430 -900
rect 2470 -970 2540 -900
rect 2580 -970 2650 -900
rect 22780 -90 22850 -20
rect 22890 -90 22960 -20
rect 23000 -90 23070 -20
rect 23110 -90 23180 -20
rect 14660 -180 14690 -140
rect 14690 -180 14730 -140
rect 14770 -180 14810 -140
rect 14810 -180 14840 -140
rect 14880 -180 14890 -140
rect 14890 -180 14930 -140
rect 14930 -180 14950 -140
rect 14990 -180 15010 -140
rect 15010 -180 15050 -140
rect 15050 -180 15060 -140
rect 14660 -210 14730 -180
rect 14770 -210 14840 -180
rect 14880 -210 14950 -180
rect 14990 -210 15060 -180
rect 22780 -200 22850 -130
rect 22890 -200 22960 -130
rect 23000 -200 23070 -130
rect 23110 -200 23180 -130
rect 14660 -300 14730 -270
rect 14770 -300 14840 -270
rect 14880 -300 14950 -270
rect 14990 -300 15060 -270
rect 14660 -340 14690 -300
rect 14690 -340 14730 -300
rect 14770 -340 14810 -300
rect 14810 -340 14840 -300
rect 14880 -340 14890 -300
rect 14890 -340 14930 -300
rect 14930 -340 14950 -300
rect 14990 -340 15010 -300
rect 15010 -340 15050 -300
rect 15050 -340 15060 -300
rect 22780 -310 22850 -240
rect 22890 -310 22960 -240
rect 23000 -310 23070 -240
rect 23110 -310 23180 -240
rect 12250 -860 12320 -790
rect 12360 -860 12430 -790
rect 12470 -860 12540 -790
rect 12580 -860 12650 -790
rect 12690 -860 12760 -790
rect 12800 -860 12870 -790
rect 12910 -860 12980 -790
rect 13020 -860 13090 -790
rect 13130 -860 13200 -790
rect 13240 -860 13310 -790
rect 13350 -860 13420 -790
rect 13460 -860 13530 -790
rect 13570 -860 13640 -790
rect 13680 -860 13750 -790
rect 12250 -970 12320 -900
rect 12360 -970 12430 -900
rect 12470 -970 12540 -900
rect 12580 -970 12650 -900
rect 12690 -970 12760 -900
rect 12800 -970 12870 -900
rect 12910 -970 12980 -900
rect 13020 -970 13090 -900
rect 13130 -970 13200 -900
rect 13240 -970 13310 -900
rect 13350 -970 13420 -900
rect 13460 -970 13530 -900
rect 13570 -970 13640 -900
rect 13680 -970 13750 -900
rect 21820 -920 21890 -850
rect 21930 -920 22000 -850
rect 21820 -1030 21890 -960
rect 21930 -1030 22000 -960
rect 21820 -1140 21890 -1070
rect 21930 -1140 22000 -1070
rect 21820 -1250 21890 -1180
rect 21930 -1250 22000 -1180
rect 21820 -1360 21890 -1290
rect 21930 -1360 22000 -1290
rect 21820 -1470 21890 -1400
rect 21930 -1470 22000 -1400
rect 27710 -1490 27770 -1430
rect 27810 -1490 27870 -1430
rect 27910 -1490 27970 -1430
rect 21820 -1580 21890 -1510
rect 21930 -1580 22000 -1510
rect 27710 -1590 27770 -1530
rect 27810 -1590 27870 -1530
rect 27910 -1590 27970 -1530
rect 21820 -1690 21890 -1620
rect 21930 -1690 22000 -1620
rect 27710 -1690 27770 -1630
rect 27810 -1690 27870 -1630
rect 27910 -1690 27970 -1630
rect 21820 -1800 21890 -1730
rect 21930 -1800 22000 -1730
rect 27710 -1790 27770 -1730
rect 27810 -1790 27870 -1730
rect 27910 -1790 27970 -1730
rect 21820 -1910 21890 -1840
rect 21930 -1910 22000 -1840
rect 27710 -1890 27770 -1830
rect 27810 -1890 27870 -1830
rect 27910 -1890 27970 -1830
rect 21820 -2020 21890 -1950
rect 21930 -2020 22000 -1950
rect 27710 -1990 27770 -1930
rect 27810 -1990 27870 -1930
rect 27910 -1990 27970 -1930
rect 27710 -2090 27770 -2030
rect 27810 -2090 27870 -2030
rect 27910 -2090 27970 -2030
rect 27710 -2190 27770 -2130
rect 27810 -2190 27870 -2130
rect 27910 -2190 27970 -2130
rect 27710 -2290 27770 -2230
rect 27810 -2290 27870 -2230
rect 27910 -2290 27970 -2230
rect 1570 -2850 1640 -2780
rect 1680 -2850 1750 -2780
rect 1790 -2850 1860 -2780
rect 1900 -2850 1970 -2780
rect 2010 -2850 2080 -2780
rect 2120 -2850 2190 -2780
rect 2230 -2850 2300 -2780
rect 2340 -2850 2410 -2780
rect 2450 -2850 2520 -2780
rect 2560 -2850 2630 -2780
rect 2670 -2850 2740 -2780
rect 2780 -2850 2850 -2780
rect 2890 -2850 2960 -2780
rect 3000 -2850 3070 -2780
rect 1570 -2960 1640 -2890
rect 1680 -2960 1750 -2890
rect 1790 -2960 1860 -2890
rect 1900 -2960 1970 -2890
rect 2010 -2960 2080 -2890
rect 2120 -2960 2190 -2890
rect 2230 -2960 2300 -2890
rect 2340 -2960 2410 -2890
rect 2450 -2960 2520 -2890
rect 2560 -2960 2630 -2890
rect 2670 -2960 2740 -2890
rect 2780 -2960 2850 -2890
rect 2890 -2960 2960 -2890
rect 3000 -2960 3070 -2890
rect 11790 -2850 11860 -2780
rect 11900 -2850 11970 -2780
rect 12010 -2850 12080 -2780
rect 12120 -2850 12190 -2780
rect 12230 -2850 12300 -2780
rect 12340 -2850 12410 -2780
rect 12450 -2850 12520 -2780
rect 12560 -2850 12630 -2780
rect 12670 -2850 12740 -2780
rect 12780 -2850 12850 -2780
rect 12890 -2850 12960 -2780
rect 13000 -2850 13070 -2780
rect 13110 -2850 13180 -2780
rect 13220 -2850 13290 -2780
rect 11790 -2960 11860 -2890
rect 11900 -2960 11970 -2890
rect 12010 -2960 12080 -2890
rect 12120 -2960 12190 -2890
rect 12230 -2960 12300 -2890
rect 12340 -2960 12410 -2890
rect 12450 -2960 12520 -2890
rect 12560 -2960 12630 -2890
rect 12670 -2960 12740 -2890
rect 12780 -2960 12850 -2890
rect 12890 -2960 12960 -2890
rect 13000 -2960 13070 -2890
rect 13110 -2960 13180 -2890
rect 13220 -2960 13290 -2890
rect 24740 -3120 24810 -3050
rect 24850 -3120 24920 -3050
rect 24960 -3120 25030 -3050
rect 24740 -3230 24810 -3160
rect 24850 -3230 24920 -3160
rect 24960 -3230 25030 -3160
rect 24740 -3340 24810 -3270
rect 24850 -3340 24920 -3270
rect 24960 -3340 25030 -3270
rect 7380 -3400 7440 -3340
rect 7480 -3400 7540 -3340
rect 7380 -3550 7440 -3440
rect 7480 -3550 7540 -3440
rect 7380 -3650 7440 -3590
rect 7480 -3650 7540 -3590
rect 22470 -3760 22540 -3690
rect 22580 -3760 22650 -3690
rect 22690 -3760 22760 -3690
rect 22800 -3760 22870 -3690
rect 7310 -3950 7380 -3880
rect 7420 -3950 7490 -3880
rect 7530 -3950 7600 -3880
rect 22470 -3870 22540 -3800
rect 22580 -3870 22650 -3800
rect 22690 -3870 22760 -3800
rect 22800 -3870 22870 -3800
rect 26950 -3760 27020 -3690
rect 27060 -3760 27130 -3690
rect 27170 -3760 27240 -3690
rect 27280 -3760 27350 -3690
rect 26950 -3870 27020 -3800
rect 27060 -3870 27130 -3800
rect 27170 -3870 27240 -3800
rect 27280 -3870 27350 -3800
rect 7310 -4060 7380 -3990
rect 7420 -4060 7490 -3990
rect 7530 -4060 7600 -3990
rect 7310 -4170 7380 -4100
rect 7420 -4170 7490 -4100
rect 7530 -4170 7600 -4100
rect -1330 -4352 -1290 -4350
rect -1290 -4352 -1260 -4350
rect -1220 -4352 -1210 -4350
rect -1210 -4352 -1170 -4350
rect -1170 -4352 -1150 -4350
rect -1110 -4352 -1090 -4350
rect -1090 -4352 -1050 -4350
rect -1050 -4352 -1040 -4350
rect -1000 -4352 -970 -4350
rect -970 -4352 -930 -4350
rect -1330 -4392 -1260 -4352
rect -1220 -4392 -1150 -4352
rect -1110 -4392 -1040 -4352
rect -1000 -4392 -930 -4352
rect -1330 -4420 -1290 -4392
rect -1290 -4420 -1260 -4392
rect -1220 -4420 -1210 -4392
rect -1210 -4420 -1170 -4392
rect -1170 -4420 -1150 -4392
rect -1110 -4420 -1090 -4392
rect -1090 -4420 -1050 -4392
rect -1050 -4420 -1040 -4392
rect -1000 -4420 -970 -4392
rect -970 -4420 -930 -4392
rect -1330 -4472 -1260 -4460
rect -1220 -4472 -1150 -4460
rect -1110 -4472 -1040 -4460
rect -1000 -4472 -930 -4460
rect -1330 -4512 -1290 -4472
rect -1290 -4512 -1260 -4472
rect -1220 -4512 -1210 -4472
rect -1210 -4512 -1170 -4472
rect -1170 -4512 -1150 -4472
rect -1110 -4512 -1090 -4472
rect -1090 -4512 -1050 -4472
rect -1050 -4512 -1040 -4472
rect -1000 -4512 -970 -4472
rect -970 -4512 -930 -4472
rect -1330 -4530 -1260 -4512
rect -1220 -4530 -1150 -4512
rect -1110 -4530 -1040 -4512
rect -1000 -4530 -930 -4512
rect -560 -4312 -490 -4290
rect -450 -4312 -380 -4290
rect -340 -4312 -270 -4290
rect -230 -4312 -160 -4290
rect -560 -4352 -530 -4312
rect -530 -4352 -490 -4312
rect -450 -4352 -410 -4312
rect -410 -4352 -380 -4312
rect -340 -4352 -330 -4312
rect -330 -4352 -290 -4312
rect -290 -4352 -270 -4312
rect -230 -4352 -210 -4312
rect -210 -4352 -170 -4312
rect -170 -4352 -160 -4312
rect -560 -4360 -490 -4352
rect -450 -4360 -380 -4352
rect -340 -4360 -270 -4352
rect -230 -4360 -160 -4352
rect -560 -4432 -530 -4400
rect -530 -4432 -490 -4400
rect -450 -4432 -410 -4400
rect -410 -4432 -380 -4400
rect -340 -4432 -330 -4400
rect -330 -4432 -290 -4400
rect -290 -4432 -270 -4400
rect -230 -4432 -210 -4400
rect -210 -4432 -170 -4400
rect -170 -4432 -160 -4400
rect -560 -4470 -490 -4432
rect -450 -4470 -380 -4432
rect -340 -4470 -270 -4432
rect -230 -4470 -160 -4432
rect 14940 -4312 15010 -4290
rect 15050 -4312 15120 -4290
rect 15160 -4312 15230 -4290
rect 15270 -4312 15340 -4290
rect 14940 -4352 14950 -4312
rect 14950 -4352 14990 -4312
rect 14990 -4352 15010 -4312
rect 15050 -4352 15070 -4312
rect 15070 -4352 15110 -4312
rect 15110 -4352 15120 -4312
rect 15160 -4352 15190 -4312
rect 15190 -4352 15230 -4312
rect 15270 -4352 15310 -4312
rect 15310 -4352 15340 -4312
rect 14940 -4360 15010 -4352
rect 15050 -4360 15120 -4352
rect 15160 -4360 15230 -4352
rect 15270 -4360 15340 -4352
rect 14940 -4432 14950 -4400
rect 14950 -4432 14990 -4400
rect 14990 -4432 15010 -4400
rect 15050 -4432 15070 -4400
rect 15070 -4432 15110 -4400
rect 15110 -4432 15120 -4400
rect 15160 -4432 15190 -4400
rect 15190 -4432 15230 -4400
rect 15270 -4432 15310 -4400
rect 15310 -4432 15340 -4400
rect 14940 -4470 15010 -4432
rect 15050 -4470 15120 -4432
rect 15160 -4470 15230 -4432
rect 15270 -4470 15340 -4432
rect 15710 -4352 15750 -4350
rect 15750 -4352 15780 -4350
rect 15820 -4352 15830 -4350
rect 15830 -4352 15870 -4350
rect 15870 -4352 15890 -4350
rect 15930 -4352 15950 -4350
rect 15950 -4352 15990 -4350
rect 15990 -4352 16000 -4350
rect 16040 -4352 16070 -4350
rect 16070 -4352 16110 -4350
rect 15710 -4392 15780 -4352
rect 15820 -4392 15890 -4352
rect 15930 -4392 16000 -4352
rect 16040 -4392 16110 -4352
rect 15710 -4420 15750 -4392
rect 15750 -4420 15780 -4392
rect 15820 -4420 15830 -4392
rect 15830 -4420 15870 -4392
rect 15870 -4420 15890 -4392
rect 15930 -4420 15950 -4392
rect 15950 -4420 15990 -4392
rect 15990 -4420 16000 -4392
rect 16040 -4420 16070 -4392
rect 16070 -4420 16110 -4392
rect 15710 -4472 15780 -4460
rect 15820 -4472 15890 -4460
rect 15930 -4472 16000 -4460
rect 16040 -4472 16110 -4460
rect 15710 -4512 15750 -4472
rect 15750 -4512 15780 -4472
rect 15820 -4512 15830 -4472
rect 15830 -4512 15870 -4472
rect 15870 -4512 15890 -4472
rect 15930 -4512 15950 -4472
rect 15950 -4512 15990 -4472
rect 15990 -4512 16000 -4472
rect 16040 -4512 16070 -4472
rect 16070 -4512 16110 -4472
rect 15710 -4530 15780 -4512
rect 15820 -4530 15890 -4512
rect 15930 -4530 16000 -4512
rect 16040 -4530 16110 -4512
rect -1710 -6530 -1700 -6520
rect -1700 -6530 -1640 -6520
rect -1710 -6570 -1640 -6530
rect -1710 -6590 -1700 -6570
rect -1700 -6590 -1640 -6570
rect 7050 -6520 7110 -6460
rect 7150 -6520 7210 -6460
rect 7250 -6520 7310 -6460
rect 7590 -6520 7650 -6460
rect 7690 -6520 7750 -6460
rect 7790 -6520 7850 -6460
rect 7050 -6620 7110 -6560
rect 7150 -6620 7210 -6560
rect 7250 -6620 7310 -6560
rect 7590 -6620 7650 -6560
rect 7690 -6620 7750 -6560
rect 7790 -6620 7850 -6560
rect -1710 -6650 -1640 -6630
rect -1710 -6690 -1700 -6650
rect -1700 -6690 -1640 -6650
rect -1710 -6700 -1640 -6690
rect 4770 -6730 4830 -6670
rect 4870 -6730 4930 -6670
rect 4970 -6730 5030 -6670
rect 7050 -6720 7110 -6660
rect 7150 -6720 7210 -6660
rect 7250 -6720 7310 -6660
rect 7590 -6720 7650 -6660
rect 7690 -6720 7750 -6660
rect 7790 -6720 7850 -6660
rect 16420 -6530 16480 -6520
rect 16480 -6530 16490 -6520
rect 16420 -6570 16490 -6530
rect 16420 -6590 16480 -6570
rect 16480 -6590 16490 -6570
rect -1710 -6770 -1700 -6740
rect -1700 -6770 -1640 -6740
rect -1710 -6810 -1640 -6770
rect -1710 -6890 -1640 -6850
rect -1710 -6920 -1700 -6890
rect -1700 -6920 -1640 -6890
rect 9870 -6730 9930 -6670
rect 9970 -6730 10030 -6670
rect 10070 -6730 10130 -6670
rect 16420 -6650 16490 -6630
rect 16420 -6690 16480 -6650
rect 16480 -6690 16490 -6650
rect 16420 -6700 16490 -6690
rect 4770 -6830 4830 -6770
rect 4870 -6830 4930 -6770
rect 4970 -6830 5030 -6770
rect 7050 -6820 7110 -6760
rect 7150 -6820 7210 -6760
rect 7250 -6820 7310 -6760
rect 7590 -6820 7650 -6760
rect 7690 -6820 7750 -6760
rect 7790 -6820 7850 -6760
rect 9870 -6830 9930 -6770
rect 9970 -6830 10030 -6770
rect 10070 -6830 10130 -6770
rect 4770 -6930 4830 -6870
rect 4870 -6930 4930 -6870
rect 4970 -6930 5030 -6870
rect 9870 -6930 9930 -6870
rect 9970 -6930 10030 -6870
rect 10070 -6930 10130 -6870
rect 16420 -6770 16480 -6740
rect 16480 -6770 16490 -6740
rect 16420 -6810 16490 -6770
rect 16420 -6890 16490 -6850
rect 16420 -6920 16480 -6890
rect 16480 -6920 16490 -6890
rect 20 -8210 90 -8140
rect 130 -8210 200 -8140
rect 230 -8210 300 -8140
rect 20 -8320 90 -8250
rect 130 -8320 200 -8250
rect 230 -8320 300 -8250
rect 20 -8430 90 -8360
rect 130 -8430 200 -8360
rect 230 -8430 300 -8360
rect 14600 -8300 14670 -8230
rect 14700 -8300 14770 -8230
rect 14810 -8300 14880 -8230
rect 14600 -8410 14670 -8340
rect 14700 -8410 14770 -8340
rect 14810 -8410 14880 -8340
rect 14600 -8520 14670 -8450
rect 14700 -8520 14770 -8450
rect 14810 -8520 14880 -8450
rect 21630 -8430 21700 -8360
rect 21730 -8430 21800 -8360
rect 21830 -8430 21900 -8360
rect 21630 -8530 21700 -8460
rect 21730 -8530 21800 -8460
rect 21830 -8530 21900 -8460
rect 21630 -8630 21700 -8560
rect 21730 -8630 21800 -8560
rect 21830 -8630 21900 -8560
rect 22650 -9080 22720 -9010
rect 22750 -9080 22820 -9010
rect 22850 -9080 22920 -9010
rect 22650 -9180 22720 -9110
rect 22750 -9180 22820 -9110
rect 22850 -9180 22920 -9110
rect 22650 -9280 22720 -9210
rect 22750 -9280 22820 -9210
rect 22850 -9280 22920 -9210
rect -240 -9700 -210 -9660
rect -210 -9700 -170 -9660
rect -130 -9700 -90 -9660
rect -90 -9700 -60 -9660
rect -20 -9700 -10 -9660
rect -10 -9700 30 -9660
rect 30 -9700 50 -9660
rect 90 -9700 110 -9660
rect 110 -9700 150 -9660
rect 150 -9700 160 -9660
rect -240 -9730 -170 -9700
rect -130 -9730 -60 -9700
rect -20 -9730 50 -9700
rect 90 -9730 160 -9700
rect -240 -9820 -170 -9790
rect -130 -9820 -60 -9790
rect -20 -9820 50 -9790
rect 90 -9820 160 -9790
rect -240 -9860 -210 -9820
rect -210 -9860 -170 -9820
rect -130 -9860 -90 -9820
rect -90 -9860 -60 -9820
rect -20 -9860 -10 -9820
rect -10 -9860 30 -9820
rect 30 -9860 50 -9820
rect 90 -9860 110 -9820
rect 110 -9860 150 -9820
rect 150 -9860 160 -9820
rect 7240 -9660 7300 -9640
rect 7340 -9660 7400 -9640
rect 7500 -9660 7560 -9640
rect 7600 -9660 7660 -9640
rect 7240 -9700 7270 -9660
rect 7270 -9700 7300 -9660
rect 7340 -9700 7350 -9660
rect 7350 -9700 7390 -9660
rect 7390 -9700 7400 -9660
rect 7500 -9700 7510 -9660
rect 7510 -9700 7550 -9660
rect 7550 -9700 7560 -9660
rect 7600 -9700 7630 -9660
rect 7630 -9700 7660 -9660
rect 7240 -9740 7300 -9730
rect 7340 -9740 7400 -9730
rect 7500 -9740 7560 -9730
rect 7600 -9740 7660 -9730
rect 7240 -9780 7270 -9740
rect 7270 -9780 7300 -9740
rect 7340 -9780 7350 -9740
rect 7350 -9780 7390 -9740
rect 7390 -9780 7400 -9740
rect 7500 -9780 7510 -9740
rect 7510 -9780 7550 -9740
rect 7550 -9780 7560 -9740
rect 7600 -9780 7630 -9740
rect 7630 -9780 7660 -9740
rect 7240 -9790 7300 -9780
rect 7340 -9790 7400 -9780
rect 7500 -9790 7560 -9780
rect 7600 -9790 7660 -9780
rect 7240 -9860 7270 -9820
rect 7270 -9860 7300 -9820
rect 7340 -9860 7350 -9820
rect 7350 -9860 7390 -9820
rect 7390 -9860 7400 -9820
rect 7500 -9860 7510 -9820
rect 7510 -9860 7550 -9820
rect 7550 -9860 7560 -9820
rect 7600 -9860 7630 -9820
rect 7630 -9860 7660 -9820
rect 7240 -9880 7300 -9860
rect 7340 -9880 7400 -9860
rect 7500 -9880 7560 -9860
rect 7600 -9880 7660 -9860
rect 1150 -10410 1220 -10340
rect 1260 -10410 1330 -10340
rect 1370 -10410 1440 -10340
rect 1480 -10410 1550 -10340
rect 1590 -10410 1660 -10340
rect 1700 -10410 1770 -10340
rect 1810 -10410 1880 -10340
rect 1920 -10410 1990 -10340
rect 2030 -10410 2100 -10340
rect 2140 -10410 2210 -10340
rect 2250 -10410 2320 -10340
rect 2360 -10410 2430 -10340
rect 2470 -10410 2540 -10340
rect 2580 -10410 2650 -10340
rect 1150 -10520 1220 -10450
rect 1260 -10520 1330 -10450
rect 1370 -10520 1440 -10450
rect 1480 -10520 1550 -10450
rect 1590 -10520 1660 -10450
rect 1700 -10520 1770 -10450
rect 1810 -10520 1880 -10450
rect 1920 -10520 1990 -10450
rect 2030 -10520 2100 -10450
rect 2140 -10520 2210 -10450
rect 2250 -10520 2320 -10450
rect 2360 -10520 2430 -10450
rect 2470 -10520 2540 -10450
rect 2580 -10520 2650 -10450
rect 14720 -9700 14750 -9660
rect 14750 -9700 14790 -9660
rect 14830 -9700 14870 -9660
rect 14870 -9700 14900 -9660
rect 14940 -9700 14950 -9660
rect 14950 -9700 14990 -9660
rect 14990 -9700 15010 -9660
rect 15050 -9700 15070 -9660
rect 15070 -9700 15110 -9660
rect 15110 -9700 15120 -9660
rect 14720 -9730 14790 -9700
rect 14830 -9730 14900 -9700
rect 14940 -9730 15010 -9700
rect 15050 -9730 15120 -9700
rect 14720 -9820 14790 -9790
rect 14830 -9820 14900 -9790
rect 14940 -9820 15010 -9790
rect 15050 -9820 15120 -9790
rect 14720 -9860 14750 -9820
rect 14750 -9860 14790 -9820
rect 14830 -9860 14870 -9820
rect 14870 -9860 14900 -9820
rect 14940 -9860 14950 -9820
rect 14950 -9860 14990 -9820
rect 14990 -9860 15010 -9820
rect 15050 -9860 15070 -9820
rect 15070 -9860 15110 -9820
rect 15110 -9860 15120 -9820
rect 12290 -10440 12360 -10370
rect 12400 -10440 12470 -10370
rect 12510 -10440 12580 -10370
rect 12620 -10440 12690 -10370
rect 12730 -10440 12800 -10370
rect 12840 -10440 12910 -10370
rect 12950 -10440 13020 -10370
rect 13060 -10440 13130 -10370
rect 13170 -10440 13240 -10370
rect 13280 -10440 13350 -10370
rect 13390 -10440 13460 -10370
rect 13500 -10440 13570 -10370
rect 13610 -10440 13680 -10370
rect 13720 -10440 13790 -10370
rect 12290 -10550 12360 -10480
rect 12400 -10550 12470 -10480
rect 12510 -10550 12580 -10480
rect 12620 -10550 12690 -10480
rect 12730 -10550 12800 -10480
rect 12840 -10550 12910 -10480
rect 12950 -10550 13020 -10480
rect 13060 -10550 13130 -10480
rect 13170 -10550 13240 -10480
rect 13280 -10550 13350 -10480
rect 13390 -10550 13460 -10480
rect 13500 -10550 13570 -10480
rect 13610 -10550 13680 -10480
rect 13720 -10550 13790 -10480
rect 1540 -12370 1610 -12300
rect 1650 -12370 1720 -12300
rect 1760 -12370 1830 -12300
rect 1870 -12370 1940 -12300
rect 1980 -12370 2050 -12300
rect 2090 -12370 2160 -12300
rect 2200 -12370 2270 -12300
rect 2310 -12370 2380 -12300
rect 2420 -12370 2490 -12300
rect 2530 -12370 2600 -12300
rect 2640 -12370 2710 -12300
rect 2750 -12370 2820 -12300
rect 2860 -12370 2930 -12300
rect 2970 -12370 3040 -12300
rect 1540 -12480 1610 -12410
rect 1650 -12480 1720 -12410
rect 1760 -12480 1830 -12410
rect 1870 -12480 1940 -12410
rect 1980 -12480 2050 -12410
rect 2090 -12480 2160 -12410
rect 2200 -12480 2270 -12410
rect 2310 -12480 2380 -12410
rect 2420 -12480 2490 -12410
rect 2530 -12480 2600 -12410
rect 2640 -12480 2710 -12410
rect 2750 -12480 2820 -12410
rect 2860 -12480 2930 -12410
rect 2970 -12480 3040 -12410
rect 11820 -12370 11890 -12300
rect 11930 -12370 12000 -12300
rect 12040 -12370 12110 -12300
rect 12150 -12370 12220 -12300
rect 12260 -12370 12330 -12300
rect 12370 -12370 12440 -12300
rect 12480 -12370 12550 -12300
rect 12590 -12370 12660 -12300
rect 12700 -12370 12770 -12300
rect 12810 -12370 12880 -12300
rect 12920 -12370 12990 -12300
rect 13030 -12370 13100 -12300
rect 13140 -12370 13210 -12300
rect 13250 -12370 13320 -12300
rect 11820 -12480 11890 -12410
rect 11930 -12480 12000 -12410
rect 12040 -12480 12110 -12410
rect 12150 -12480 12220 -12410
rect 12260 -12480 12330 -12410
rect 12370 -12480 12440 -12410
rect 12480 -12480 12550 -12410
rect 12590 -12480 12660 -12410
rect 12700 -12480 12770 -12410
rect 12810 -12480 12880 -12410
rect 12920 -12480 12990 -12410
rect 13030 -12480 13100 -12410
rect 13140 -12480 13210 -12410
rect 13250 -12480 13320 -12410
rect 6310 -13310 6370 -13250
rect 6410 -13310 6470 -13250
rect 6510 -13310 6570 -13250
rect 8330 -13310 8390 -13250
rect 8430 -13310 8490 -13250
rect 8530 -13310 8590 -13250
rect 6310 -13400 6370 -13340
rect 6410 -13400 6470 -13340
rect 6510 -13400 6570 -13340
rect 8330 -13400 8390 -13340
rect 8430 -13400 8490 -13340
rect 8530 -13400 8590 -13340
rect 6310 -13490 6370 -13430
rect 6410 -13490 6470 -13430
rect 6510 -13490 6570 -13430
rect 8330 -13490 8390 -13430
rect 8430 -13490 8490 -13430
rect 8530 -13490 8590 -13430
rect 6310 -13590 6370 -13530
rect 6410 -13590 6470 -13530
rect 6510 -13590 6570 -13530
rect 8330 -13590 8390 -13530
rect 8430 -13590 8490 -13530
rect 8530 -13590 8590 -13530
rect 6310 -13680 6370 -13620
rect 6410 -13680 6470 -13620
rect 6510 -13680 6570 -13620
rect 8330 -13680 8390 -13620
rect 8430 -13680 8490 -13620
rect 8530 -13680 8590 -13620
rect 6310 -13770 6370 -13710
rect 6410 -13770 6470 -13710
rect 6510 -13770 6570 -13710
rect 8330 -13770 8390 -13710
rect 8430 -13770 8490 -13710
rect 8530 -13770 8590 -13710
rect 21630 -14090 21700 -14020
rect 21730 -14090 21800 -14020
rect 21830 -14090 21900 -14020
rect 21630 -14190 21700 -14120
rect 21730 -14190 21800 -14120
rect 21830 -14190 21900 -14120
rect 21630 -14290 21700 -14220
rect 21730 -14290 21800 -14220
rect 21830 -14290 21900 -14220
rect 22920 -14940 22990 -14870
rect 23020 -14940 23090 -14870
rect 23120 -14940 23190 -14870
rect 22920 -15040 22990 -14970
rect 23020 -15040 23090 -14970
rect 23120 -15040 23190 -14970
rect 22920 -15140 22990 -15070
rect 23020 -15140 23090 -15070
rect 23120 -15140 23190 -15070
rect 4980 -17160 5040 -17100
rect 5080 -17160 5140 -17100
rect 5180 -17160 5240 -17100
rect 9660 -17160 9720 -17100
rect 9760 -17160 9820 -17100
rect 9860 -17160 9920 -17100
rect 4980 -17260 5040 -17200
rect 5080 -17260 5140 -17200
rect 5180 -17260 5240 -17200
rect 9660 -17260 9720 -17200
rect 9760 -17260 9820 -17200
rect 9860 -17260 9920 -17200
rect 4980 -17360 5040 -17300
rect 5080 -17360 5140 -17300
rect 5180 -17360 5240 -17300
rect 9660 -17360 9720 -17300
rect 9760 -17360 9820 -17300
rect 9860 -17360 9920 -17300
rect 6460 -17820 6530 -17750
rect 6560 -17820 6630 -17750
rect 6660 -17820 6730 -17750
rect 6460 -17930 6530 -17860
rect 6560 -17930 6630 -17860
rect 6660 -17930 6730 -17860
rect 6460 -18040 6530 -17970
rect 6560 -18040 6630 -17970
rect 6660 -18040 6730 -17970
rect 6460 -18150 6530 -18080
rect 6560 -18150 6630 -18080
rect 6660 -18150 6730 -18080
rect 8170 -17820 8240 -17750
rect 8270 -17820 8340 -17750
rect 8370 -17820 8440 -17750
rect 8170 -17930 8240 -17860
rect 8270 -17930 8340 -17860
rect 8370 -17930 8440 -17860
rect 8170 -18040 8240 -17970
rect 8270 -18040 8340 -17970
rect 8370 -18040 8440 -17970
rect 8170 -18150 8240 -18080
rect 8270 -18150 8340 -18080
rect 8370 -18150 8440 -18080
rect 21630 -20170 21700 -20100
rect 21730 -20170 21800 -20100
rect 21830 -20170 21900 -20100
rect 21630 -20270 21700 -20200
rect 21730 -20270 21800 -20200
rect 21830 -20270 21900 -20200
rect 21630 -20370 21700 -20300
rect 21730 -20370 21800 -20300
rect 21830 -20370 21900 -20300
rect 22700 -20800 22770 -20730
rect 22800 -20800 22870 -20730
rect 22900 -20800 22970 -20730
rect 22700 -20900 22770 -20830
rect 22800 -20900 22870 -20830
rect 22900 -20900 22970 -20830
rect 22700 -21000 22770 -20930
rect 22800 -21000 22870 -20930
rect 22900 -21000 22970 -20930
rect 1620 -22730 1690 -22660
rect 1730 -22730 1800 -22660
rect 1840 -22730 1910 -22660
rect 1950 -22730 2020 -22660
rect 2060 -22730 2130 -22660
rect 2170 -22730 2240 -22660
rect 2280 -22730 2350 -22660
rect 2390 -22730 2460 -22660
rect 2500 -22730 2570 -22660
rect 2610 -22730 2680 -22660
rect 2720 -22730 2790 -22660
rect 2830 -22730 2900 -22660
rect 2940 -22730 3010 -22660
rect 3050 -22730 3120 -22660
rect 1620 -22840 1690 -22770
rect 1730 -22840 1800 -22770
rect 1840 -22840 1910 -22770
rect 1950 -22840 2020 -22770
rect 2060 -22840 2130 -22770
rect 2170 -22840 2240 -22770
rect 2280 -22840 2350 -22770
rect 2390 -22840 2460 -22770
rect 2500 -22840 2570 -22770
rect 2610 -22840 2680 -22770
rect 2720 -22840 2790 -22770
rect 2830 -22840 2900 -22770
rect 2940 -22840 3010 -22770
rect 3050 -22840 3120 -22770
rect 11820 -22730 11890 -22660
rect 11930 -22730 12000 -22660
rect 12040 -22730 12110 -22660
rect 12150 -22730 12220 -22660
rect 12260 -22730 12330 -22660
rect 12370 -22730 12440 -22660
rect 12480 -22730 12550 -22660
rect 12590 -22730 12660 -22660
rect 12700 -22730 12770 -22660
rect 12810 -22730 12880 -22660
rect 12920 -22730 12990 -22660
rect 13030 -22730 13100 -22660
rect 13140 -22730 13210 -22660
rect 13250 -22730 13320 -22660
rect 11820 -22840 11890 -22770
rect 11930 -22840 12000 -22770
rect 12040 -22840 12110 -22770
rect 12150 -22840 12220 -22770
rect 12260 -22840 12330 -22770
rect 12370 -22840 12440 -22770
rect 12480 -22840 12550 -22770
rect 12590 -22840 12660 -22770
rect 12700 -22840 12770 -22770
rect 12810 -22840 12880 -22770
rect 12920 -22840 12990 -22770
rect 13030 -22840 13100 -22770
rect 13140 -22840 13210 -22770
rect 13250 -22840 13320 -22770
<< metal2 >>
rect 23460 7210 23940 7260
rect 23460 7140 23490 7210
rect 23560 7140 23600 7210
rect 23670 7140 23710 7210
rect 23780 7140 23820 7210
rect 23890 7140 23940 7210
rect 23460 7100 23940 7140
rect 23460 7030 23490 7100
rect 23560 7030 23600 7100
rect 23670 7030 23710 7100
rect 23780 7030 23820 7100
rect 23890 7030 23940 7100
rect 23460 7000 23940 7030
rect 25860 7210 26340 7260
rect 25860 7140 25890 7210
rect 25960 7140 26000 7210
rect 26070 7140 26110 7210
rect 26180 7140 26220 7210
rect 26290 7140 26340 7210
rect 25860 7100 26340 7140
rect 25860 7030 25890 7100
rect 25960 7030 26000 7100
rect 26070 7030 26110 7100
rect 26180 7030 26220 7100
rect 26290 7030 26340 7100
rect 25860 7000 26340 7030
rect 1540 6850 3140 6900
rect 1540 6780 1570 6850
rect 1640 6780 1680 6850
rect 1750 6780 1790 6850
rect 1860 6780 1900 6850
rect 1970 6780 2010 6850
rect 2080 6780 2120 6850
rect 2190 6780 2230 6850
rect 2300 6780 2340 6850
rect 2410 6780 2450 6850
rect 2520 6780 2560 6850
rect 2630 6780 2670 6850
rect 2740 6780 2780 6850
rect 2850 6780 2890 6850
rect 2960 6780 3000 6850
rect 3070 6780 3140 6850
rect 1540 6740 3140 6780
rect 1540 6670 1570 6740
rect 1640 6670 1680 6740
rect 1750 6670 1790 6740
rect 1860 6670 1900 6740
rect 1970 6670 2010 6740
rect 2080 6670 2120 6740
rect 2190 6670 2230 6740
rect 2300 6670 2340 6740
rect 2410 6670 2450 6740
rect 2520 6670 2560 6740
rect 2630 6670 2670 6740
rect 2740 6670 2780 6740
rect 2850 6670 2890 6740
rect 2960 6670 3000 6740
rect 3070 6670 3140 6740
rect 11760 6880 13360 6930
rect 11760 6810 11790 6880
rect 11860 6810 11900 6880
rect 11970 6810 12010 6880
rect 12080 6810 12120 6880
rect 12190 6810 12230 6880
rect 12300 6810 12340 6880
rect 12410 6810 12450 6880
rect 12520 6810 12560 6880
rect 12630 6810 12670 6880
rect 12740 6810 12780 6880
rect 12850 6810 12890 6880
rect 12960 6810 13000 6880
rect 13070 6810 13110 6880
rect 13180 6810 13220 6880
rect 13290 6810 13360 6880
rect 11760 6770 13360 6810
rect 11760 6700 11790 6770
rect 11860 6700 11900 6770
rect 11970 6700 12010 6770
rect 12080 6700 12120 6770
rect 12190 6700 12230 6770
rect 12300 6700 12340 6770
rect 12410 6700 12450 6770
rect 12520 6700 12560 6770
rect 12630 6700 12670 6770
rect 12740 6700 12780 6770
rect 12850 6700 12890 6770
rect 12960 6700 13000 6770
rect 13070 6700 13110 6770
rect 13180 6700 13220 6770
rect 13290 6700 13360 6770
rect 11760 6670 13360 6700
rect 1540 6640 3140 6670
rect -7150 6300 30940 6320
rect -7150 6290 30740 6300
rect -7150 6230 7380 6290
rect 7440 6230 7480 6290
rect 7540 6280 30740 6290
rect 7540 6230 22780 6280
rect -7150 6210 22780 6230
rect 22850 6210 22890 6280
rect 22960 6210 23000 6280
rect 23070 6210 23110 6280
rect 23180 6230 30740 6280
rect 30810 6230 30850 6300
rect 30920 6230 30940 6300
rect 23180 6210 30940 6230
rect -7150 6190 30940 6210
rect -7150 6080 7380 6190
rect 7440 6080 7480 6190
rect 7540 6170 30940 6190
rect 7540 6100 22780 6170
rect 22850 6100 22890 6170
rect 22960 6100 23000 6170
rect 23070 6100 23110 6170
rect 23180 6100 30740 6170
rect 30810 6100 30850 6170
rect 30920 6100 30940 6170
rect 7540 6080 30940 6100
rect -7150 6060 30940 6080
rect -7150 6040 22780 6060
rect -7150 5980 7380 6040
rect 7440 5980 7480 6040
rect 7540 5990 22780 6040
rect 22850 5990 22890 6060
rect 22960 5990 23000 6060
rect 23070 5990 23110 6060
rect 23180 6040 30940 6060
rect 23180 5990 30740 6040
rect 7540 5980 30740 5990
rect -7150 5970 30740 5980
rect 30810 5970 30850 6040
rect 30920 5970 30940 6040
rect -7150 5950 30940 5970
rect 21800 5670 22020 5690
rect 21800 5600 21820 5670
rect 21890 5600 21930 5670
rect 22000 5600 22020 5670
rect 21800 5560 22020 5600
rect 21800 5490 21820 5560
rect 21890 5490 21930 5560
rect 22000 5490 22020 5560
rect 21800 5450 22020 5490
rect 7400 5390 7490 5410
rect 7400 5320 7410 5390
rect 7480 5320 7490 5390
rect 7400 5280 7490 5320
rect 7400 5210 7410 5280
rect 7480 5210 7490 5280
rect 7400 5170 7490 5210
rect 7400 5100 7410 5170
rect 7480 5100 7490 5170
rect 7400 5060 7490 5100
rect 7400 4990 7410 5060
rect 7480 4990 7490 5060
rect 7400 4950 7490 4990
rect 7400 4880 7410 4950
rect 7480 4880 7490 4950
rect 7400 4860 7490 4880
rect 21800 5380 21820 5450
rect 21890 5380 21930 5450
rect 22000 5380 22020 5450
rect 21800 5340 22020 5380
rect 21800 5270 21820 5340
rect 21890 5270 21930 5340
rect 22000 5270 22020 5340
rect 21800 5230 22020 5270
rect 21800 5160 21820 5230
rect 21890 5160 21930 5230
rect 22000 5160 22020 5230
rect 21800 5120 22020 5160
rect 21800 5050 21820 5120
rect 21890 5050 21930 5120
rect 22000 5050 22020 5120
rect 21800 5010 22020 5050
rect 21800 4940 21820 5010
rect 21890 4940 21930 5010
rect 22000 4940 22020 5010
rect 21800 4900 22020 4940
rect 21800 4830 21820 4900
rect 21890 4830 21930 4900
rect 22000 4830 22020 4900
rect 21800 4790 22020 4830
rect 8140 4760 8460 4790
rect 8140 4700 8170 4760
rect 8230 4700 8270 4760
rect 8330 4700 8370 4760
rect 8430 4700 8460 4760
rect 8140 4610 8460 4700
rect 21800 4720 21820 4790
rect 21890 4720 21930 4790
rect 22000 4720 22020 4790
rect 21800 4680 22020 4720
rect 21800 4610 21820 4680
rect 21890 4610 21930 4680
rect 22000 4610 22020 4680
rect -2520 4580 -2380 4610
rect -2520 4510 -2490 4580
rect -2420 4510 -2380 4580
rect -2520 4470 -2380 4510
rect -2520 4400 -2490 4470
rect -2420 4400 -2380 4470
rect -2520 4360 -2380 4400
rect -2520 4290 -2490 4360
rect -2420 4290 -2380 4360
rect -2520 4250 -2380 4290
rect -2520 4180 -2490 4250
rect -2420 4180 -2380 4250
rect -2520 4130 -2380 4180
rect 6090 4580 8460 4610
rect 6090 4520 6120 4580
rect 6180 4520 8460 4580
rect 6090 4460 8460 4520
rect 6090 4400 6120 4460
rect 6180 4400 8460 4460
rect 6090 4340 8460 4400
rect 6090 4280 6120 4340
rect 6180 4280 8460 4340
rect 6090 4220 8460 4280
rect 6090 4160 6120 4220
rect 6180 4160 8460 4220
rect 6090 4130 8460 4160
rect 17160 4580 17300 4610
rect 17160 4510 17200 4580
rect 17270 4510 17300 4580
rect 17160 4470 17300 4510
rect 21800 4570 22020 4610
rect 21800 4500 21820 4570
rect 21890 4500 21930 4570
rect 22000 4500 22020 4570
rect 21800 4480 22020 4500
rect 27680 4870 28280 4900
rect 27680 4810 27710 4870
rect 27770 4810 27810 4870
rect 27870 4810 27910 4870
rect 27970 4810 28280 4870
rect 27680 4770 28280 4810
rect 27680 4710 27710 4770
rect 27770 4710 27810 4770
rect 27870 4710 27910 4770
rect 27970 4710 28280 4770
rect 27680 4670 28280 4710
rect 27680 4610 27710 4670
rect 27770 4610 27810 4670
rect 27870 4610 27910 4670
rect 27970 4610 28280 4670
rect 27680 4570 28280 4610
rect 27680 4510 27710 4570
rect 27770 4510 27810 4570
rect 27870 4510 27910 4570
rect 27970 4510 28280 4570
rect 17160 4400 17200 4470
rect 17270 4400 17300 4470
rect 17160 4360 17300 4400
rect 17160 4290 17200 4360
rect 17270 4290 17300 4360
rect 17160 4250 17300 4290
rect 17160 4180 17200 4250
rect 17270 4180 17300 4250
rect 17160 4130 17300 4180
rect 27680 4470 28280 4510
rect 27680 4410 27710 4470
rect 27770 4410 27810 4470
rect 27870 4410 27910 4470
rect 27970 4410 28280 4470
rect 27680 4370 28280 4410
rect 27680 4310 27710 4370
rect 27770 4310 27810 4370
rect 27870 4310 27910 4370
rect 27970 4310 28280 4370
rect 27680 4270 28280 4310
rect 27680 4210 27710 4270
rect 27770 4210 27810 4270
rect 27870 4210 27910 4270
rect 27970 4210 28280 4270
rect 27680 4170 28280 4210
rect 8140 3310 8460 4130
rect 27680 4110 27710 4170
rect 27770 4110 27810 4170
rect 27870 4110 27910 4170
rect 27970 4110 28280 4170
rect 27680 4070 28280 4110
rect 27680 4010 27710 4070
rect 27770 4010 27810 4070
rect 27870 4010 27910 4070
rect 27970 4010 28280 4070
rect 27680 3980 28280 4010
rect 7020 3280 7340 3310
rect 7020 3220 7050 3280
rect 7110 3220 7150 3280
rect 7210 3220 7250 3280
rect 7310 3220 7340 3280
rect 7020 3180 7340 3220
rect 7020 3120 7050 3180
rect 7110 3120 7150 3180
rect 7210 3120 7250 3180
rect 7310 3120 7340 3180
rect 7020 3080 7340 3120
rect 7020 3020 7050 3080
rect 7110 3020 7150 3080
rect 7210 3020 7250 3080
rect 7310 3020 7340 3080
rect 7020 3000 7340 3020
rect 7560 3280 8460 3310
rect 7560 3220 7590 3280
rect 7650 3220 7690 3280
rect 7750 3220 7790 3280
rect 7850 3220 8460 3280
rect 7560 3180 8460 3220
rect 7560 3120 7590 3180
rect 7650 3120 7690 3180
rect 7750 3120 7790 3180
rect 7850 3120 8460 3180
rect 7560 3080 8460 3120
rect 7560 3020 7590 3080
rect 7650 3020 7690 3080
rect 7750 3020 7790 3080
rect 7850 3020 8460 3080
rect 24700 3360 25030 3380
rect 24700 3290 24720 3360
rect 24790 3290 24830 3360
rect 24900 3290 24940 3360
rect 25010 3290 25030 3360
rect 24700 3250 25030 3290
rect 24700 3180 24720 3250
rect 24790 3180 24830 3250
rect 24900 3180 24940 3250
rect 25010 3180 25030 3250
rect 24700 3140 25030 3180
rect 24700 3070 24720 3140
rect 24790 3070 24830 3140
rect 24900 3070 24940 3140
rect 25010 3070 25030 3140
rect 24700 3050 25030 3070
rect 7560 3000 8460 3020
rect 4740 2890 5060 2920
rect 4740 2830 4770 2890
rect 4830 2830 4870 2890
rect 4930 2830 4970 2890
rect 5030 2830 5060 2890
rect 4740 2790 5060 2830
rect 4740 2730 4770 2790
rect 4830 2730 4870 2790
rect 4930 2730 4970 2790
rect 5030 2730 5060 2790
rect 4740 2690 5060 2730
rect 4740 2630 4770 2690
rect 4830 2630 4870 2690
rect 4930 2630 4970 2690
rect 5030 2630 5060 2690
rect 4740 2610 5060 2630
rect 9840 2890 10160 2920
rect 9840 2830 9870 2890
rect 9930 2830 9970 2890
rect 10030 2830 10070 2890
rect 10130 2830 10160 2890
rect 9840 2790 10160 2830
rect 9840 2730 9870 2790
rect 9930 2730 9970 2790
rect 10030 2730 10070 2790
rect 10130 2730 10160 2790
rect 9840 2690 10160 2730
rect 9840 2630 9870 2690
rect 9930 2630 9970 2690
rect 10030 2630 10070 2690
rect 10130 2630 10160 2690
rect 9840 2610 10160 2630
rect 22420 2600 22900 2630
rect 22420 2530 22470 2600
rect 22540 2530 22580 2600
rect 22650 2530 22690 2600
rect 22760 2530 22800 2600
rect 22870 2530 22900 2600
rect 22420 2490 22900 2530
rect 22420 2420 22470 2490
rect 22540 2420 22580 2490
rect 22650 2420 22690 2490
rect 22760 2420 22800 2490
rect 22870 2420 22900 2490
rect 22420 2370 22900 2420
rect 26900 2600 27380 2630
rect 26900 2530 26950 2600
rect 27020 2530 27060 2600
rect 27130 2530 27170 2600
rect 27240 2530 27280 2600
rect 27350 2530 27380 2600
rect 26900 2490 27380 2530
rect 26900 2420 26950 2490
rect 27020 2420 27060 2490
rect 27130 2420 27170 2490
rect 27240 2420 27280 2490
rect 27350 2420 27380 2490
rect 26900 2370 27380 2420
rect 28040 1980 28280 3980
rect -7150 1740 -1740 1980
rect -1600 1740 28280 1980
rect 0 1160 310 1180
rect 0 1090 20 1160
rect 90 1090 130 1160
rect 200 1090 230 1160
rect 300 1090 310 1160
rect 0 1050 310 1090
rect 0 980 20 1050
rect 90 980 130 1050
rect 200 980 230 1050
rect 300 980 310 1050
rect 0 940 310 980
rect 0 870 20 940
rect 90 870 130 940
rect 200 870 230 940
rect 300 870 310 940
rect 0 850 310 870
rect -330 -140 150 -100
rect -330 -210 -300 -140
rect -230 -210 -190 -140
rect -120 -210 -80 -140
rect -10 -210 30 -140
rect 100 -210 150 -140
rect -330 -270 150 -210
rect -330 -340 -300 -270
rect -230 -340 -190 -270
rect -120 -340 -80 -270
rect -10 -340 30 -270
rect 100 -340 150 -270
rect -330 -380 150 -340
rect 7150 -120 7630 1740
rect 14590 1160 14900 1180
rect 14590 1090 14600 1160
rect 14670 1090 14700 1160
rect 14770 1090 14810 1160
rect 14880 1090 14900 1160
rect 14590 1050 14900 1090
rect 14590 980 14600 1050
rect 14670 980 14700 1050
rect 14770 980 14810 1050
rect 14880 980 14900 1050
rect 14590 940 14900 980
rect 14590 870 14600 940
rect 14670 870 14700 940
rect 14770 870 14810 940
rect 14880 870 14900 940
rect 14590 850 14900 870
rect 23460 920 23940 970
rect 23460 850 23490 920
rect 23560 850 23600 920
rect 23670 850 23710 920
rect 23780 850 23820 920
rect 23890 850 23940 920
rect 23460 810 23940 850
rect 23460 740 23490 810
rect 23560 740 23600 810
rect 23670 740 23710 810
rect 23780 740 23820 810
rect 23890 740 23940 810
rect 23460 710 23940 740
rect 25860 920 26340 970
rect 25860 850 25890 920
rect 25960 850 26000 920
rect 26070 850 26110 920
rect 26180 850 26220 920
rect 26290 850 26340 920
rect 25860 810 26340 850
rect 25860 740 25890 810
rect 25960 740 26000 810
rect 26070 740 26110 810
rect 26180 740 26220 810
rect 26290 740 26340 810
rect 25860 710 26340 740
rect 19440 0 30940 20
rect 19440 -20 30740 0
rect 19440 -90 22780 -20
rect 22850 -90 22890 -20
rect 22960 -90 23000 -20
rect 23070 -90 23110 -20
rect 23180 -70 30740 -20
rect 30810 -70 30850 0
rect 30920 -70 30940 0
rect 23180 -90 30940 -70
rect 7150 -180 7180 -120
rect 7240 -180 7280 -120
rect 7340 -180 7440 -120
rect 7500 -180 7540 -120
rect 7600 -180 7630 -120
rect 7150 -210 7630 -180
rect 7150 -270 7180 -210
rect 7240 -270 7280 -210
rect 7340 -270 7440 -210
rect 7500 -270 7540 -210
rect 7600 -270 7630 -210
rect 7150 -300 7630 -270
rect 7150 -360 7180 -300
rect 7240 -360 7280 -300
rect 7340 -360 7440 -300
rect 7500 -360 7540 -300
rect 7600 -360 7630 -300
rect 7150 -380 7630 -360
rect 14630 -140 15110 -100
rect 14630 -210 14660 -140
rect 14730 -210 14770 -140
rect 14840 -210 14880 -140
rect 14950 -210 14990 -140
rect 15060 -210 15110 -140
rect 14630 -270 15110 -210
rect 14630 -340 14660 -270
rect 14730 -340 14770 -270
rect 14840 -340 14880 -270
rect 14950 -340 14990 -270
rect 15060 -340 15110 -270
rect 14630 -380 15110 -340
rect 19440 -130 30940 -90
rect 19440 -200 22780 -130
rect 22850 -200 22890 -130
rect 22960 -200 23000 -130
rect 23070 -200 23110 -130
rect 23180 -200 30740 -130
rect 30810 -200 30850 -130
rect 30920 -200 30940 -130
rect 19440 -240 30940 -200
rect 19440 -310 22780 -240
rect 22850 -310 22890 -240
rect 22960 -310 23000 -240
rect 23070 -310 23110 -240
rect 23180 -260 30940 -240
rect 23180 -310 30740 -260
rect 19440 -330 30740 -310
rect 30810 -330 30850 -260
rect 30920 -330 30940 -260
rect 19440 -350 30940 -330
rect 1080 -790 2680 -760
rect 1080 -860 1150 -790
rect 1220 -860 1260 -790
rect 1330 -860 1370 -790
rect 1440 -860 1480 -790
rect 1550 -860 1590 -790
rect 1660 -860 1700 -790
rect 1770 -860 1810 -790
rect 1880 -860 1920 -790
rect 1990 -860 2030 -790
rect 2100 -860 2140 -790
rect 2210 -860 2250 -790
rect 2320 -860 2360 -790
rect 2430 -860 2470 -790
rect 2540 -860 2580 -790
rect 2650 -860 2680 -790
rect 1080 -900 2680 -860
rect 1080 -970 1150 -900
rect 1220 -970 1260 -900
rect 1330 -970 1370 -900
rect 1440 -970 1480 -900
rect 1550 -970 1590 -900
rect 1660 -970 1700 -900
rect 1770 -970 1810 -900
rect 1880 -970 1920 -900
rect 1990 -970 2030 -900
rect 2100 -970 2140 -900
rect 2210 -970 2250 -900
rect 2320 -970 2360 -900
rect 2430 -970 2470 -900
rect 2540 -970 2580 -900
rect 2650 -970 2680 -900
rect 1080 -1020 2680 -970
rect 12220 -790 13820 -760
rect 12220 -860 12250 -790
rect 12320 -860 12360 -790
rect 12430 -860 12470 -790
rect 12540 -860 12580 -790
rect 12650 -860 12690 -790
rect 12760 -860 12800 -790
rect 12870 -860 12910 -790
rect 12980 -860 13020 -790
rect 13090 -860 13130 -790
rect 13200 -860 13240 -790
rect 13310 -860 13350 -790
rect 13420 -860 13460 -790
rect 13530 -860 13570 -790
rect 13640 -860 13680 -790
rect 13750 -860 13820 -790
rect 12220 -900 13820 -860
rect 12220 -970 12250 -900
rect 12320 -970 12360 -900
rect 12430 -970 12470 -900
rect 12540 -970 12580 -900
rect 12650 -970 12690 -900
rect 12760 -970 12800 -900
rect 12870 -970 12910 -900
rect 12980 -970 13020 -900
rect 13090 -970 13130 -900
rect 13200 -970 13240 -900
rect 13310 -970 13350 -900
rect 13420 -970 13460 -900
rect 13530 -970 13570 -900
rect 13640 -970 13680 -900
rect 13750 -970 13820 -900
rect 12220 -1020 13820 -970
rect 1540 -2780 3140 -2730
rect 1540 -2850 1570 -2780
rect 1640 -2850 1680 -2780
rect 1750 -2850 1790 -2780
rect 1860 -2850 1900 -2780
rect 1970 -2850 2010 -2780
rect 2080 -2850 2120 -2780
rect 2190 -2850 2230 -2780
rect 2300 -2850 2340 -2780
rect 2410 -2850 2450 -2780
rect 2520 -2850 2560 -2780
rect 2630 -2850 2670 -2780
rect 2740 -2850 2780 -2780
rect 2850 -2850 2890 -2780
rect 2960 -2850 3000 -2780
rect 3070 -2850 3140 -2780
rect 1540 -2890 3140 -2850
rect 1540 -2960 1570 -2890
rect 1640 -2960 1680 -2890
rect 1750 -2960 1790 -2890
rect 1860 -2960 1900 -2890
rect 1970 -2960 2010 -2890
rect 2080 -2960 2120 -2890
rect 2190 -2960 2230 -2890
rect 2300 -2960 2340 -2890
rect 2410 -2960 2450 -2890
rect 2520 -2960 2560 -2890
rect 2630 -2960 2670 -2890
rect 2740 -2960 2780 -2890
rect 2850 -2960 2890 -2890
rect 2960 -2960 3000 -2890
rect 3070 -2960 3140 -2890
rect 1540 -2990 3140 -2960
rect 11760 -2780 13360 -2730
rect 11760 -2850 11790 -2780
rect 11860 -2850 11900 -2780
rect 11970 -2850 12010 -2780
rect 12080 -2850 12120 -2780
rect 12190 -2850 12230 -2780
rect 12300 -2850 12340 -2780
rect 12410 -2850 12450 -2780
rect 12520 -2850 12560 -2780
rect 12630 -2850 12670 -2780
rect 12740 -2850 12780 -2780
rect 12850 -2850 12890 -2780
rect 12960 -2850 13000 -2780
rect 13070 -2850 13110 -2780
rect 13180 -2850 13220 -2780
rect 13290 -2850 13360 -2780
rect 11760 -2890 13360 -2850
rect 11760 -2960 11790 -2890
rect 11860 -2960 11900 -2890
rect 11970 -2960 12010 -2890
rect 12080 -2960 12120 -2890
rect 12190 -2960 12230 -2890
rect 12300 -2960 12340 -2890
rect 12410 -2960 12450 -2890
rect 12520 -2960 12560 -2890
rect 12630 -2960 12670 -2890
rect 12740 -2960 12780 -2890
rect 12850 -2960 12890 -2890
rect 12960 -2960 13000 -2890
rect 13070 -2960 13110 -2890
rect 13180 -2960 13220 -2890
rect 13290 -2960 13360 -2890
rect 11760 -2990 13360 -2960
rect 19440 -3310 19680 -350
rect 21800 -850 22020 -830
rect 21800 -920 21820 -850
rect 21890 -920 21930 -850
rect 22000 -920 22020 -850
rect 21800 -960 22020 -920
rect 21800 -1030 21820 -960
rect 21890 -1030 21930 -960
rect 22000 -1030 22020 -960
rect 21800 -1070 22020 -1030
rect 21800 -1140 21820 -1070
rect 21890 -1140 21930 -1070
rect 22000 -1140 22020 -1070
rect 21800 -1180 22020 -1140
rect 21800 -1250 21820 -1180
rect 21890 -1250 21930 -1180
rect 22000 -1250 22020 -1180
rect 21800 -1290 22020 -1250
rect 21800 -1360 21820 -1290
rect 21890 -1360 21930 -1290
rect 22000 -1360 22020 -1290
rect 21800 -1400 22020 -1360
rect 21800 -1470 21820 -1400
rect 21890 -1470 21930 -1400
rect 22000 -1470 22020 -1400
rect 21800 -1510 22020 -1470
rect 21800 -1580 21820 -1510
rect 21890 -1580 21930 -1510
rect 22000 -1580 22020 -1510
rect 21800 -1620 22020 -1580
rect 21800 -1690 21820 -1620
rect 21890 -1690 21930 -1620
rect 22000 -1690 22020 -1620
rect 21800 -1730 22020 -1690
rect 21800 -1800 21820 -1730
rect 21890 -1800 21930 -1730
rect 22000 -1800 22020 -1730
rect 21800 -1840 22020 -1800
rect 21800 -1910 21820 -1840
rect 21890 -1910 21930 -1840
rect 22000 -1910 22020 -1840
rect 21800 -1950 22020 -1910
rect 21800 -2020 21820 -1950
rect 21890 -2020 21930 -1950
rect 22000 -2020 22020 -1950
rect 21800 -2040 22020 -2020
rect 27680 -1430 28280 -1400
rect 27680 -1490 27710 -1430
rect 27770 -1490 27810 -1430
rect 27870 -1490 27910 -1430
rect 27970 -1490 28280 -1430
rect 27680 -1530 28280 -1490
rect 27680 -1590 27710 -1530
rect 27770 -1590 27810 -1530
rect 27870 -1590 27910 -1530
rect 27970 -1590 28280 -1530
rect 27680 -1630 28280 -1590
rect 27680 -1690 27710 -1630
rect 27770 -1690 27810 -1630
rect 27870 -1690 27910 -1630
rect 27970 -1690 28280 -1630
rect 27680 -1730 28280 -1690
rect 27680 -1790 27710 -1730
rect 27770 -1790 27810 -1730
rect 27870 -1790 27910 -1730
rect 27970 -1790 28280 -1730
rect 27680 -1830 28280 -1790
rect 27680 -1890 27710 -1830
rect 27770 -1890 27810 -1830
rect 27870 -1890 27910 -1830
rect 27970 -1890 28280 -1830
rect 27680 -1930 28280 -1890
rect 27680 -1990 27710 -1930
rect 27770 -1990 27810 -1930
rect 27870 -1990 27910 -1930
rect 27970 -1990 28280 -1930
rect 27680 -2030 28280 -1990
rect 27680 -2090 27710 -2030
rect 27770 -2090 27810 -2030
rect 27870 -2090 27910 -2030
rect 27970 -2090 28280 -2030
rect 27680 -2130 28280 -2090
rect 27680 -2190 27710 -2130
rect 27770 -2190 27810 -2130
rect 27870 -2190 27910 -2130
rect 27970 -2190 28280 -2130
rect 27680 -2230 28280 -2190
rect 27680 -2290 27710 -2230
rect 27770 -2290 27810 -2230
rect 27870 -2290 27910 -2230
rect 27970 -2290 28280 -2230
rect 27680 -2320 28280 -2290
rect -7150 -3340 19680 -3310
rect -7150 -3400 7380 -3340
rect 7440 -3400 7480 -3340
rect 7540 -3400 19680 -3340
rect 24720 -3050 25050 -3030
rect 24720 -3120 24740 -3050
rect 24810 -3120 24850 -3050
rect 24920 -3120 24960 -3050
rect 25030 -3120 25050 -3050
rect 24720 -3160 25050 -3120
rect 24720 -3230 24740 -3160
rect 24810 -3230 24850 -3160
rect 24920 -3230 24960 -3160
rect 25030 -3230 25050 -3160
rect 24720 -3270 25050 -3230
rect 24720 -3340 24740 -3270
rect 24810 -3340 24850 -3270
rect 24920 -3340 24960 -3270
rect 25030 -3340 25050 -3270
rect 24720 -3360 25050 -3340
rect -7150 -3440 19680 -3400
rect -7150 -3550 7380 -3440
rect 7440 -3550 7480 -3440
rect 7540 -3550 19680 -3440
rect -7150 -3590 19680 -3550
rect -7150 -3650 7380 -3590
rect 7440 -3650 7480 -3590
rect 7540 -3650 19680 -3590
rect -7150 -3680 19680 -3650
rect 22420 -3690 22900 -3660
rect 22420 -3760 22470 -3690
rect 22540 -3760 22580 -3690
rect 22650 -3760 22690 -3690
rect 22760 -3760 22800 -3690
rect 22870 -3760 22900 -3690
rect 22420 -3800 22900 -3760
rect 7290 -3880 7620 -3860
rect 7290 -3950 7310 -3880
rect 7380 -3950 7420 -3880
rect 7490 -3950 7530 -3880
rect 7600 -3950 7620 -3880
rect 22420 -3870 22470 -3800
rect 22540 -3870 22580 -3800
rect 22650 -3870 22690 -3800
rect 22760 -3870 22800 -3800
rect 22870 -3870 22900 -3800
rect 22420 -3920 22900 -3870
rect 26900 -3690 27380 -3660
rect 26900 -3760 26950 -3690
rect 27020 -3760 27060 -3690
rect 27130 -3760 27170 -3690
rect 27240 -3760 27280 -3690
rect 27350 -3760 27380 -3690
rect 26900 -3800 27380 -3760
rect 26900 -3870 26950 -3800
rect 27020 -3870 27060 -3800
rect 27130 -3870 27170 -3800
rect 27240 -3870 27280 -3800
rect 27350 -3870 27380 -3800
rect 26900 -3920 27380 -3870
rect 7290 -3990 7620 -3950
rect 7290 -4060 7310 -3990
rect 7380 -4060 7420 -3990
rect 7490 -4060 7530 -3990
rect 7600 -4060 7620 -3990
rect 7290 -4100 7620 -4060
rect 7290 -4170 7310 -4100
rect 7380 -4170 7420 -4100
rect 7490 -4170 7530 -4100
rect 7600 -4170 7620 -4100
rect 7290 -4190 7620 -4170
rect -580 -4290 -140 -4270
rect -1350 -4350 -910 -4330
rect -1350 -4420 -1330 -4350
rect -1260 -4420 -1220 -4350
rect -1150 -4420 -1110 -4350
rect -1040 -4420 -1000 -4350
rect -930 -4420 -910 -4350
rect -1350 -4460 -910 -4420
rect -1350 -4530 -1330 -4460
rect -1260 -4530 -1220 -4460
rect -1150 -4530 -1110 -4460
rect -1040 -4530 -1000 -4460
rect -930 -4530 -910 -4460
rect -580 -4360 -560 -4290
rect -490 -4360 -450 -4290
rect -380 -4360 -340 -4290
rect -270 -4360 -230 -4290
rect -160 -4360 -140 -4290
rect -580 -4400 -140 -4360
rect -580 -4470 -560 -4400
rect -490 -4470 -450 -4400
rect -380 -4470 -340 -4400
rect -270 -4470 -230 -4400
rect -160 -4470 -140 -4400
rect -580 -4490 -140 -4470
rect 14920 -4290 15360 -4270
rect 14920 -4360 14940 -4290
rect 15010 -4360 15050 -4290
rect 15120 -4360 15160 -4290
rect 15230 -4360 15270 -4290
rect 15340 -4360 15360 -4290
rect 14920 -4400 15360 -4360
rect 14920 -4470 14940 -4400
rect 15010 -4470 15050 -4400
rect 15120 -4470 15160 -4400
rect 15230 -4470 15270 -4400
rect 15340 -4470 15360 -4400
rect 14920 -4490 15360 -4470
rect 15690 -4350 16130 -4330
rect 15690 -4420 15710 -4350
rect 15780 -4420 15820 -4350
rect 15890 -4420 15930 -4350
rect 16000 -4420 16040 -4350
rect 16110 -4420 16130 -4350
rect 28080 -4370 28280 -2320
rect 15690 -4460 16130 -4420
rect -1350 -4550 -910 -4530
rect 15690 -4530 15710 -4460
rect 15780 -4530 15820 -4460
rect 15890 -4530 15930 -4460
rect 16000 -4530 16040 -4460
rect 16110 -4530 16130 -4460
rect 15690 -4550 16130 -4530
rect 20180 -4600 28280 -4370
rect 7030 -6460 7340 -6420
rect -1740 -6520 -1600 -6470
rect -1740 -6590 -1710 -6520
rect -1640 -6590 -1600 -6520
rect -1740 -6630 -1600 -6590
rect -1740 -6700 -1710 -6630
rect -1640 -6700 -1600 -6630
rect 7030 -6520 7050 -6460
rect 7110 -6520 7150 -6460
rect 7210 -6520 7250 -6460
rect 7310 -6520 7340 -6460
rect 7030 -6560 7340 -6520
rect 7030 -6620 7050 -6560
rect 7110 -6620 7150 -6560
rect 7210 -6620 7250 -6560
rect 7310 -6620 7340 -6560
rect -1740 -6740 -1600 -6700
rect -1740 -6810 -1710 -6740
rect -1640 -6810 -1600 -6740
rect -1740 -6850 -1600 -6810
rect -1740 -6920 -1710 -6850
rect -1640 -6920 -1600 -6850
rect -1740 -6950 -1600 -6920
rect 4740 -6670 5060 -6640
rect 4740 -6730 4770 -6670
rect 4830 -6730 4870 -6670
rect 4930 -6730 4970 -6670
rect 5030 -6730 5060 -6670
rect 4740 -6770 5060 -6730
rect 4740 -6830 4770 -6770
rect 4830 -6830 4870 -6770
rect 4930 -6830 4970 -6770
rect 5030 -6830 5060 -6770
rect 4740 -6870 5060 -6830
rect 7030 -6660 7340 -6620
rect 7030 -6720 7050 -6660
rect 7110 -6720 7150 -6660
rect 7210 -6720 7250 -6660
rect 7310 -6720 7340 -6660
rect 7030 -6760 7340 -6720
rect 7030 -6820 7050 -6760
rect 7110 -6820 7150 -6760
rect 7210 -6820 7250 -6760
rect 7310 -6820 7340 -6760
rect 7030 -6850 7340 -6820
rect 7570 -6460 7870 -6420
rect 7570 -6520 7590 -6460
rect 7650 -6520 7690 -6460
rect 7750 -6520 7790 -6460
rect 7850 -6520 7870 -6460
rect 7570 -6560 7870 -6520
rect 7570 -6620 7590 -6560
rect 7650 -6620 7690 -6560
rect 7750 -6620 7790 -6560
rect 7850 -6620 7870 -6560
rect 7570 -6660 7870 -6620
rect 16380 -6520 16520 -6470
rect 16380 -6590 16420 -6520
rect 16490 -6590 16520 -6520
rect 16380 -6630 16520 -6590
rect 7570 -6720 7590 -6660
rect 7650 -6720 7690 -6660
rect 7750 -6720 7790 -6660
rect 7850 -6720 7870 -6660
rect 7570 -6760 7870 -6720
rect 7570 -6820 7590 -6760
rect 7650 -6820 7690 -6760
rect 7750 -6820 7790 -6760
rect 7850 -6820 7870 -6760
rect 7570 -6850 7870 -6820
rect 9840 -6670 10160 -6640
rect 9840 -6730 9870 -6670
rect 9930 -6730 9970 -6670
rect 10030 -6730 10070 -6670
rect 10130 -6730 10160 -6670
rect 9840 -6770 10160 -6730
rect 9840 -6830 9870 -6770
rect 9930 -6830 9970 -6770
rect 10030 -6830 10070 -6770
rect 10130 -6830 10160 -6770
rect 4740 -6930 4770 -6870
rect 4830 -6930 4870 -6870
rect 4930 -6930 4970 -6870
rect 5030 -6930 5060 -6870
rect 4740 -6950 5060 -6930
rect 9840 -6870 10160 -6830
rect 9840 -6930 9870 -6870
rect 9930 -6930 9970 -6870
rect 10030 -6930 10070 -6870
rect 10130 -6930 10160 -6870
rect 9840 -6950 10160 -6930
rect 16380 -6700 16420 -6630
rect 16490 -6700 16520 -6630
rect 16380 -6740 16520 -6700
rect 16380 -6810 16420 -6740
rect 16490 -6810 16520 -6740
rect 16380 -6850 16520 -6810
rect 16380 -6920 16420 -6850
rect 16490 -6920 16520 -6850
rect 16380 -6950 16520 -6920
rect 0 -8140 310 -8120
rect 0 -8210 20 -8140
rect 90 -8210 130 -8140
rect 200 -8210 230 -8140
rect 300 -8210 310 -8140
rect 0 -8250 310 -8210
rect 0 -8320 20 -8250
rect 90 -8320 130 -8250
rect 200 -8320 230 -8250
rect 300 -8320 310 -8250
rect 0 -8360 310 -8320
rect 0 -8430 20 -8360
rect 90 -8430 130 -8360
rect 200 -8430 230 -8360
rect 300 -8430 310 -8360
rect 0 -8450 310 -8430
rect 14590 -8230 14900 -8210
rect 14590 -8300 14600 -8230
rect 14670 -8300 14700 -8230
rect 14770 -8300 14810 -8230
rect 14880 -8300 14900 -8230
rect 14590 -8340 14900 -8300
rect 14590 -8410 14600 -8340
rect 14670 -8410 14700 -8340
rect 14770 -8410 14810 -8340
rect 14880 -8410 14900 -8340
rect 14590 -8450 14900 -8410
rect 14590 -8520 14600 -8450
rect 14670 -8520 14700 -8450
rect 14770 -8520 14810 -8450
rect 14880 -8520 14900 -8450
rect 14590 -8540 14900 -8520
rect 20180 -9160 20490 -4600
rect 21610 -8360 21930 -8330
rect 21610 -8430 21630 -8360
rect 21700 -8430 21730 -8360
rect 21800 -8430 21830 -8360
rect 21900 -8430 21930 -8360
rect 21610 -8460 21930 -8430
rect 21610 -8530 21630 -8460
rect 21700 -8530 21730 -8460
rect 21800 -8530 21830 -8460
rect 21900 -8530 21930 -8460
rect 21610 -8560 21930 -8530
rect 21610 -8630 21630 -8560
rect 21700 -8630 21730 -8560
rect 21800 -8630 21830 -8560
rect 21900 -8630 21930 -8560
rect 21610 -8650 21930 -8630
rect -7150 -9440 20490 -9160
rect 22630 -9010 22950 -8980
rect 22630 -9080 22650 -9010
rect 22720 -9080 22750 -9010
rect 22820 -9080 22850 -9010
rect 22920 -9080 22950 -9010
rect 22630 -9110 22950 -9080
rect 22630 -9180 22650 -9110
rect 22720 -9180 22750 -9110
rect 22820 -9180 22850 -9110
rect 22920 -9180 22950 -9110
rect 22630 -9210 22950 -9180
rect 22630 -9280 22650 -9210
rect 22720 -9280 22750 -9210
rect 22820 -9280 22850 -9210
rect 22920 -9280 22950 -9210
rect 22630 -9300 22950 -9280
rect -270 -9660 210 -9620
rect -270 -9730 -240 -9660
rect -170 -9730 -130 -9660
rect -60 -9730 -20 -9660
rect 50 -9730 90 -9660
rect 160 -9730 210 -9660
rect -270 -9790 210 -9730
rect -270 -9860 -240 -9790
rect -170 -9860 -130 -9790
rect -60 -9860 -20 -9790
rect 50 -9860 90 -9790
rect 160 -9860 210 -9790
rect -270 -9900 210 -9860
rect 7210 -9640 7690 -9440
rect 7210 -9700 7240 -9640
rect 7300 -9700 7340 -9640
rect 7400 -9700 7500 -9640
rect 7560 -9700 7600 -9640
rect 7660 -9700 7690 -9640
rect 7210 -9730 7690 -9700
rect 7210 -9790 7240 -9730
rect 7300 -9790 7340 -9730
rect 7400 -9790 7500 -9730
rect 7560 -9790 7600 -9730
rect 7660 -9790 7690 -9730
rect 7210 -9820 7690 -9790
rect 7210 -9880 7240 -9820
rect 7300 -9880 7340 -9820
rect 7400 -9880 7500 -9820
rect 7560 -9880 7600 -9820
rect 7660 -9880 7690 -9820
rect 7210 -9900 7690 -9880
rect 14690 -9660 15170 -9620
rect 14690 -9730 14720 -9660
rect 14790 -9730 14830 -9660
rect 14900 -9730 14940 -9660
rect 15010 -9730 15050 -9660
rect 15120 -9730 15170 -9660
rect 14690 -9790 15170 -9730
rect 14690 -9860 14720 -9790
rect 14790 -9860 14830 -9790
rect 14900 -9860 14940 -9790
rect 15010 -9860 15050 -9790
rect 15120 -9860 15170 -9790
rect 14690 -9900 15170 -9860
rect 1080 -10340 2680 -10310
rect 1080 -10410 1150 -10340
rect 1220 -10410 1260 -10340
rect 1330 -10410 1370 -10340
rect 1440 -10410 1480 -10340
rect 1550 -10410 1590 -10340
rect 1660 -10410 1700 -10340
rect 1770 -10410 1810 -10340
rect 1880 -10410 1920 -10340
rect 1990 -10410 2030 -10340
rect 2100 -10410 2140 -10340
rect 2210 -10410 2250 -10340
rect 2320 -10410 2360 -10340
rect 2430 -10410 2470 -10340
rect 2540 -10410 2580 -10340
rect 2650 -10410 2680 -10340
rect 1080 -10450 2680 -10410
rect 1080 -10520 1150 -10450
rect 1220 -10520 1260 -10450
rect 1330 -10520 1370 -10450
rect 1440 -10520 1480 -10450
rect 1550 -10520 1590 -10450
rect 1660 -10520 1700 -10450
rect 1770 -10520 1810 -10450
rect 1880 -10520 1920 -10450
rect 1990 -10520 2030 -10450
rect 2100 -10520 2140 -10450
rect 2210 -10520 2250 -10450
rect 2320 -10520 2360 -10450
rect 2430 -10520 2470 -10450
rect 2540 -10520 2580 -10450
rect 2650 -10520 2680 -10450
rect 1080 -10570 2680 -10520
rect 12220 -10370 13820 -10340
rect 12220 -10440 12290 -10370
rect 12360 -10440 12400 -10370
rect 12470 -10440 12510 -10370
rect 12580 -10440 12620 -10370
rect 12690 -10440 12730 -10370
rect 12800 -10440 12840 -10370
rect 12910 -10440 12950 -10370
rect 13020 -10440 13060 -10370
rect 13130 -10440 13170 -10370
rect 13240 -10440 13280 -10370
rect 13350 -10440 13390 -10370
rect 13460 -10440 13500 -10370
rect 13570 -10440 13610 -10370
rect 13680 -10440 13720 -10370
rect 13790 -10440 13820 -10370
rect 12220 -10480 13820 -10440
rect 12220 -10550 12290 -10480
rect 12360 -10550 12400 -10480
rect 12470 -10550 12510 -10480
rect 12580 -10550 12620 -10480
rect 12690 -10550 12730 -10480
rect 12800 -10550 12840 -10480
rect 12910 -10550 12950 -10480
rect 13020 -10550 13060 -10480
rect 13130 -10550 13170 -10480
rect 13240 -10550 13280 -10480
rect 13350 -10550 13390 -10480
rect 13460 -10550 13500 -10480
rect 13570 -10550 13610 -10480
rect 13680 -10550 13720 -10480
rect 13790 -10550 13820 -10480
rect 12220 -10600 13820 -10550
rect 1510 -12300 3110 -12250
rect 1510 -12370 1540 -12300
rect 1610 -12370 1650 -12300
rect 1720 -12370 1760 -12300
rect 1830 -12370 1870 -12300
rect 1940 -12370 1980 -12300
rect 2050 -12370 2090 -12300
rect 2160 -12370 2200 -12300
rect 2270 -12370 2310 -12300
rect 2380 -12370 2420 -12300
rect 2490 -12370 2530 -12300
rect 2600 -12370 2640 -12300
rect 2710 -12370 2750 -12300
rect 2820 -12370 2860 -12300
rect 2930 -12370 2970 -12300
rect 3040 -12370 3110 -12300
rect 1510 -12410 3110 -12370
rect 1510 -12480 1540 -12410
rect 1610 -12480 1650 -12410
rect 1720 -12480 1760 -12410
rect 1830 -12480 1870 -12410
rect 1940 -12480 1980 -12410
rect 2050 -12480 2090 -12410
rect 2160 -12480 2200 -12410
rect 2270 -12480 2310 -12410
rect 2380 -12480 2420 -12410
rect 2490 -12480 2530 -12410
rect 2600 -12480 2640 -12410
rect 2710 -12480 2750 -12410
rect 2820 -12480 2860 -12410
rect 2930 -12480 2970 -12410
rect 3040 -12480 3110 -12410
rect 1510 -12510 3110 -12480
rect 11790 -12300 13390 -12250
rect 11790 -12370 11820 -12300
rect 11890 -12370 11930 -12300
rect 12000 -12370 12040 -12300
rect 12110 -12370 12150 -12300
rect 12220 -12370 12260 -12300
rect 12330 -12370 12370 -12300
rect 12440 -12370 12480 -12300
rect 12550 -12370 12590 -12300
rect 12660 -12370 12700 -12300
rect 12770 -12370 12810 -12300
rect 12880 -12370 12920 -12300
rect 12990 -12370 13030 -12300
rect 13100 -12370 13140 -12300
rect 13210 -12370 13250 -12300
rect 13320 -12370 13390 -12300
rect 11790 -12410 13390 -12370
rect 11790 -12480 11820 -12410
rect 11890 -12480 11930 -12410
rect 12000 -12480 12040 -12410
rect 12110 -12480 12150 -12410
rect 12220 -12480 12260 -12410
rect 12330 -12480 12370 -12410
rect 12440 -12480 12480 -12410
rect 12550 -12480 12590 -12410
rect 12660 -12480 12700 -12410
rect 12770 -12480 12810 -12410
rect 12880 -12480 12920 -12410
rect 12990 -12480 13030 -12410
rect 13100 -12480 13140 -12410
rect 13210 -12480 13250 -12410
rect 13320 -12480 13390 -12410
rect 11790 -12510 13390 -12480
rect 6280 -13250 6610 -13220
rect 6280 -13310 6310 -13250
rect 6370 -13310 6410 -13250
rect 6470 -13310 6510 -13250
rect 6570 -13310 6610 -13250
rect 6280 -13340 6610 -13310
rect 6280 -13400 6310 -13340
rect 6370 -13400 6410 -13340
rect 6470 -13400 6510 -13340
rect 6570 -13400 6610 -13340
rect 6280 -13430 6610 -13400
rect 6280 -13490 6310 -13430
rect 6370 -13490 6410 -13430
rect 6470 -13490 6510 -13430
rect 6570 -13490 6610 -13430
rect 6280 -13530 6610 -13490
rect 6280 -13590 6310 -13530
rect 6370 -13590 6410 -13530
rect 6470 -13590 6510 -13530
rect 6570 -13590 6610 -13530
rect 6280 -13620 6610 -13590
rect 6280 -13680 6310 -13620
rect 6370 -13680 6410 -13620
rect 6470 -13680 6510 -13620
rect 6570 -13680 6610 -13620
rect 6280 -13710 6610 -13680
rect 6280 -13770 6310 -13710
rect 6370 -13770 6410 -13710
rect 6470 -13770 6510 -13710
rect 6570 -13770 6610 -13710
rect 6280 -13800 6610 -13770
rect 8290 -13250 8620 -13220
rect 8290 -13310 8330 -13250
rect 8390 -13310 8430 -13250
rect 8490 -13310 8530 -13250
rect 8590 -13310 8620 -13250
rect 8290 -13340 8620 -13310
rect 8290 -13400 8330 -13340
rect 8390 -13400 8430 -13340
rect 8490 -13400 8530 -13340
rect 8590 -13400 8620 -13340
rect 8290 -13430 8620 -13400
rect 8290 -13490 8330 -13430
rect 8390 -13490 8430 -13430
rect 8490 -13490 8530 -13430
rect 8590 -13490 8620 -13430
rect 8290 -13530 8620 -13490
rect 8290 -13590 8330 -13530
rect 8390 -13590 8430 -13530
rect 8490 -13590 8530 -13530
rect 8590 -13590 8620 -13530
rect 8290 -13620 8620 -13590
rect 8290 -13680 8330 -13620
rect 8390 -13680 8430 -13620
rect 8490 -13680 8530 -13620
rect 8590 -13680 8620 -13620
rect 8290 -13710 8620 -13680
rect 8290 -13770 8330 -13710
rect 8390 -13770 8430 -13710
rect 8490 -13770 8530 -13710
rect 8590 -13770 8620 -13710
rect 8290 -13800 8620 -13770
rect 21610 -14020 21930 -13990
rect 21610 -14090 21630 -14020
rect 21700 -14090 21730 -14020
rect 21800 -14090 21830 -14020
rect 21900 -14090 21930 -14020
rect 21610 -14120 21930 -14090
rect 21610 -14190 21630 -14120
rect 21700 -14190 21730 -14120
rect 21800 -14190 21830 -14120
rect 21900 -14190 21930 -14120
rect 21610 -14220 21930 -14190
rect 21610 -14290 21630 -14220
rect 21700 -14290 21730 -14220
rect 21800 -14290 21830 -14220
rect 21900 -14290 21930 -14220
rect 21610 -14310 21930 -14290
rect 22900 -14870 23220 -14840
rect 22900 -14940 22920 -14870
rect 22990 -14940 23020 -14870
rect 23090 -14940 23120 -14870
rect 23190 -14940 23220 -14870
rect 22900 -14970 23220 -14940
rect 22900 -15040 22920 -14970
rect 22990 -15040 23020 -14970
rect 23090 -15040 23120 -14970
rect 23190 -15040 23220 -14970
rect 22900 -15070 23220 -15040
rect 22900 -15140 22920 -15070
rect 22990 -15140 23020 -15070
rect 23090 -15140 23120 -15070
rect 23190 -15140 23220 -15070
rect 22900 -15160 23220 -15140
rect 4950 -17100 5270 -17070
rect 4950 -17160 4980 -17100
rect 5040 -17160 5080 -17100
rect 5140 -17160 5180 -17100
rect 5240 -17160 5270 -17100
rect 4950 -17200 5270 -17160
rect 4950 -17260 4980 -17200
rect 5040 -17260 5080 -17200
rect 5140 -17260 5180 -17200
rect 5240 -17260 5270 -17200
rect 4950 -17300 5270 -17260
rect 4950 -17360 4980 -17300
rect 5040 -17360 5080 -17300
rect 5140 -17360 5180 -17300
rect 5240 -17360 5270 -17300
rect 4950 -17380 5270 -17360
rect 9630 -17100 9950 -17070
rect 9630 -17160 9660 -17100
rect 9720 -17160 9760 -17100
rect 9820 -17160 9860 -17100
rect 9920 -17160 9950 -17100
rect 9630 -17200 9950 -17160
rect 9630 -17260 9660 -17200
rect 9720 -17260 9760 -17200
rect 9820 -17260 9860 -17200
rect 9920 -17260 9950 -17200
rect 9630 -17300 9950 -17260
rect 9630 -17360 9660 -17300
rect 9720 -17360 9760 -17300
rect 9820 -17360 9860 -17300
rect 9920 -17360 9950 -17300
rect 9630 -17380 9950 -17360
rect 6440 -17750 6750 -17730
rect 6440 -17820 6460 -17750
rect 6530 -17820 6560 -17750
rect 6630 -17820 6660 -17750
rect 6730 -17820 6750 -17750
rect 6440 -17860 6750 -17820
rect 6440 -17930 6460 -17860
rect 6530 -17930 6560 -17860
rect 6630 -17930 6660 -17860
rect 6730 -17930 6750 -17860
rect 6440 -17970 6750 -17930
rect 6440 -18040 6460 -17970
rect 6530 -18040 6560 -17970
rect 6630 -18040 6660 -17970
rect 6730 -18040 6750 -17970
rect 6440 -18080 6750 -18040
rect 6440 -18150 6460 -18080
rect 6530 -18150 6560 -18080
rect 6630 -18150 6660 -18080
rect 6730 -18150 6750 -18080
rect 6440 -18170 6750 -18150
rect 8150 -17750 8460 -17730
rect 8150 -17820 8170 -17750
rect 8240 -17820 8270 -17750
rect 8340 -17820 8370 -17750
rect 8440 -17820 8460 -17750
rect 8150 -17860 8460 -17820
rect 8150 -17930 8170 -17860
rect 8240 -17930 8270 -17860
rect 8340 -17930 8370 -17860
rect 8440 -17930 8460 -17860
rect 8150 -17970 8460 -17930
rect 8150 -18040 8170 -17970
rect 8240 -18040 8270 -17970
rect 8340 -18040 8370 -17970
rect 8440 -18040 8460 -17970
rect 8150 -18080 8460 -18040
rect 8150 -18150 8170 -18080
rect 8240 -18150 8270 -18080
rect 8340 -18150 8370 -18080
rect 8440 -18150 8460 -18080
rect 8150 -18170 8460 -18150
rect 21610 -20100 21930 -20070
rect 21610 -20170 21630 -20100
rect 21700 -20170 21730 -20100
rect 21800 -20170 21830 -20100
rect 21900 -20170 21930 -20100
rect 21610 -20200 21930 -20170
rect 21610 -20270 21630 -20200
rect 21700 -20270 21730 -20200
rect 21800 -20270 21830 -20200
rect 21900 -20270 21930 -20200
rect 21610 -20300 21930 -20270
rect 21610 -20370 21630 -20300
rect 21700 -20370 21730 -20300
rect 21800 -20370 21830 -20300
rect 21900 -20370 21930 -20300
rect 21610 -20390 21930 -20370
rect 22680 -20730 23000 -20700
rect 22680 -20800 22700 -20730
rect 22770 -20800 22800 -20730
rect 22870 -20800 22900 -20730
rect 22970 -20800 23000 -20730
rect 22680 -20830 23000 -20800
rect 22680 -20900 22700 -20830
rect 22770 -20900 22800 -20830
rect 22870 -20900 22900 -20830
rect 22970 -20900 23000 -20830
rect 22680 -20930 23000 -20900
rect 22680 -21000 22700 -20930
rect 22770 -21000 22800 -20930
rect 22870 -21000 22900 -20930
rect 22970 -21000 23000 -20930
rect 22680 -21020 23000 -21000
rect 1550 -22660 3150 -22630
rect 1550 -22730 1620 -22660
rect 1690 -22730 1730 -22660
rect 1800 -22730 1840 -22660
rect 1910 -22730 1950 -22660
rect 2020 -22730 2060 -22660
rect 2130 -22730 2170 -22660
rect 2240 -22730 2280 -22660
rect 2350 -22730 2390 -22660
rect 2460 -22730 2500 -22660
rect 2570 -22730 2610 -22660
rect 2680 -22730 2720 -22660
rect 2790 -22730 2830 -22660
rect 2900 -22730 2940 -22660
rect 3010 -22730 3050 -22660
rect 3120 -22730 3150 -22660
rect 1550 -22770 3150 -22730
rect 1550 -22840 1620 -22770
rect 1690 -22840 1730 -22770
rect 1800 -22840 1840 -22770
rect 1910 -22840 1950 -22770
rect 2020 -22840 2060 -22770
rect 2130 -22840 2170 -22770
rect 2240 -22840 2280 -22770
rect 2350 -22840 2390 -22770
rect 2460 -22840 2500 -22770
rect 2570 -22840 2610 -22770
rect 2680 -22840 2720 -22770
rect 2790 -22840 2830 -22770
rect 2900 -22840 2940 -22770
rect 3010 -22840 3050 -22770
rect 3120 -22840 3150 -22770
rect 1550 -22890 3150 -22840
rect 11750 -22660 13350 -22630
rect 11750 -22730 11820 -22660
rect 11890 -22730 11930 -22660
rect 12000 -22730 12040 -22660
rect 12110 -22730 12150 -22660
rect 12220 -22730 12260 -22660
rect 12330 -22730 12370 -22660
rect 12440 -22730 12480 -22660
rect 12550 -22730 12590 -22660
rect 12660 -22730 12700 -22660
rect 12770 -22730 12810 -22660
rect 12880 -22730 12920 -22660
rect 12990 -22730 13030 -22660
rect 13100 -22730 13140 -22660
rect 13210 -22730 13250 -22660
rect 13320 -22730 13350 -22660
rect 11750 -22770 13350 -22730
rect 11750 -22840 11820 -22770
rect 11890 -22840 11930 -22770
rect 12000 -22840 12040 -22770
rect 12110 -22840 12150 -22770
rect 12220 -22840 12260 -22770
rect 12330 -22840 12370 -22770
rect 12440 -22840 12480 -22770
rect 12550 -22840 12590 -22770
rect 12660 -22840 12700 -22770
rect 12770 -22840 12810 -22770
rect 12880 -22840 12920 -22770
rect 12990 -22840 13030 -22770
rect 13100 -22840 13140 -22770
rect 13210 -22840 13250 -22770
rect 13320 -22840 13350 -22770
rect 11750 -22890 13350 -22840
<< via2 >>
rect 23490 7140 23560 7210
rect 23600 7140 23670 7210
rect 23710 7140 23780 7210
rect 23820 7140 23890 7210
rect 23490 7030 23560 7100
rect 23600 7030 23670 7100
rect 23710 7030 23780 7100
rect 23820 7030 23890 7100
rect 25890 7140 25960 7210
rect 26000 7140 26070 7210
rect 26110 7140 26180 7210
rect 26220 7140 26290 7210
rect 25890 7030 25960 7100
rect 26000 7030 26070 7100
rect 26110 7030 26180 7100
rect 26220 7030 26290 7100
rect 1570 6780 1640 6850
rect 1680 6780 1750 6850
rect 1790 6780 1860 6850
rect 1900 6780 1970 6850
rect 2010 6780 2080 6850
rect 2120 6780 2190 6850
rect 2230 6780 2300 6850
rect 2340 6780 2410 6850
rect 2450 6780 2520 6850
rect 2560 6780 2630 6850
rect 2670 6780 2740 6850
rect 2780 6780 2850 6850
rect 2890 6780 2960 6850
rect 3000 6780 3070 6850
rect 1570 6670 1640 6740
rect 1680 6670 1750 6740
rect 1790 6670 1860 6740
rect 1900 6670 1970 6740
rect 2010 6670 2080 6740
rect 2120 6670 2190 6740
rect 2230 6670 2300 6740
rect 2340 6670 2410 6740
rect 2450 6670 2520 6740
rect 2560 6670 2630 6740
rect 2670 6670 2740 6740
rect 2780 6670 2850 6740
rect 2890 6670 2960 6740
rect 3000 6670 3070 6740
rect 11790 6810 11860 6880
rect 11900 6810 11970 6880
rect 12010 6810 12080 6880
rect 12120 6810 12190 6880
rect 12230 6810 12300 6880
rect 12340 6810 12410 6880
rect 12450 6810 12520 6880
rect 12560 6810 12630 6880
rect 12670 6810 12740 6880
rect 12780 6810 12850 6880
rect 12890 6810 12960 6880
rect 13000 6810 13070 6880
rect 13110 6810 13180 6880
rect 13220 6810 13290 6880
rect 11790 6700 11860 6770
rect 11900 6700 11970 6770
rect 12010 6700 12080 6770
rect 12120 6700 12190 6770
rect 12230 6700 12300 6770
rect 12340 6700 12410 6770
rect 12450 6700 12520 6770
rect 12560 6700 12630 6770
rect 12670 6700 12740 6770
rect 12780 6700 12850 6770
rect 12890 6700 12960 6770
rect 13000 6700 13070 6770
rect 13110 6700 13180 6770
rect 13220 6700 13290 6770
rect 30740 6230 30810 6300
rect 30850 6230 30920 6300
rect 30740 6100 30810 6170
rect 30850 6100 30920 6170
rect 30740 5970 30810 6040
rect 30850 5970 30920 6040
rect 21820 5600 21890 5670
rect 21930 5600 22000 5670
rect 21820 5490 21890 5560
rect 21930 5490 22000 5560
rect 7410 5320 7480 5390
rect 7410 5210 7480 5280
rect 7410 5100 7480 5170
rect 7410 4990 7480 5060
rect 7410 4880 7480 4950
rect 21820 5380 21890 5450
rect 21930 5380 22000 5450
rect 21820 5270 21890 5340
rect 21930 5270 22000 5340
rect 21820 5160 21890 5230
rect 21930 5160 22000 5230
rect 21820 5050 21890 5120
rect 21930 5050 22000 5120
rect 21820 4940 21890 5010
rect 21930 4940 22000 5010
rect 21820 4830 21890 4900
rect 21930 4830 22000 4900
rect 8170 4700 8230 4760
rect 8270 4700 8330 4760
rect 8370 4700 8430 4760
rect 21820 4720 21890 4790
rect 21930 4720 22000 4790
rect 21820 4610 21890 4680
rect 21930 4610 22000 4680
rect -2490 4510 -2420 4580
rect -2490 4400 -2420 4470
rect -2490 4290 -2420 4360
rect -2490 4180 -2420 4250
rect 6120 4520 6180 4580
rect 6120 4400 6180 4460
rect 6120 4280 6180 4340
rect 6120 4160 6180 4220
rect 17200 4510 17270 4580
rect 21820 4500 21890 4570
rect 21930 4500 22000 4570
rect 17200 4400 17270 4470
rect 17200 4290 17270 4360
rect 17200 4180 17270 4250
rect 7050 3220 7110 3280
rect 7150 3220 7210 3280
rect 7250 3220 7310 3280
rect 7050 3120 7110 3180
rect 7150 3120 7210 3180
rect 7250 3120 7310 3180
rect 7050 3020 7110 3080
rect 7150 3020 7210 3080
rect 7250 3020 7310 3080
rect 24720 3290 24790 3360
rect 24830 3290 24900 3360
rect 24940 3290 25010 3360
rect 24720 3180 24790 3250
rect 24830 3180 24900 3250
rect 24940 3180 25010 3250
rect 24720 3070 24790 3140
rect 24830 3070 24900 3140
rect 24940 3070 25010 3140
rect 4770 2830 4830 2890
rect 4870 2830 4930 2890
rect 4970 2830 5030 2890
rect 4770 2730 4830 2790
rect 4870 2730 4930 2790
rect 4970 2730 5030 2790
rect 4770 2630 4830 2690
rect 4870 2630 4930 2690
rect 4970 2630 5030 2690
rect 9870 2830 9930 2890
rect 9970 2830 10030 2890
rect 10070 2830 10130 2890
rect 9870 2730 9930 2790
rect 9970 2730 10030 2790
rect 10070 2730 10130 2790
rect 9870 2630 9930 2690
rect 9970 2630 10030 2690
rect 10070 2630 10130 2690
rect 22470 2530 22540 2600
rect 22580 2530 22650 2600
rect 22690 2530 22760 2600
rect 22800 2530 22870 2600
rect 22470 2420 22540 2490
rect 22580 2420 22650 2490
rect 22690 2420 22760 2490
rect 22800 2420 22870 2490
rect 26950 2530 27020 2600
rect 27060 2530 27130 2600
rect 27170 2530 27240 2600
rect 27280 2530 27350 2600
rect 26950 2420 27020 2490
rect 27060 2420 27130 2490
rect 27170 2420 27240 2490
rect 27280 2420 27350 2490
rect 20 1090 90 1160
rect 130 1090 200 1160
rect 230 1090 300 1160
rect 20 980 90 1050
rect 130 980 200 1050
rect 230 980 300 1050
rect 20 870 90 940
rect 130 870 200 940
rect 230 870 300 940
rect -300 -210 -230 -140
rect -190 -210 -120 -140
rect -80 -210 -10 -140
rect 30 -210 100 -140
rect -300 -340 -230 -270
rect -190 -340 -120 -270
rect -80 -340 -10 -270
rect 30 -340 100 -270
rect 14600 1090 14670 1160
rect 14700 1090 14770 1160
rect 14810 1090 14880 1160
rect 14600 980 14670 1050
rect 14700 980 14770 1050
rect 14810 980 14880 1050
rect 14600 870 14670 940
rect 14700 870 14770 940
rect 14810 870 14880 940
rect 23490 850 23560 920
rect 23600 850 23670 920
rect 23710 850 23780 920
rect 23820 850 23890 920
rect 23490 740 23560 810
rect 23600 740 23670 810
rect 23710 740 23780 810
rect 23820 740 23890 810
rect 25890 850 25960 920
rect 26000 850 26070 920
rect 26110 850 26180 920
rect 26220 850 26290 920
rect 25890 740 25960 810
rect 26000 740 26070 810
rect 26110 740 26180 810
rect 26220 740 26290 810
rect 30740 -70 30810 0
rect 30850 -70 30920 0
rect 14660 -210 14730 -140
rect 14770 -210 14840 -140
rect 14880 -210 14950 -140
rect 14990 -210 15060 -140
rect 14660 -340 14730 -270
rect 14770 -340 14840 -270
rect 14880 -340 14950 -270
rect 14990 -340 15060 -270
rect 30740 -200 30810 -130
rect 30850 -200 30920 -130
rect 30740 -330 30810 -260
rect 30850 -330 30920 -260
rect 1150 -860 1220 -790
rect 1260 -860 1330 -790
rect 1370 -860 1440 -790
rect 1480 -860 1550 -790
rect 1590 -860 1660 -790
rect 1700 -860 1770 -790
rect 1810 -860 1880 -790
rect 1920 -860 1990 -790
rect 2030 -860 2100 -790
rect 2140 -860 2210 -790
rect 2250 -860 2320 -790
rect 2360 -860 2430 -790
rect 2470 -860 2540 -790
rect 2580 -860 2650 -790
rect 1150 -970 1220 -900
rect 1260 -970 1330 -900
rect 1370 -970 1440 -900
rect 1480 -970 1550 -900
rect 1590 -970 1660 -900
rect 1700 -970 1770 -900
rect 1810 -970 1880 -900
rect 1920 -970 1990 -900
rect 2030 -970 2100 -900
rect 2140 -970 2210 -900
rect 2250 -970 2320 -900
rect 2360 -970 2430 -900
rect 2470 -970 2540 -900
rect 2580 -970 2650 -900
rect 12250 -860 12320 -790
rect 12360 -860 12430 -790
rect 12470 -860 12540 -790
rect 12580 -860 12650 -790
rect 12690 -860 12760 -790
rect 12800 -860 12870 -790
rect 12910 -860 12980 -790
rect 13020 -860 13090 -790
rect 13130 -860 13200 -790
rect 13240 -860 13310 -790
rect 13350 -860 13420 -790
rect 13460 -860 13530 -790
rect 13570 -860 13640 -790
rect 13680 -860 13750 -790
rect 12250 -970 12320 -900
rect 12360 -970 12430 -900
rect 12470 -970 12540 -900
rect 12580 -970 12650 -900
rect 12690 -970 12760 -900
rect 12800 -970 12870 -900
rect 12910 -970 12980 -900
rect 13020 -970 13090 -900
rect 13130 -970 13200 -900
rect 13240 -970 13310 -900
rect 13350 -970 13420 -900
rect 13460 -970 13530 -900
rect 13570 -970 13640 -900
rect 13680 -970 13750 -900
rect 1570 -2850 1640 -2780
rect 1680 -2850 1750 -2780
rect 1790 -2850 1860 -2780
rect 1900 -2850 1970 -2780
rect 2010 -2850 2080 -2780
rect 2120 -2850 2190 -2780
rect 2230 -2850 2300 -2780
rect 2340 -2850 2410 -2780
rect 2450 -2850 2520 -2780
rect 2560 -2850 2630 -2780
rect 2670 -2850 2740 -2780
rect 2780 -2850 2850 -2780
rect 2890 -2850 2960 -2780
rect 3000 -2850 3070 -2780
rect 1570 -2960 1640 -2890
rect 1680 -2960 1750 -2890
rect 1790 -2960 1860 -2890
rect 1900 -2960 1970 -2890
rect 2010 -2960 2080 -2890
rect 2120 -2960 2190 -2890
rect 2230 -2960 2300 -2890
rect 2340 -2960 2410 -2890
rect 2450 -2960 2520 -2890
rect 2560 -2960 2630 -2890
rect 2670 -2960 2740 -2890
rect 2780 -2960 2850 -2890
rect 2890 -2960 2960 -2890
rect 3000 -2960 3070 -2890
rect 11790 -2850 11860 -2780
rect 11900 -2850 11970 -2780
rect 12010 -2850 12080 -2780
rect 12120 -2850 12190 -2780
rect 12230 -2850 12300 -2780
rect 12340 -2850 12410 -2780
rect 12450 -2850 12520 -2780
rect 12560 -2850 12630 -2780
rect 12670 -2850 12740 -2780
rect 12780 -2850 12850 -2780
rect 12890 -2850 12960 -2780
rect 13000 -2850 13070 -2780
rect 13110 -2850 13180 -2780
rect 13220 -2850 13290 -2780
rect 11790 -2960 11860 -2890
rect 11900 -2960 11970 -2890
rect 12010 -2960 12080 -2890
rect 12120 -2960 12190 -2890
rect 12230 -2960 12300 -2890
rect 12340 -2960 12410 -2890
rect 12450 -2960 12520 -2890
rect 12560 -2960 12630 -2890
rect 12670 -2960 12740 -2890
rect 12780 -2960 12850 -2890
rect 12890 -2960 12960 -2890
rect 13000 -2960 13070 -2890
rect 13110 -2960 13180 -2890
rect 13220 -2960 13290 -2890
rect 21820 -920 21890 -850
rect 21930 -920 22000 -850
rect 21820 -1030 21890 -960
rect 21930 -1030 22000 -960
rect 21820 -1140 21890 -1070
rect 21930 -1140 22000 -1070
rect 21820 -1250 21890 -1180
rect 21930 -1250 22000 -1180
rect 21820 -1360 21890 -1290
rect 21930 -1360 22000 -1290
rect 21820 -1470 21890 -1400
rect 21930 -1470 22000 -1400
rect 21820 -1580 21890 -1510
rect 21930 -1580 22000 -1510
rect 21820 -1690 21890 -1620
rect 21930 -1690 22000 -1620
rect 21820 -1800 21890 -1730
rect 21930 -1800 22000 -1730
rect 21820 -1910 21890 -1840
rect 21930 -1910 22000 -1840
rect 21820 -2020 21890 -1950
rect 21930 -2020 22000 -1950
rect 24740 -3120 24810 -3050
rect 24850 -3120 24920 -3050
rect 24960 -3120 25030 -3050
rect 24740 -3230 24810 -3160
rect 24850 -3230 24920 -3160
rect 24960 -3230 25030 -3160
rect 24740 -3340 24810 -3270
rect 24850 -3340 24920 -3270
rect 24960 -3340 25030 -3270
rect 22470 -3760 22540 -3690
rect 22580 -3760 22650 -3690
rect 22690 -3760 22760 -3690
rect 22800 -3760 22870 -3690
rect 7310 -3950 7380 -3880
rect 7420 -3950 7490 -3880
rect 7530 -3950 7600 -3880
rect 22470 -3870 22540 -3800
rect 22580 -3870 22650 -3800
rect 22690 -3870 22760 -3800
rect 22800 -3870 22870 -3800
rect 26950 -3760 27020 -3690
rect 27060 -3760 27130 -3690
rect 27170 -3760 27240 -3690
rect 27280 -3760 27350 -3690
rect 26950 -3870 27020 -3800
rect 27060 -3870 27130 -3800
rect 27170 -3870 27240 -3800
rect 27280 -3870 27350 -3800
rect 7310 -4060 7380 -3990
rect 7420 -4060 7490 -3990
rect 7530 -4060 7600 -3990
rect 7310 -4170 7380 -4100
rect 7420 -4170 7490 -4100
rect 7530 -4170 7600 -4100
rect -1330 -4420 -1260 -4350
rect -1220 -4420 -1150 -4350
rect -1110 -4420 -1040 -4350
rect -1000 -4420 -930 -4350
rect -1330 -4530 -1260 -4460
rect -1220 -4530 -1150 -4460
rect -1110 -4530 -1040 -4460
rect -1000 -4530 -930 -4460
rect -560 -4360 -490 -4290
rect -450 -4360 -380 -4290
rect -340 -4360 -270 -4290
rect -230 -4360 -160 -4290
rect -560 -4470 -490 -4400
rect -450 -4470 -380 -4400
rect -340 -4470 -270 -4400
rect -230 -4470 -160 -4400
rect 14940 -4360 15010 -4290
rect 15050 -4360 15120 -4290
rect 15160 -4360 15230 -4290
rect 15270 -4360 15340 -4290
rect 14940 -4470 15010 -4400
rect 15050 -4470 15120 -4400
rect 15160 -4470 15230 -4400
rect 15270 -4470 15340 -4400
rect 15710 -4420 15780 -4350
rect 15820 -4420 15890 -4350
rect 15930 -4420 16000 -4350
rect 16040 -4420 16110 -4350
rect 15710 -4530 15780 -4460
rect 15820 -4530 15890 -4460
rect 15930 -4530 16000 -4460
rect 16040 -4530 16110 -4460
rect -1710 -6590 -1640 -6520
rect -1710 -6700 -1640 -6630
rect 7050 -6520 7110 -6460
rect 7150 -6520 7210 -6460
rect 7250 -6520 7310 -6460
rect 7050 -6620 7110 -6560
rect 7150 -6620 7210 -6560
rect 7250 -6620 7310 -6560
rect -1710 -6810 -1640 -6740
rect -1710 -6920 -1640 -6850
rect 4770 -6730 4830 -6670
rect 4870 -6730 4930 -6670
rect 4970 -6730 5030 -6670
rect 4770 -6830 4830 -6770
rect 4870 -6830 4930 -6770
rect 4970 -6830 5030 -6770
rect 7050 -6720 7110 -6660
rect 7150 -6720 7210 -6660
rect 7250 -6720 7310 -6660
rect 7050 -6820 7110 -6760
rect 7150 -6820 7210 -6760
rect 7250 -6820 7310 -6760
rect 7590 -6520 7650 -6460
rect 7690 -6520 7750 -6460
rect 7790 -6520 7850 -6460
rect 7590 -6620 7650 -6560
rect 7690 -6620 7750 -6560
rect 7790 -6620 7850 -6560
rect 16420 -6590 16490 -6520
rect 7590 -6720 7650 -6660
rect 7690 -6720 7750 -6660
rect 7790 -6720 7850 -6660
rect 7590 -6820 7650 -6760
rect 7690 -6820 7750 -6760
rect 7790 -6820 7850 -6760
rect 9870 -6730 9930 -6670
rect 9970 -6730 10030 -6670
rect 10070 -6730 10130 -6670
rect 9870 -6830 9930 -6770
rect 9970 -6830 10030 -6770
rect 10070 -6830 10130 -6770
rect 4770 -6930 4830 -6870
rect 4870 -6930 4930 -6870
rect 4970 -6930 5030 -6870
rect 9870 -6930 9930 -6870
rect 9970 -6930 10030 -6870
rect 10070 -6930 10130 -6870
rect 16420 -6700 16490 -6630
rect 16420 -6810 16490 -6740
rect 16420 -6920 16490 -6850
rect 20 -8210 90 -8140
rect 130 -8210 200 -8140
rect 230 -8210 300 -8140
rect 20 -8320 90 -8250
rect 130 -8320 200 -8250
rect 230 -8320 300 -8250
rect 20 -8430 90 -8360
rect 130 -8430 200 -8360
rect 230 -8430 300 -8360
rect 14600 -8300 14670 -8230
rect 14700 -8300 14770 -8230
rect 14810 -8300 14880 -8230
rect 14600 -8410 14670 -8340
rect 14700 -8410 14770 -8340
rect 14810 -8410 14880 -8340
rect 14600 -8520 14670 -8450
rect 14700 -8520 14770 -8450
rect 14810 -8520 14880 -8450
rect 21630 -8430 21700 -8360
rect 21730 -8430 21800 -8360
rect 21830 -8430 21900 -8360
rect 21630 -8530 21700 -8460
rect 21730 -8530 21800 -8460
rect 21830 -8530 21900 -8460
rect 21630 -8630 21700 -8560
rect 21730 -8630 21800 -8560
rect 21830 -8630 21900 -8560
rect 22650 -9080 22720 -9010
rect 22750 -9080 22820 -9010
rect 22850 -9080 22920 -9010
rect 22650 -9180 22720 -9110
rect 22750 -9180 22820 -9110
rect 22850 -9180 22920 -9110
rect 22650 -9280 22720 -9210
rect 22750 -9280 22820 -9210
rect 22850 -9280 22920 -9210
rect -240 -9730 -170 -9660
rect -130 -9730 -60 -9660
rect -20 -9730 50 -9660
rect 90 -9730 160 -9660
rect -240 -9860 -170 -9790
rect -130 -9860 -60 -9790
rect -20 -9860 50 -9790
rect 90 -9860 160 -9790
rect 14720 -9730 14790 -9660
rect 14830 -9730 14900 -9660
rect 14940 -9730 15010 -9660
rect 15050 -9730 15120 -9660
rect 14720 -9860 14790 -9790
rect 14830 -9860 14900 -9790
rect 14940 -9860 15010 -9790
rect 15050 -9860 15120 -9790
rect 1150 -10410 1220 -10340
rect 1260 -10410 1330 -10340
rect 1370 -10410 1440 -10340
rect 1480 -10410 1550 -10340
rect 1590 -10410 1660 -10340
rect 1700 -10410 1770 -10340
rect 1810 -10410 1880 -10340
rect 1920 -10410 1990 -10340
rect 2030 -10410 2100 -10340
rect 2140 -10410 2210 -10340
rect 2250 -10410 2320 -10340
rect 2360 -10410 2430 -10340
rect 2470 -10410 2540 -10340
rect 2580 -10410 2650 -10340
rect 1150 -10520 1220 -10450
rect 1260 -10520 1330 -10450
rect 1370 -10520 1440 -10450
rect 1480 -10520 1550 -10450
rect 1590 -10520 1660 -10450
rect 1700 -10520 1770 -10450
rect 1810 -10520 1880 -10450
rect 1920 -10520 1990 -10450
rect 2030 -10520 2100 -10450
rect 2140 -10520 2210 -10450
rect 2250 -10520 2320 -10450
rect 2360 -10520 2430 -10450
rect 2470 -10520 2540 -10450
rect 2580 -10520 2650 -10450
rect 12290 -10440 12360 -10370
rect 12400 -10440 12470 -10370
rect 12510 -10440 12580 -10370
rect 12620 -10440 12690 -10370
rect 12730 -10440 12800 -10370
rect 12840 -10440 12910 -10370
rect 12950 -10440 13020 -10370
rect 13060 -10440 13130 -10370
rect 13170 -10440 13240 -10370
rect 13280 -10440 13350 -10370
rect 13390 -10440 13460 -10370
rect 13500 -10440 13570 -10370
rect 13610 -10440 13680 -10370
rect 13720 -10440 13790 -10370
rect 12290 -10550 12360 -10480
rect 12400 -10550 12470 -10480
rect 12510 -10550 12580 -10480
rect 12620 -10550 12690 -10480
rect 12730 -10550 12800 -10480
rect 12840 -10550 12910 -10480
rect 12950 -10550 13020 -10480
rect 13060 -10550 13130 -10480
rect 13170 -10550 13240 -10480
rect 13280 -10550 13350 -10480
rect 13390 -10550 13460 -10480
rect 13500 -10550 13570 -10480
rect 13610 -10550 13680 -10480
rect 13720 -10550 13790 -10480
rect 1540 -12370 1610 -12300
rect 1650 -12370 1720 -12300
rect 1760 -12370 1830 -12300
rect 1870 -12370 1940 -12300
rect 1980 -12370 2050 -12300
rect 2090 -12370 2160 -12300
rect 2200 -12370 2270 -12300
rect 2310 -12370 2380 -12300
rect 2420 -12370 2490 -12300
rect 2530 -12370 2600 -12300
rect 2640 -12370 2710 -12300
rect 2750 -12370 2820 -12300
rect 2860 -12370 2930 -12300
rect 2970 -12370 3040 -12300
rect 1540 -12480 1610 -12410
rect 1650 -12480 1720 -12410
rect 1760 -12480 1830 -12410
rect 1870 -12480 1940 -12410
rect 1980 -12480 2050 -12410
rect 2090 -12480 2160 -12410
rect 2200 -12480 2270 -12410
rect 2310 -12480 2380 -12410
rect 2420 -12480 2490 -12410
rect 2530 -12480 2600 -12410
rect 2640 -12480 2710 -12410
rect 2750 -12480 2820 -12410
rect 2860 -12480 2930 -12410
rect 2970 -12480 3040 -12410
rect 11820 -12370 11890 -12300
rect 11930 -12370 12000 -12300
rect 12040 -12370 12110 -12300
rect 12150 -12370 12220 -12300
rect 12260 -12370 12330 -12300
rect 12370 -12370 12440 -12300
rect 12480 -12370 12550 -12300
rect 12590 -12370 12660 -12300
rect 12700 -12370 12770 -12300
rect 12810 -12370 12880 -12300
rect 12920 -12370 12990 -12300
rect 13030 -12370 13100 -12300
rect 13140 -12370 13210 -12300
rect 13250 -12370 13320 -12300
rect 11820 -12480 11890 -12410
rect 11930 -12480 12000 -12410
rect 12040 -12480 12110 -12410
rect 12150 -12480 12220 -12410
rect 12260 -12480 12330 -12410
rect 12370 -12480 12440 -12410
rect 12480 -12480 12550 -12410
rect 12590 -12480 12660 -12410
rect 12700 -12480 12770 -12410
rect 12810 -12480 12880 -12410
rect 12920 -12480 12990 -12410
rect 13030 -12480 13100 -12410
rect 13140 -12480 13210 -12410
rect 13250 -12480 13320 -12410
rect 6310 -13310 6370 -13250
rect 6410 -13310 6470 -13250
rect 6510 -13310 6570 -13250
rect 6310 -13400 6370 -13340
rect 6410 -13400 6470 -13340
rect 6510 -13400 6570 -13340
rect 6310 -13490 6370 -13430
rect 6410 -13490 6470 -13430
rect 6510 -13490 6570 -13430
rect 6310 -13590 6370 -13530
rect 6410 -13590 6470 -13530
rect 6510 -13590 6570 -13530
rect 6310 -13680 6370 -13620
rect 6410 -13680 6470 -13620
rect 6510 -13680 6570 -13620
rect 6310 -13770 6370 -13710
rect 6410 -13770 6470 -13710
rect 6510 -13770 6570 -13710
rect 8330 -13310 8390 -13250
rect 8430 -13310 8490 -13250
rect 8530 -13310 8590 -13250
rect 8330 -13400 8390 -13340
rect 8430 -13400 8490 -13340
rect 8530 -13400 8590 -13340
rect 8330 -13490 8390 -13430
rect 8430 -13490 8490 -13430
rect 8530 -13490 8590 -13430
rect 8330 -13590 8390 -13530
rect 8430 -13590 8490 -13530
rect 8530 -13590 8590 -13530
rect 8330 -13680 8390 -13620
rect 8430 -13680 8490 -13620
rect 8530 -13680 8590 -13620
rect 8330 -13770 8390 -13710
rect 8430 -13770 8490 -13710
rect 8530 -13770 8590 -13710
rect 21630 -14090 21700 -14020
rect 21730 -14090 21800 -14020
rect 21830 -14090 21900 -14020
rect 21630 -14190 21700 -14120
rect 21730 -14190 21800 -14120
rect 21830 -14190 21900 -14120
rect 21630 -14290 21700 -14220
rect 21730 -14290 21800 -14220
rect 21830 -14290 21900 -14220
rect 22920 -14940 22990 -14870
rect 23020 -14940 23090 -14870
rect 23120 -14940 23190 -14870
rect 22920 -15040 22990 -14970
rect 23020 -15040 23090 -14970
rect 23120 -15040 23190 -14970
rect 22920 -15140 22990 -15070
rect 23020 -15140 23090 -15070
rect 23120 -15140 23190 -15070
rect 4980 -17160 5040 -17100
rect 5080 -17160 5140 -17100
rect 5180 -17160 5240 -17100
rect 4980 -17260 5040 -17200
rect 5080 -17260 5140 -17200
rect 5180 -17260 5240 -17200
rect 4980 -17360 5040 -17300
rect 5080 -17360 5140 -17300
rect 5180 -17360 5240 -17300
rect 9660 -17160 9720 -17100
rect 9760 -17160 9820 -17100
rect 9860 -17160 9920 -17100
rect 9660 -17260 9720 -17200
rect 9760 -17260 9820 -17200
rect 9860 -17260 9920 -17200
rect 9660 -17360 9720 -17300
rect 9760 -17360 9820 -17300
rect 9860 -17360 9920 -17300
rect 6460 -17820 6530 -17750
rect 6560 -17820 6630 -17750
rect 6660 -17820 6730 -17750
rect 6460 -17930 6530 -17860
rect 6560 -17930 6630 -17860
rect 6660 -17930 6730 -17860
rect 6460 -18040 6530 -17970
rect 6560 -18040 6630 -17970
rect 6660 -18040 6730 -17970
rect 6460 -18150 6530 -18080
rect 6560 -18150 6630 -18080
rect 6660 -18150 6730 -18080
rect 8170 -17820 8240 -17750
rect 8270 -17820 8340 -17750
rect 8370 -17820 8440 -17750
rect 8170 -17930 8240 -17860
rect 8270 -17930 8340 -17860
rect 8370 -17930 8440 -17860
rect 8170 -18040 8240 -17970
rect 8270 -18040 8340 -17970
rect 8370 -18040 8440 -17970
rect 8170 -18150 8240 -18080
rect 8270 -18150 8340 -18080
rect 8370 -18150 8440 -18080
rect 21630 -20170 21700 -20100
rect 21730 -20170 21800 -20100
rect 21830 -20170 21900 -20100
rect 21630 -20270 21700 -20200
rect 21730 -20270 21800 -20200
rect 21830 -20270 21900 -20200
rect 21630 -20370 21700 -20300
rect 21730 -20370 21800 -20300
rect 21830 -20370 21900 -20300
rect 22700 -20800 22770 -20730
rect 22800 -20800 22870 -20730
rect 22900 -20800 22970 -20730
rect 22700 -20900 22770 -20830
rect 22800 -20900 22870 -20830
rect 22900 -20900 22970 -20830
rect 22700 -21000 22770 -20930
rect 22800 -21000 22870 -20930
rect 22900 -21000 22970 -20930
rect 1620 -22730 1690 -22660
rect 1730 -22730 1800 -22660
rect 1840 -22730 1910 -22660
rect 1950 -22730 2020 -22660
rect 2060 -22730 2130 -22660
rect 2170 -22730 2240 -22660
rect 2280 -22730 2350 -22660
rect 2390 -22730 2460 -22660
rect 2500 -22730 2570 -22660
rect 2610 -22730 2680 -22660
rect 2720 -22730 2790 -22660
rect 2830 -22730 2900 -22660
rect 2940 -22730 3010 -22660
rect 3050 -22730 3120 -22660
rect 1620 -22840 1690 -22770
rect 1730 -22840 1800 -22770
rect 1840 -22840 1910 -22770
rect 1950 -22840 2020 -22770
rect 2060 -22840 2130 -22770
rect 2170 -22840 2240 -22770
rect 2280 -22840 2350 -22770
rect 2390 -22840 2460 -22770
rect 2500 -22840 2570 -22770
rect 2610 -22840 2680 -22770
rect 2720 -22840 2790 -22770
rect 2830 -22840 2900 -22770
rect 2940 -22840 3010 -22770
rect 3050 -22840 3120 -22770
rect 11820 -22730 11890 -22660
rect 11930 -22730 12000 -22660
rect 12040 -22730 12110 -22660
rect 12150 -22730 12220 -22660
rect 12260 -22730 12330 -22660
rect 12370 -22730 12440 -22660
rect 12480 -22730 12550 -22660
rect 12590 -22730 12660 -22660
rect 12700 -22730 12770 -22660
rect 12810 -22730 12880 -22660
rect 12920 -22730 12990 -22660
rect 13030 -22730 13100 -22660
rect 13140 -22730 13210 -22660
rect 13250 -22730 13320 -22660
rect 11820 -22840 11890 -22770
rect 11930 -22840 12000 -22770
rect 12040 -22840 12110 -22770
rect 12150 -22840 12220 -22770
rect 12260 -22840 12330 -22770
rect 12370 -22840 12440 -22770
rect 12480 -22840 12550 -22770
rect 12590 -22840 12660 -22770
rect 12700 -22840 12770 -22770
rect 12810 -22840 12880 -22770
rect 12920 -22840 12990 -22770
rect 13030 -22840 13100 -22770
rect 13140 -22840 13210 -22770
rect 13250 -22840 13320 -22770
<< metal3 >>
rect -5550 21580 6760 21640
rect -5550 21510 -5260 21580
rect -5190 21510 -5170 21580
rect -5100 21510 -5080 21580
rect -5010 21510 -4990 21580
rect -4920 21510 -4900 21580
rect -4830 21510 -4810 21580
rect -4740 21510 -4720 21580
rect -4650 21510 -4630 21580
rect -4560 21510 -4540 21580
rect -4470 21510 -4450 21580
rect -4380 21510 -4360 21580
rect -4290 21510 -4270 21580
rect -4200 21510 -4180 21580
rect -4110 21510 -4090 21580
rect -4020 21510 -4000 21580
rect -3930 21510 -3910 21580
rect -3840 21510 -3820 21580
rect -3750 21510 -3730 21580
rect -3660 21510 -3640 21580
rect -3570 21510 -3550 21580
rect -3480 21510 -3460 21580
rect -3390 21510 -3370 21580
rect -3300 21510 -3280 21580
rect -3210 21510 -3190 21580
rect -3120 21510 -3100 21580
rect -3030 21510 -3010 21580
rect -2940 21510 -2920 21580
rect -2850 21510 -2830 21580
rect -2760 21510 -2740 21580
rect -2670 21510 -2650 21580
rect -2580 21510 -2560 21580
rect -2490 21510 -2470 21580
rect -2400 21510 -2380 21580
rect -2310 21510 -2250 21580
rect -2180 21510 -2160 21580
rect -2090 21510 -2070 21580
rect -2000 21510 -1980 21580
rect -1910 21510 -1890 21580
rect -1820 21510 -1800 21580
rect -1730 21510 -1710 21580
rect -1640 21510 -1620 21580
rect -1550 21510 -1530 21580
rect -1460 21510 -1440 21580
rect -1370 21510 -1350 21580
rect -1280 21510 -1260 21580
rect -1190 21510 -1170 21580
rect -1100 21510 -1080 21580
rect -1010 21510 -990 21580
rect -920 21510 -900 21580
rect -830 21510 -810 21580
rect -740 21510 -720 21580
rect -650 21510 -630 21580
rect -560 21510 -540 21580
rect -470 21510 -450 21580
rect -380 21510 -360 21580
rect -290 21510 -270 21580
rect -200 21510 -180 21580
rect -110 21510 -90 21580
rect -20 21510 0 21580
rect 70 21510 90 21580
rect 160 21510 180 21580
rect 250 21510 270 21580
rect 340 21510 360 21580
rect 430 21510 450 21580
rect 520 21510 540 21580
rect 610 21510 630 21580
rect 700 21510 760 21580
rect 830 21510 850 21580
rect 920 21510 940 21580
rect 1010 21510 1030 21580
rect 1100 21510 1120 21580
rect 1190 21510 1210 21580
rect 1280 21510 1300 21580
rect 1370 21510 1390 21580
rect 1460 21510 1480 21580
rect 1550 21510 1570 21580
rect 1640 21510 1660 21580
rect 1730 21510 1750 21580
rect 1820 21510 1840 21580
rect 1910 21510 1930 21580
rect 2000 21510 2020 21580
rect 2090 21510 2110 21580
rect 2180 21510 2200 21580
rect 2270 21510 2290 21580
rect 2360 21510 2380 21580
rect 2450 21510 2470 21580
rect 2540 21510 2560 21580
rect 2630 21510 2650 21580
rect 2720 21510 2740 21580
rect 2810 21510 2830 21580
rect 2900 21510 2920 21580
rect 2990 21510 3010 21580
rect 3080 21510 3100 21580
rect 3170 21510 3190 21580
rect 3260 21510 3280 21580
rect 3350 21510 3370 21580
rect 3440 21510 3460 21580
rect 3530 21510 3550 21580
rect 3620 21510 3640 21580
rect 3710 21510 3770 21580
rect 3840 21510 3860 21580
rect 3930 21510 3950 21580
rect 4020 21510 4040 21580
rect 4110 21510 4130 21580
rect 4200 21510 4220 21580
rect 4290 21510 4310 21580
rect 4380 21510 4400 21580
rect 4470 21510 4490 21580
rect 4560 21510 4580 21580
rect 4650 21510 4670 21580
rect 4740 21510 4760 21580
rect 4830 21510 4850 21580
rect 4920 21510 4940 21580
rect 5010 21510 5030 21580
rect 5100 21510 5120 21580
rect 5190 21510 5210 21580
rect 5280 21510 5300 21580
rect 5370 21510 5390 21580
rect 5460 21510 5480 21580
rect 5550 21510 5570 21580
rect 5640 21510 5660 21580
rect 5730 21510 5750 21580
rect 5820 21510 5840 21580
rect 5910 21510 5930 21580
rect 6000 21510 6020 21580
rect 6090 21510 6110 21580
rect 6180 21510 6200 21580
rect 6270 21510 6290 21580
rect 6360 21510 6380 21580
rect 6450 21510 6470 21580
rect 6540 21510 6560 21580
rect 6630 21510 6650 21580
rect 6720 21510 6760 21580
rect -5550 21490 6760 21510
rect -5550 21420 -5260 21490
rect -5190 21420 -5170 21490
rect -5100 21420 -5080 21490
rect -5010 21420 -4990 21490
rect -4920 21420 -4900 21490
rect -4830 21420 -4810 21490
rect -4740 21420 -4720 21490
rect -4650 21420 -4630 21490
rect -4560 21420 -4540 21490
rect -4470 21420 -4450 21490
rect -4380 21420 -4360 21490
rect -4290 21420 -4270 21490
rect -4200 21420 -4180 21490
rect -4110 21420 -4090 21490
rect -4020 21420 -4000 21490
rect -3930 21420 -3910 21490
rect -3840 21420 -3820 21490
rect -3750 21420 -3730 21490
rect -3660 21420 -3640 21490
rect -3570 21420 -3550 21490
rect -3480 21420 -3460 21490
rect -3390 21420 -3370 21490
rect -3300 21420 -3280 21490
rect -3210 21420 -3190 21490
rect -3120 21420 -3100 21490
rect -3030 21420 -3010 21490
rect -2940 21420 -2920 21490
rect -2850 21420 -2830 21490
rect -2760 21420 -2740 21490
rect -2670 21420 -2650 21490
rect -2580 21420 -2560 21490
rect -2490 21420 -2470 21490
rect -2400 21420 -2380 21490
rect -2310 21420 -2250 21490
rect -2180 21420 -2160 21490
rect -2090 21420 -2070 21490
rect -2000 21420 -1980 21490
rect -1910 21420 -1890 21490
rect -1820 21420 -1800 21490
rect -1730 21420 -1710 21490
rect -1640 21420 -1620 21490
rect -1550 21420 -1530 21490
rect -1460 21420 -1440 21490
rect -1370 21420 -1350 21490
rect -1280 21420 -1260 21490
rect -1190 21420 -1170 21490
rect -1100 21420 -1080 21490
rect -1010 21420 -990 21490
rect -920 21420 -900 21490
rect -830 21420 -810 21490
rect -740 21420 -720 21490
rect -650 21420 -630 21490
rect -560 21420 -540 21490
rect -470 21420 -450 21490
rect -380 21420 -360 21490
rect -290 21420 -270 21490
rect -200 21420 -180 21490
rect -110 21420 -90 21490
rect -20 21420 0 21490
rect 70 21420 90 21490
rect 160 21420 180 21490
rect 250 21420 270 21490
rect 340 21420 360 21490
rect 430 21420 450 21490
rect 520 21420 540 21490
rect 610 21420 630 21490
rect 700 21420 760 21490
rect 830 21420 850 21490
rect 920 21420 940 21490
rect 1010 21420 1030 21490
rect 1100 21420 1120 21490
rect 1190 21420 1210 21490
rect 1280 21420 1300 21490
rect 1370 21420 1390 21490
rect 1460 21420 1480 21490
rect 1550 21420 1570 21490
rect 1640 21420 1660 21490
rect 1730 21420 1750 21490
rect 1820 21420 1840 21490
rect 1910 21420 1930 21490
rect 2000 21420 2020 21490
rect 2090 21420 2110 21490
rect 2180 21420 2200 21490
rect 2270 21420 2290 21490
rect 2360 21420 2380 21490
rect 2450 21420 2470 21490
rect 2540 21420 2560 21490
rect 2630 21420 2650 21490
rect 2720 21420 2740 21490
rect 2810 21420 2830 21490
rect 2900 21420 2920 21490
rect 2990 21420 3010 21490
rect 3080 21420 3100 21490
rect 3170 21420 3190 21490
rect 3260 21420 3280 21490
rect 3350 21420 3370 21490
rect 3440 21420 3460 21490
rect 3530 21420 3550 21490
rect 3620 21420 3640 21490
rect 3710 21420 3770 21490
rect 3840 21420 3860 21490
rect 3930 21420 3950 21490
rect 4020 21420 4040 21490
rect 4110 21420 4130 21490
rect 4200 21420 4220 21490
rect 4290 21420 4310 21490
rect 4380 21420 4400 21490
rect 4470 21420 4490 21490
rect 4560 21420 4580 21490
rect 4650 21420 4670 21490
rect 4740 21420 4760 21490
rect 4830 21420 4850 21490
rect 4920 21420 4940 21490
rect 5010 21420 5030 21490
rect 5100 21420 5120 21490
rect 5190 21420 5210 21490
rect 5280 21420 5300 21490
rect 5370 21420 5390 21490
rect 5460 21420 5480 21490
rect 5550 21420 5570 21490
rect 5640 21420 5660 21490
rect 5730 21420 5750 21490
rect 5820 21420 5840 21490
rect 5910 21420 5930 21490
rect 6000 21420 6020 21490
rect 6090 21420 6110 21490
rect 6180 21420 6200 21490
rect 6270 21420 6290 21490
rect 6360 21420 6380 21490
rect 6450 21420 6470 21490
rect 6540 21420 6560 21490
rect 6630 21420 6650 21490
rect 6720 21420 6760 21490
rect -5550 21400 6760 21420
rect -5550 21330 -5260 21400
rect -5190 21330 -5170 21400
rect -5100 21330 -5080 21400
rect -5010 21330 -4990 21400
rect -4920 21330 -4900 21400
rect -4830 21330 -4810 21400
rect -4740 21330 -4720 21400
rect -4650 21330 -4630 21400
rect -4560 21330 -4540 21400
rect -4470 21330 -4450 21400
rect -4380 21330 -4360 21400
rect -4290 21330 -4270 21400
rect -4200 21330 -4180 21400
rect -4110 21330 -4090 21400
rect -4020 21330 -4000 21400
rect -3930 21330 -3910 21400
rect -3840 21330 -3820 21400
rect -3750 21330 -3730 21400
rect -3660 21330 -3640 21400
rect -3570 21330 -3550 21400
rect -3480 21330 -3460 21400
rect -3390 21330 -3370 21400
rect -3300 21330 -3280 21400
rect -3210 21330 -3190 21400
rect -3120 21330 -3100 21400
rect -3030 21330 -3010 21400
rect -2940 21330 -2920 21400
rect -2850 21330 -2830 21400
rect -2760 21330 -2740 21400
rect -2670 21330 -2650 21400
rect -2580 21330 -2560 21400
rect -2490 21330 -2470 21400
rect -2400 21330 -2380 21400
rect -2310 21330 -2250 21400
rect -2180 21330 -2160 21400
rect -2090 21330 -2070 21400
rect -2000 21330 -1980 21400
rect -1910 21330 -1890 21400
rect -1820 21330 -1800 21400
rect -1730 21330 -1710 21400
rect -1640 21330 -1620 21400
rect -1550 21330 -1530 21400
rect -1460 21330 -1440 21400
rect -1370 21330 -1350 21400
rect -1280 21330 -1260 21400
rect -1190 21330 -1170 21400
rect -1100 21330 -1080 21400
rect -1010 21330 -990 21400
rect -920 21330 -900 21400
rect -830 21330 -810 21400
rect -740 21330 -720 21400
rect -650 21330 -630 21400
rect -560 21330 -540 21400
rect -470 21330 -450 21400
rect -380 21330 -360 21400
rect -290 21330 -270 21400
rect -200 21330 -180 21400
rect -110 21330 -90 21400
rect -20 21330 0 21400
rect 70 21330 90 21400
rect 160 21330 180 21400
rect 250 21330 270 21400
rect 340 21330 360 21400
rect 430 21330 450 21400
rect 520 21330 540 21400
rect 610 21330 630 21400
rect 700 21330 760 21400
rect 830 21330 850 21400
rect 920 21330 940 21400
rect 1010 21330 1030 21400
rect 1100 21330 1120 21400
rect 1190 21330 1210 21400
rect 1280 21330 1300 21400
rect 1370 21330 1390 21400
rect 1460 21330 1480 21400
rect 1550 21330 1570 21400
rect 1640 21330 1660 21400
rect 1730 21330 1750 21400
rect 1820 21330 1840 21400
rect 1910 21330 1930 21400
rect 2000 21330 2020 21400
rect 2090 21330 2110 21400
rect 2180 21330 2200 21400
rect 2270 21330 2290 21400
rect 2360 21330 2380 21400
rect 2450 21330 2470 21400
rect 2540 21330 2560 21400
rect 2630 21330 2650 21400
rect 2720 21330 2740 21400
rect 2810 21330 2830 21400
rect 2900 21330 2920 21400
rect 2990 21330 3010 21400
rect 3080 21330 3100 21400
rect 3170 21330 3190 21400
rect 3260 21330 3280 21400
rect 3350 21330 3370 21400
rect 3440 21330 3460 21400
rect 3530 21330 3550 21400
rect 3620 21330 3640 21400
rect 3710 21330 3770 21400
rect 3840 21330 3860 21400
rect 3930 21330 3950 21400
rect 4020 21330 4040 21400
rect 4110 21330 4130 21400
rect 4200 21330 4220 21400
rect 4290 21330 4310 21400
rect 4380 21330 4400 21400
rect 4470 21330 4490 21400
rect 4560 21330 4580 21400
rect 4650 21330 4670 21400
rect 4740 21330 4760 21400
rect 4830 21330 4850 21400
rect 4920 21330 4940 21400
rect 5010 21330 5030 21400
rect 5100 21330 5120 21400
rect 5190 21330 5210 21400
rect 5280 21330 5300 21400
rect 5370 21330 5390 21400
rect 5460 21330 5480 21400
rect 5550 21330 5570 21400
rect 5640 21330 5660 21400
rect 5730 21330 5750 21400
rect 5820 21330 5840 21400
rect 5910 21330 5930 21400
rect 6000 21330 6020 21400
rect 6090 21330 6110 21400
rect 6180 21330 6200 21400
rect 6270 21330 6290 21400
rect 6360 21330 6380 21400
rect 6450 21330 6470 21400
rect 6540 21330 6560 21400
rect 6630 21330 6650 21400
rect 6720 21330 6760 21400
rect -5550 8690 6760 21330
rect 8140 21580 20450 21640
rect 8140 21510 8180 21580
rect 8250 21510 8270 21580
rect 8340 21510 8360 21580
rect 8430 21510 8450 21580
rect 8520 21510 8540 21580
rect 8610 21510 8630 21580
rect 8700 21510 8720 21580
rect 8790 21510 8810 21580
rect 8880 21510 8900 21580
rect 8970 21510 8990 21580
rect 9060 21510 9080 21580
rect 9150 21510 9170 21580
rect 9240 21510 9260 21580
rect 9330 21510 9350 21580
rect 9420 21510 9440 21580
rect 9510 21510 9530 21580
rect 9600 21510 9620 21580
rect 9690 21510 9710 21580
rect 9780 21510 9800 21580
rect 9870 21510 9890 21580
rect 9960 21510 9980 21580
rect 10050 21510 10070 21580
rect 10140 21510 10160 21580
rect 10230 21510 10250 21580
rect 10320 21510 10340 21580
rect 10410 21510 10430 21580
rect 10500 21510 10520 21580
rect 10590 21510 10610 21580
rect 10680 21510 10700 21580
rect 10770 21510 10790 21580
rect 10860 21510 10880 21580
rect 10950 21510 10970 21580
rect 11040 21510 11060 21580
rect 11130 21510 11190 21580
rect 11260 21510 11280 21580
rect 11350 21510 11370 21580
rect 11440 21510 11460 21580
rect 11530 21510 11550 21580
rect 11620 21510 11640 21580
rect 11710 21510 11730 21580
rect 11800 21510 11820 21580
rect 11890 21510 11910 21580
rect 11980 21510 12000 21580
rect 12070 21510 12090 21580
rect 12160 21510 12180 21580
rect 12250 21510 12270 21580
rect 12340 21510 12360 21580
rect 12430 21510 12450 21580
rect 12520 21510 12540 21580
rect 12610 21510 12630 21580
rect 12700 21510 12720 21580
rect 12790 21510 12810 21580
rect 12880 21510 12900 21580
rect 12970 21510 12990 21580
rect 13060 21510 13080 21580
rect 13150 21510 13170 21580
rect 13240 21510 13260 21580
rect 13330 21510 13350 21580
rect 13420 21510 13440 21580
rect 13510 21510 13530 21580
rect 13600 21510 13620 21580
rect 13690 21510 13710 21580
rect 13780 21510 13800 21580
rect 13870 21510 13890 21580
rect 13960 21510 13980 21580
rect 14050 21510 14070 21580
rect 14140 21510 14200 21580
rect 14270 21510 14290 21580
rect 14360 21510 14380 21580
rect 14450 21510 14470 21580
rect 14540 21510 14560 21580
rect 14630 21510 14650 21580
rect 14720 21510 14740 21580
rect 14810 21510 14830 21580
rect 14900 21510 14920 21580
rect 14990 21510 15010 21580
rect 15080 21510 15100 21580
rect 15170 21510 15190 21580
rect 15260 21510 15280 21580
rect 15350 21510 15370 21580
rect 15440 21510 15460 21580
rect 15530 21510 15550 21580
rect 15620 21510 15640 21580
rect 15710 21510 15730 21580
rect 15800 21510 15820 21580
rect 15890 21510 15910 21580
rect 15980 21510 16000 21580
rect 16070 21510 16090 21580
rect 16160 21510 16180 21580
rect 16250 21510 16270 21580
rect 16340 21510 16360 21580
rect 16430 21510 16450 21580
rect 16520 21510 16540 21580
rect 16610 21510 16630 21580
rect 16700 21510 16720 21580
rect 16790 21510 16810 21580
rect 16880 21510 16900 21580
rect 16970 21510 16990 21580
rect 17060 21510 17080 21580
rect 17150 21510 17210 21580
rect 17280 21510 17300 21580
rect 17370 21510 17390 21580
rect 17460 21510 17480 21580
rect 17550 21510 17570 21580
rect 17640 21510 17660 21580
rect 17730 21510 17750 21580
rect 17820 21510 17840 21580
rect 17910 21510 17930 21580
rect 18000 21510 18020 21580
rect 18090 21510 18110 21580
rect 18180 21510 18200 21580
rect 18270 21510 18290 21580
rect 18360 21510 18380 21580
rect 18450 21510 18470 21580
rect 18540 21510 18560 21580
rect 18630 21510 18650 21580
rect 18720 21510 18740 21580
rect 18810 21510 18830 21580
rect 18900 21510 18920 21580
rect 18990 21510 19010 21580
rect 19080 21510 19100 21580
rect 19170 21510 19190 21580
rect 19260 21510 19280 21580
rect 19350 21510 19370 21580
rect 19440 21510 19460 21580
rect 19530 21510 19550 21580
rect 19620 21510 19640 21580
rect 19710 21510 19730 21580
rect 19800 21510 19820 21580
rect 19890 21510 19910 21580
rect 19980 21510 20000 21580
rect 20070 21510 20090 21580
rect 20160 21510 20450 21580
rect 8140 21490 20450 21510
rect 8140 21420 8180 21490
rect 8250 21420 8270 21490
rect 8340 21420 8360 21490
rect 8430 21420 8450 21490
rect 8520 21420 8540 21490
rect 8610 21420 8630 21490
rect 8700 21420 8720 21490
rect 8790 21420 8810 21490
rect 8880 21420 8900 21490
rect 8970 21420 8990 21490
rect 9060 21420 9080 21490
rect 9150 21420 9170 21490
rect 9240 21420 9260 21490
rect 9330 21420 9350 21490
rect 9420 21420 9440 21490
rect 9510 21420 9530 21490
rect 9600 21420 9620 21490
rect 9690 21420 9710 21490
rect 9780 21420 9800 21490
rect 9870 21420 9890 21490
rect 9960 21420 9980 21490
rect 10050 21420 10070 21490
rect 10140 21420 10160 21490
rect 10230 21420 10250 21490
rect 10320 21420 10340 21490
rect 10410 21420 10430 21490
rect 10500 21420 10520 21490
rect 10590 21420 10610 21490
rect 10680 21420 10700 21490
rect 10770 21420 10790 21490
rect 10860 21420 10880 21490
rect 10950 21420 10970 21490
rect 11040 21420 11060 21490
rect 11130 21420 11190 21490
rect 11260 21420 11280 21490
rect 11350 21420 11370 21490
rect 11440 21420 11460 21490
rect 11530 21420 11550 21490
rect 11620 21420 11640 21490
rect 11710 21420 11730 21490
rect 11800 21420 11820 21490
rect 11890 21420 11910 21490
rect 11980 21420 12000 21490
rect 12070 21420 12090 21490
rect 12160 21420 12180 21490
rect 12250 21420 12270 21490
rect 12340 21420 12360 21490
rect 12430 21420 12450 21490
rect 12520 21420 12540 21490
rect 12610 21420 12630 21490
rect 12700 21420 12720 21490
rect 12790 21420 12810 21490
rect 12880 21420 12900 21490
rect 12970 21420 12990 21490
rect 13060 21420 13080 21490
rect 13150 21420 13170 21490
rect 13240 21420 13260 21490
rect 13330 21420 13350 21490
rect 13420 21420 13440 21490
rect 13510 21420 13530 21490
rect 13600 21420 13620 21490
rect 13690 21420 13710 21490
rect 13780 21420 13800 21490
rect 13870 21420 13890 21490
rect 13960 21420 13980 21490
rect 14050 21420 14070 21490
rect 14140 21420 14200 21490
rect 14270 21420 14290 21490
rect 14360 21420 14380 21490
rect 14450 21420 14470 21490
rect 14540 21420 14560 21490
rect 14630 21420 14650 21490
rect 14720 21420 14740 21490
rect 14810 21420 14830 21490
rect 14900 21420 14920 21490
rect 14990 21420 15010 21490
rect 15080 21420 15100 21490
rect 15170 21420 15190 21490
rect 15260 21420 15280 21490
rect 15350 21420 15370 21490
rect 15440 21420 15460 21490
rect 15530 21420 15550 21490
rect 15620 21420 15640 21490
rect 15710 21420 15730 21490
rect 15800 21420 15820 21490
rect 15890 21420 15910 21490
rect 15980 21420 16000 21490
rect 16070 21420 16090 21490
rect 16160 21420 16180 21490
rect 16250 21420 16270 21490
rect 16340 21420 16360 21490
rect 16430 21420 16450 21490
rect 16520 21420 16540 21490
rect 16610 21420 16630 21490
rect 16700 21420 16720 21490
rect 16790 21420 16810 21490
rect 16880 21420 16900 21490
rect 16970 21420 16990 21490
rect 17060 21420 17080 21490
rect 17150 21420 17210 21490
rect 17280 21420 17300 21490
rect 17370 21420 17390 21490
rect 17460 21420 17480 21490
rect 17550 21420 17570 21490
rect 17640 21420 17660 21490
rect 17730 21420 17750 21490
rect 17820 21420 17840 21490
rect 17910 21420 17930 21490
rect 18000 21420 18020 21490
rect 18090 21420 18110 21490
rect 18180 21420 18200 21490
rect 18270 21420 18290 21490
rect 18360 21420 18380 21490
rect 18450 21420 18470 21490
rect 18540 21420 18560 21490
rect 18630 21420 18650 21490
rect 18720 21420 18740 21490
rect 18810 21420 18830 21490
rect 18900 21420 18920 21490
rect 18990 21420 19010 21490
rect 19080 21420 19100 21490
rect 19170 21420 19190 21490
rect 19260 21420 19280 21490
rect 19350 21420 19370 21490
rect 19440 21420 19460 21490
rect 19530 21420 19550 21490
rect 19620 21420 19640 21490
rect 19710 21420 19730 21490
rect 19800 21420 19820 21490
rect 19890 21420 19910 21490
rect 19980 21420 20000 21490
rect 20070 21420 20090 21490
rect 20160 21420 20450 21490
rect 8140 21400 20450 21420
rect 8140 21330 8180 21400
rect 8250 21330 8270 21400
rect 8340 21330 8360 21400
rect 8430 21330 8450 21400
rect 8520 21330 8540 21400
rect 8610 21330 8630 21400
rect 8700 21330 8720 21400
rect 8790 21330 8810 21400
rect 8880 21330 8900 21400
rect 8970 21330 8990 21400
rect 9060 21330 9080 21400
rect 9150 21330 9170 21400
rect 9240 21330 9260 21400
rect 9330 21330 9350 21400
rect 9420 21330 9440 21400
rect 9510 21330 9530 21400
rect 9600 21330 9620 21400
rect 9690 21330 9710 21400
rect 9780 21330 9800 21400
rect 9870 21330 9890 21400
rect 9960 21330 9980 21400
rect 10050 21330 10070 21400
rect 10140 21330 10160 21400
rect 10230 21330 10250 21400
rect 10320 21330 10340 21400
rect 10410 21330 10430 21400
rect 10500 21330 10520 21400
rect 10590 21330 10610 21400
rect 10680 21330 10700 21400
rect 10770 21330 10790 21400
rect 10860 21330 10880 21400
rect 10950 21330 10970 21400
rect 11040 21330 11060 21400
rect 11130 21330 11190 21400
rect 11260 21330 11280 21400
rect 11350 21330 11370 21400
rect 11440 21330 11460 21400
rect 11530 21330 11550 21400
rect 11620 21330 11640 21400
rect 11710 21330 11730 21400
rect 11800 21330 11820 21400
rect 11890 21330 11910 21400
rect 11980 21330 12000 21400
rect 12070 21330 12090 21400
rect 12160 21330 12180 21400
rect 12250 21330 12270 21400
rect 12340 21330 12360 21400
rect 12430 21330 12450 21400
rect 12520 21330 12540 21400
rect 12610 21330 12630 21400
rect 12700 21330 12720 21400
rect 12790 21330 12810 21400
rect 12880 21330 12900 21400
rect 12970 21330 12990 21400
rect 13060 21330 13080 21400
rect 13150 21330 13170 21400
rect 13240 21330 13260 21400
rect 13330 21330 13350 21400
rect 13420 21330 13440 21400
rect 13510 21330 13530 21400
rect 13600 21330 13620 21400
rect 13690 21330 13710 21400
rect 13780 21330 13800 21400
rect 13870 21330 13890 21400
rect 13960 21330 13980 21400
rect 14050 21330 14070 21400
rect 14140 21330 14200 21400
rect 14270 21330 14290 21400
rect 14360 21330 14380 21400
rect 14450 21330 14470 21400
rect 14540 21330 14560 21400
rect 14630 21330 14650 21400
rect 14720 21330 14740 21400
rect 14810 21330 14830 21400
rect 14900 21330 14920 21400
rect 14990 21330 15010 21400
rect 15080 21330 15100 21400
rect 15170 21330 15190 21400
rect 15260 21330 15280 21400
rect 15350 21330 15370 21400
rect 15440 21330 15460 21400
rect 15530 21330 15550 21400
rect 15620 21330 15640 21400
rect 15710 21330 15730 21400
rect 15800 21330 15820 21400
rect 15890 21330 15910 21400
rect 15980 21330 16000 21400
rect 16070 21330 16090 21400
rect 16160 21330 16180 21400
rect 16250 21330 16270 21400
rect 16340 21330 16360 21400
rect 16430 21330 16450 21400
rect 16520 21330 16540 21400
rect 16610 21330 16630 21400
rect 16700 21330 16720 21400
rect 16790 21330 16810 21400
rect 16880 21330 16900 21400
rect 16970 21330 16990 21400
rect 17060 21330 17080 21400
rect 17150 21330 17210 21400
rect 17280 21330 17300 21400
rect 17370 21330 17390 21400
rect 17460 21330 17480 21400
rect 17550 21330 17570 21400
rect 17640 21330 17660 21400
rect 17730 21330 17750 21400
rect 17820 21330 17840 21400
rect 17910 21330 17930 21400
rect 18000 21330 18020 21400
rect 18090 21330 18110 21400
rect 18180 21330 18200 21400
rect 18270 21330 18290 21400
rect 18360 21330 18380 21400
rect 18450 21330 18470 21400
rect 18540 21330 18560 21400
rect 18630 21330 18650 21400
rect 18720 21330 18740 21400
rect 18810 21330 18830 21400
rect 18900 21330 18920 21400
rect 18990 21330 19010 21400
rect 19080 21330 19100 21400
rect 19170 21330 19190 21400
rect 19260 21330 19280 21400
rect 19350 21330 19370 21400
rect 19440 21330 19460 21400
rect 19530 21330 19550 21400
rect 19620 21330 19640 21400
rect 19710 21330 19730 21400
rect 19800 21330 19820 21400
rect 19890 21330 19910 21400
rect 19980 21330 20000 21400
rect 20070 21330 20090 21400
rect 20160 21330 20450 21400
rect 8140 8690 20450 21330
rect 6440 8410 6760 8430
rect 6440 8340 6470 8410
rect 6540 8340 6560 8410
rect 6630 8340 6650 8410
rect 6720 8340 6760 8410
rect 6440 8320 6760 8340
rect 6440 8250 6470 8320
rect 6540 8250 6560 8320
rect 6630 8250 6650 8320
rect 6720 8250 6760 8320
rect 1540 6850 3140 6900
rect 1540 6780 1570 6850
rect 1640 6780 1680 6850
rect 1750 6780 1790 6850
rect 1860 6780 1900 6850
rect 1970 6780 2010 6850
rect 2080 6780 2120 6850
rect 2190 6780 2230 6850
rect 2300 6780 2340 6850
rect 2410 6780 2450 6850
rect 2520 6780 2560 6850
rect 2630 6780 2670 6850
rect 2740 6780 2780 6850
rect 2850 6780 2890 6850
rect 2960 6780 3000 6850
rect 3070 6780 3140 6850
rect 1540 6740 3140 6780
rect 1540 6670 1570 6740
rect 1640 6670 1680 6740
rect 1750 6670 1790 6740
rect 1860 6670 1900 6740
rect 1970 6670 2010 6740
rect 2080 6670 2120 6740
rect 2190 6670 2230 6740
rect 2300 6670 2340 6740
rect 2410 6670 2450 6740
rect 2520 6670 2560 6740
rect 2630 6670 2670 6740
rect 2740 6670 2780 6740
rect 2850 6670 2890 6740
rect 2960 6670 3000 6740
rect 3070 6670 3140 6740
rect 1540 6640 3140 6670
rect 6440 4610 6760 8250
rect 8140 8410 8460 8430
rect 8140 8340 8180 8410
rect 8250 8340 8270 8410
rect 8340 8340 8360 8410
rect 8430 8340 8460 8410
rect 8140 8320 8460 8340
rect 8140 8250 8180 8320
rect 8250 8250 8270 8320
rect 8340 8250 8360 8320
rect 8430 8250 8460 8320
rect 7400 5390 7490 5410
rect 7400 5320 7410 5390
rect 7480 5320 7490 5390
rect 7400 5280 7490 5320
rect 7400 5210 7410 5280
rect 7480 5210 7490 5280
rect 7400 5170 7490 5210
rect 7400 5100 7410 5170
rect 7480 5100 7490 5170
rect 7400 5060 7490 5100
rect 7400 4990 7410 5060
rect 7480 4990 7490 5060
rect 7400 4950 7490 4990
rect 7400 4880 7410 4950
rect 7480 4880 7490 4950
rect 7400 4860 7490 4880
rect 8140 4760 8460 8250
rect 31100 7820 38500 7910
rect 31100 7750 38190 7820
rect 38260 7750 38280 7820
rect 38350 7750 38370 7820
rect 38440 7750 38500 7820
rect 31100 7730 38500 7750
rect 31100 7660 38190 7730
rect 38260 7660 38280 7730
rect 38350 7660 38370 7730
rect 38440 7660 38500 7730
rect 31100 7640 38500 7660
rect 31100 7570 38190 7640
rect 38260 7570 38280 7640
rect 38350 7570 38370 7640
rect 38440 7570 38500 7640
rect 31100 7550 38500 7570
rect 31100 7480 38190 7550
rect 38260 7480 38280 7550
rect 38350 7480 38370 7550
rect 38440 7480 38500 7550
rect 31100 7460 38500 7480
rect 31100 7390 38190 7460
rect 38260 7390 38280 7460
rect 38350 7390 38370 7460
rect 38440 7390 38500 7460
rect 31100 7370 38500 7390
rect 31100 7300 38190 7370
rect 38260 7300 38280 7370
rect 38350 7300 38370 7370
rect 38440 7300 38500 7370
rect 31100 7280 38500 7300
rect 23460 7210 23940 7260
rect 23460 7140 23490 7210
rect 23560 7140 23600 7210
rect 23670 7140 23710 7210
rect 23780 7140 23820 7210
rect 23890 7140 23940 7210
rect 23460 7100 23940 7140
rect 23460 7030 23490 7100
rect 23560 7030 23600 7100
rect 23670 7030 23710 7100
rect 23780 7030 23820 7100
rect 23890 7030 23940 7100
rect 23460 7000 23940 7030
rect 25860 7210 26340 7260
rect 25860 7140 25890 7210
rect 25960 7140 26000 7210
rect 26070 7140 26110 7210
rect 26180 7140 26220 7210
rect 26290 7140 26340 7210
rect 25860 7100 26340 7140
rect 25860 7030 25890 7100
rect 25960 7030 26000 7100
rect 26070 7030 26110 7100
rect 26180 7030 26220 7100
rect 26290 7030 26340 7100
rect 25860 7000 26340 7030
rect 31100 7210 38190 7280
rect 38260 7210 38280 7280
rect 38350 7210 38370 7280
rect 38440 7210 38500 7280
rect 31100 7150 38500 7210
rect 31100 7080 38190 7150
rect 38260 7080 38280 7150
rect 38350 7080 38370 7150
rect 38440 7080 38500 7150
rect 31100 7060 38500 7080
rect 31100 6990 38190 7060
rect 38260 6990 38280 7060
rect 38350 6990 38370 7060
rect 38440 6990 38500 7060
rect 31100 6970 38500 6990
rect 11760 6880 13360 6930
rect 11760 6810 11790 6880
rect 11860 6810 11900 6880
rect 11970 6810 12010 6880
rect 12080 6810 12120 6880
rect 12190 6810 12230 6880
rect 12300 6810 12340 6880
rect 12410 6810 12450 6880
rect 12520 6810 12560 6880
rect 12630 6810 12670 6880
rect 12740 6810 12780 6880
rect 12850 6810 12890 6880
rect 12960 6810 13000 6880
rect 13070 6810 13110 6880
rect 13180 6810 13220 6880
rect 13290 6810 13360 6880
rect 11760 6770 13360 6810
rect 11760 6700 11790 6770
rect 11860 6700 11900 6770
rect 11970 6700 12010 6770
rect 12080 6700 12120 6770
rect 12190 6700 12230 6770
rect 12300 6700 12340 6770
rect 12410 6700 12450 6770
rect 12520 6700 12560 6770
rect 12630 6700 12670 6770
rect 12740 6700 12780 6770
rect 12850 6700 12890 6770
rect 12960 6700 13000 6770
rect 13070 6700 13110 6770
rect 13180 6700 13220 6770
rect 13290 6700 13360 6770
rect 11760 6670 13360 6700
rect 31100 6900 38190 6970
rect 38260 6900 38280 6970
rect 38350 6900 38370 6970
rect 38440 6900 38500 6970
rect 31100 6880 38500 6900
rect 31100 6810 38190 6880
rect 38260 6810 38280 6880
rect 38350 6810 38370 6880
rect 38440 6810 38500 6880
rect 31100 6790 38500 6810
rect 31100 6720 38190 6790
rect 38260 6720 38280 6790
rect 38350 6720 38370 6790
rect 38440 6720 38500 6790
rect 31100 6700 38500 6720
rect 31100 6630 38190 6700
rect 38260 6630 38280 6700
rect 38350 6630 38370 6700
rect 38440 6630 38500 6700
rect 31100 6610 38500 6630
rect 31100 6540 38190 6610
rect 38260 6540 38280 6610
rect 38350 6540 38370 6610
rect 38440 6540 38500 6610
rect 31100 6520 38500 6540
rect 31100 6450 38190 6520
rect 38260 6450 38280 6520
rect 38350 6450 38370 6520
rect 38440 6450 38500 6520
rect 31100 6430 38500 6450
rect 31100 6360 38190 6430
rect 38260 6360 38280 6430
rect 38350 6360 38370 6430
rect 38440 6360 38500 6430
rect 31100 6340 38500 6360
rect 30720 6300 30940 6320
rect 30720 6230 30740 6300
rect 30810 6230 30850 6300
rect 30920 6230 30940 6300
rect 30720 6170 30940 6230
rect 30720 6100 30740 6170
rect 30810 6100 30850 6170
rect 30920 6100 30940 6170
rect 30720 6040 30940 6100
rect 30720 5970 30740 6040
rect 30810 5970 30850 6040
rect 30920 5970 30940 6040
rect 30720 5950 30940 5970
rect 31100 6270 38190 6340
rect 38260 6270 38280 6340
rect 38350 6270 38370 6340
rect 38440 6270 38500 6340
rect 31100 6250 38500 6270
rect 31100 6180 38190 6250
rect 38260 6180 38280 6250
rect 38350 6180 38370 6250
rect 38440 6180 38500 6250
rect 31100 6160 38500 6180
rect 31100 6090 38190 6160
rect 38260 6090 38280 6160
rect 38350 6090 38370 6160
rect 38440 6090 38500 6160
rect 31100 6070 38500 6090
rect 31100 6000 38190 6070
rect 38260 6000 38280 6070
rect 38350 6000 38370 6070
rect 38440 6000 38500 6070
rect 31100 5980 38500 6000
rect 31100 5910 38190 5980
rect 38260 5910 38280 5980
rect 38350 5910 38370 5980
rect 38440 5910 38500 5980
rect 31100 5890 38500 5910
rect 31100 5820 38190 5890
rect 38260 5820 38280 5890
rect 38350 5820 38370 5890
rect 38440 5820 38500 5890
rect 31100 5800 38500 5820
rect 31100 5730 38190 5800
rect 38260 5730 38280 5800
rect 38350 5730 38370 5800
rect 38440 5730 38500 5800
rect 31100 5710 38500 5730
rect 8140 4700 8170 4760
rect 8230 4700 8270 4760
rect 8330 4700 8370 4760
rect 8430 4700 8460 4760
rect 8140 4670 8460 4700
rect 21800 5670 22020 5690
rect 21800 5600 21820 5670
rect 21890 5600 21930 5670
rect 22000 5600 22020 5670
rect 21800 5560 22020 5600
rect 21800 5490 21820 5560
rect 21890 5490 21930 5560
rect 22000 5490 22020 5560
rect 21800 5450 22020 5490
rect 21800 5380 21820 5450
rect 21890 5380 21930 5450
rect 22000 5380 22020 5450
rect 21800 5340 22020 5380
rect 21800 5270 21820 5340
rect 21890 5270 21930 5340
rect 22000 5270 22020 5340
rect 21800 5230 22020 5270
rect 21800 5160 21820 5230
rect 21890 5160 21930 5230
rect 22000 5160 22020 5230
rect 21800 5120 22020 5160
rect 21800 5050 21820 5120
rect 21890 5050 21930 5120
rect 22000 5050 22020 5120
rect 21800 5010 22020 5050
rect 21800 4940 21820 5010
rect 21890 4940 21930 5010
rect 22000 4940 22020 5010
rect 21800 4900 22020 4940
rect 21800 4830 21820 4900
rect 21890 4830 21930 4900
rect 22000 4830 22020 4900
rect 21800 4790 22020 4830
rect 21800 4720 21820 4790
rect 21890 4720 21930 4790
rect 22000 4720 22020 4790
rect 21800 4680 22020 4720
rect 21800 4610 21820 4680
rect 21890 4610 21930 4680
rect 22000 4610 22020 4680
rect -2520 4580 6210 4610
rect -2520 4510 -2490 4580
rect -2420 4520 6120 4580
rect 6180 4520 6210 4580
rect -2420 4510 6210 4520
rect -2520 4470 6210 4510
rect -2520 4400 -2490 4470
rect -2420 4460 6210 4470
rect -2420 4400 6120 4460
rect 6180 4400 6210 4460
rect -2520 4360 6210 4400
rect -2520 4290 -2490 4360
rect -2420 4340 6210 4360
rect -2420 4290 6120 4340
rect -2520 4280 6120 4290
rect 6180 4280 6210 4340
rect -2520 4250 6210 4280
rect -2520 4180 -2490 4250
rect -2420 4220 6210 4250
rect -2420 4180 6120 4220
rect -2520 4160 6120 4180
rect 6180 4160 6210 4220
rect -2520 4130 6210 4160
rect 6440 4580 17300 4610
rect 6440 4510 17200 4580
rect 17270 4510 17300 4580
rect 6440 4470 17300 4510
rect 21800 4570 22020 4610
rect 21800 4500 21820 4570
rect 21890 4500 21930 4570
rect 22000 4500 22020 4570
rect 21800 4480 22020 4500
rect 31100 5640 38190 5710
rect 38260 5640 38280 5710
rect 38350 5640 38370 5710
rect 38440 5640 38500 5710
rect 31100 5620 38500 5640
rect 31100 5550 38190 5620
rect 38260 5550 38280 5620
rect 38350 5550 38370 5620
rect 38440 5550 38500 5620
rect 31100 5530 38500 5550
rect 31100 5460 38190 5530
rect 38260 5460 38280 5530
rect 38350 5460 38370 5530
rect 38440 5460 38500 5530
rect 31100 5440 38500 5460
rect 31100 5370 38190 5440
rect 38260 5370 38280 5440
rect 38350 5370 38370 5440
rect 38440 5370 38500 5440
rect 31100 5350 38500 5370
rect 31100 5280 38190 5350
rect 38260 5280 38280 5350
rect 38350 5280 38370 5350
rect 38440 5280 38500 5350
rect 31100 5260 38500 5280
rect 31100 5190 38190 5260
rect 38260 5190 38280 5260
rect 38350 5190 38370 5260
rect 38440 5190 38500 5260
rect 31100 5170 38500 5190
rect 31100 5100 38190 5170
rect 38260 5100 38280 5170
rect 38350 5100 38370 5170
rect 38440 5100 38500 5170
rect 31100 5080 38500 5100
rect 31100 5010 38190 5080
rect 38260 5010 38280 5080
rect 38350 5010 38370 5080
rect 38440 5010 38500 5080
rect 31100 4990 38500 5010
rect 31100 4920 38190 4990
rect 38260 4920 38280 4990
rect 38350 4920 38370 4990
rect 38440 4920 38500 4990
rect 31100 4900 38500 4920
rect 31100 4830 38190 4900
rect 38260 4830 38280 4900
rect 38350 4830 38370 4900
rect 38440 4830 38500 4900
rect 31100 4810 38500 4830
rect 31100 4740 38190 4810
rect 38260 4740 38280 4810
rect 38350 4740 38370 4810
rect 38440 4740 38500 4810
rect 31100 4720 38500 4740
rect 31100 4650 38190 4720
rect 38260 4650 38280 4720
rect 38350 4650 38370 4720
rect 38440 4650 38500 4720
rect 31100 4630 38500 4650
rect 31100 4560 38190 4630
rect 38260 4560 38280 4630
rect 38350 4560 38370 4630
rect 38440 4560 38500 4630
rect 31100 4540 38500 4560
rect 6440 4400 17200 4470
rect 17270 4400 17300 4470
rect 6440 4360 17300 4400
rect 6440 4290 17200 4360
rect 17270 4290 17300 4360
rect 6440 4250 17300 4290
rect 6440 4180 17200 4250
rect 17270 4180 17300 4250
rect 6440 4130 17300 4180
rect 31100 4470 38190 4540
rect 38260 4470 38280 4540
rect 38350 4470 38370 4540
rect 38440 4470 38500 4540
rect 31100 4450 38500 4470
rect 31100 4380 38190 4450
rect 38260 4380 38280 4450
rect 38350 4380 38370 4450
rect 38440 4380 38500 4450
rect 31100 4360 38500 4380
rect 31100 4290 38190 4360
rect 38260 4290 38280 4360
rect 38350 4290 38370 4360
rect 38440 4290 38500 4360
rect 31100 4270 38500 4290
rect 31100 4200 38190 4270
rect 38260 4200 38280 4270
rect 38350 4200 38370 4270
rect 38440 4200 38500 4270
rect 31100 4140 38500 4200
rect 6440 3310 6760 4130
rect 31100 4070 38190 4140
rect 38260 4070 38280 4140
rect 38350 4070 38370 4140
rect 38440 4070 38500 4140
rect 31100 4050 38500 4070
rect 31100 3980 38190 4050
rect 38260 3980 38280 4050
rect 38350 3980 38370 4050
rect 38440 3980 38500 4050
rect 31100 3960 38500 3980
rect 31100 3890 38190 3960
rect 38260 3890 38280 3960
rect 38350 3890 38370 3960
rect 38440 3890 38500 3960
rect 31100 3870 38500 3890
rect 31100 3800 38190 3870
rect 38260 3800 38280 3870
rect 38350 3800 38370 3870
rect 38440 3800 38500 3870
rect 31100 3780 38500 3800
rect 31100 3710 38190 3780
rect 38260 3710 38280 3780
rect 38350 3710 38370 3780
rect 38440 3710 38500 3780
rect 31100 3690 38500 3710
rect 31100 3620 38190 3690
rect 38260 3620 38280 3690
rect 38350 3620 38370 3690
rect 38440 3620 38500 3690
rect 31100 3600 38500 3620
rect 31100 3530 38190 3600
rect 38260 3530 38280 3600
rect 38350 3530 38370 3600
rect 38440 3530 38500 3600
rect 31100 3510 38500 3530
rect 31100 3440 38190 3510
rect 38260 3440 38280 3510
rect 38350 3440 38370 3510
rect 38440 3440 38500 3510
rect 31100 3420 38500 3440
rect 24700 3360 25030 3380
rect 6440 3280 7340 3310
rect 6440 3220 7050 3280
rect 7110 3220 7150 3280
rect 7210 3220 7250 3280
rect 7310 3220 7340 3280
rect 6440 3180 7340 3220
rect 6440 3120 7050 3180
rect 7110 3120 7150 3180
rect 7210 3120 7250 3180
rect 7310 3120 7340 3180
rect 6440 3080 7340 3120
rect 6440 3020 7050 3080
rect 7110 3020 7150 3080
rect 7210 3020 7250 3080
rect 7310 3020 7340 3080
rect 24700 3290 24720 3360
rect 24790 3290 24830 3360
rect 24900 3290 24940 3360
rect 25010 3290 25030 3360
rect 24700 3250 25030 3290
rect 24700 3180 24720 3250
rect 24790 3180 24830 3250
rect 24900 3180 24940 3250
rect 25010 3180 25030 3250
rect 24700 3140 25030 3180
rect 24700 3070 24720 3140
rect 24790 3070 24830 3140
rect 24900 3070 24940 3140
rect 25010 3070 25030 3140
rect 24700 3050 25030 3070
rect 31100 3350 38190 3420
rect 38260 3350 38280 3420
rect 38350 3350 38370 3420
rect 38440 3350 38500 3420
rect 31100 3330 38500 3350
rect 31100 3260 38190 3330
rect 38260 3260 38280 3330
rect 38350 3260 38370 3330
rect 38440 3260 38500 3330
rect 31100 3240 38500 3260
rect 31100 3170 38190 3240
rect 38260 3170 38280 3240
rect 38350 3170 38370 3240
rect 38440 3170 38500 3240
rect 31100 3150 38500 3170
rect 31100 3080 38190 3150
rect 38260 3080 38280 3150
rect 38350 3080 38370 3150
rect 38440 3080 38500 3150
rect 31100 3060 38500 3080
rect 6440 3000 7340 3020
rect 31100 2990 38190 3060
rect 38260 2990 38280 3060
rect 38350 2990 38370 3060
rect 38440 2990 38500 3060
rect 31100 2970 38500 2990
rect 4740 2890 6750 2920
rect 4740 2830 4770 2890
rect 4830 2830 4870 2890
rect 4930 2830 4970 2890
rect 5030 2830 6750 2890
rect 4740 2790 6750 2830
rect 4740 2730 4770 2790
rect 4830 2730 4870 2790
rect 4930 2730 4970 2790
rect 5030 2730 6750 2790
rect 4740 2690 6750 2730
rect 4740 2630 4770 2690
rect 4830 2630 4870 2690
rect 4930 2630 4970 2690
rect 5030 2630 6750 2690
rect 4740 2610 6750 2630
rect -2920 1160 310 1180
rect -2920 1090 20 1160
rect 90 1090 130 1160
rect 200 1090 230 1160
rect 300 1090 310 1160
rect -2920 1050 310 1090
rect -2920 980 20 1050
rect 90 980 130 1050
rect 200 980 230 1050
rect 300 980 310 1050
rect -2920 940 310 980
rect -2920 870 20 940
rect 90 870 130 940
rect 200 870 230 940
rect 300 870 310 940
rect -2920 850 310 870
rect 6440 -100 6750 2610
rect -330 -140 6750 -100
rect -330 -210 -300 -140
rect -230 -210 -190 -140
rect -120 -210 -80 -140
rect -10 -210 30 -140
rect 100 -210 6750 -140
rect -330 -270 6750 -210
rect -330 -340 -300 -270
rect -230 -340 -190 -270
rect -120 -340 -80 -270
rect -10 -340 30 -270
rect 100 -340 6750 -270
rect -330 -380 6750 -340
rect 1080 -790 2680 -760
rect 1080 -860 1150 -790
rect 1220 -860 1260 -790
rect 1330 -860 1370 -790
rect 1440 -860 1480 -790
rect 1550 -860 1590 -790
rect 1660 -860 1700 -790
rect 1770 -860 1810 -790
rect 1880 -860 1920 -790
rect 1990 -860 2030 -790
rect 2100 -860 2140 -790
rect 2210 -860 2250 -790
rect 2320 -860 2360 -790
rect 2430 -860 2470 -790
rect 2540 -860 2580 -790
rect 2650 -860 2680 -790
rect 1080 -900 2680 -860
rect 1080 -970 1150 -900
rect 1220 -970 1260 -900
rect 1330 -970 1370 -900
rect 1440 -970 1480 -900
rect 1550 -970 1590 -900
rect 1660 -970 1700 -900
rect 1770 -970 1810 -900
rect 1880 -970 1920 -900
rect 1990 -970 2030 -900
rect 2100 -970 2140 -900
rect 2210 -970 2250 -900
rect 2320 -970 2360 -900
rect 2430 -970 2470 -900
rect 2540 -970 2580 -900
rect 2650 -970 2680 -900
rect 1080 -1020 2680 -970
rect 1540 -2780 3140 -2730
rect 1540 -2850 1570 -2780
rect 1640 -2850 1680 -2780
rect 1750 -2850 1790 -2780
rect 1860 -2850 1900 -2780
rect 1970 -2850 2010 -2780
rect 2080 -2850 2120 -2780
rect 2190 -2850 2230 -2780
rect 2300 -2850 2340 -2780
rect 2410 -2850 2450 -2780
rect 2520 -2850 2560 -2780
rect 2630 -2850 2670 -2780
rect 2740 -2850 2780 -2780
rect 2850 -2850 2890 -2780
rect 2960 -2850 3000 -2780
rect 3070 -2850 3140 -2780
rect 1540 -2890 3140 -2850
rect 1540 -2960 1570 -2890
rect 1640 -2960 1680 -2890
rect 1750 -2960 1790 -2890
rect 1860 -2960 1900 -2890
rect 1970 -2960 2010 -2890
rect 2080 -2960 2120 -2890
rect 2190 -2960 2230 -2890
rect 2300 -2960 2340 -2890
rect 2410 -2960 2450 -2890
rect 2520 -2960 2560 -2890
rect 2630 -2960 2670 -2890
rect 2740 -2960 2780 -2890
rect 2850 -2960 2890 -2890
rect 2960 -2960 3000 -2890
rect 3070 -2960 3140 -2890
rect 1540 -2990 3140 -2960
rect 6440 -4270 6750 -380
rect 8180 2890 10160 2920
rect 8180 2830 9870 2890
rect 9930 2830 9970 2890
rect 10030 2830 10070 2890
rect 10130 2830 10160 2890
rect 8180 2790 10160 2830
rect 8180 2730 9870 2790
rect 9930 2730 9970 2790
rect 10030 2730 10070 2790
rect 10130 2730 10160 2790
rect 8180 2690 10160 2730
rect 8180 2630 9870 2690
rect 9930 2630 9970 2690
rect 10030 2630 10070 2690
rect 10130 2630 10160 2690
rect 31100 2900 38190 2970
rect 38260 2900 38280 2970
rect 38350 2900 38370 2970
rect 38440 2900 38500 2970
rect 31100 2880 38500 2900
rect 31100 2810 38190 2880
rect 38260 2810 38280 2880
rect 38350 2810 38370 2880
rect 38440 2810 38500 2880
rect 31100 2790 38500 2810
rect 31100 2720 38190 2790
rect 38260 2720 38280 2790
rect 38350 2720 38370 2790
rect 38440 2720 38500 2790
rect 31100 2700 38500 2720
rect 31100 2630 38190 2700
rect 38260 2630 38280 2700
rect 38350 2630 38370 2700
rect 38440 2630 38500 2700
rect 8180 2610 10160 2630
rect 8180 -100 8490 2610
rect 22420 2600 22900 2630
rect 22420 2530 22470 2600
rect 22540 2530 22580 2600
rect 22650 2530 22690 2600
rect 22760 2530 22800 2600
rect 22870 2530 22900 2600
rect 22420 2490 22900 2530
rect 22420 2420 22470 2490
rect 22540 2420 22580 2490
rect 22650 2420 22690 2490
rect 22760 2420 22800 2490
rect 22870 2420 22900 2490
rect 22420 2370 22900 2420
rect 26900 2600 27380 2630
rect 26900 2530 26950 2600
rect 27020 2530 27060 2600
rect 27130 2530 27170 2600
rect 27240 2530 27280 2600
rect 27350 2530 27380 2600
rect 26900 2490 27380 2530
rect 26900 2420 26950 2490
rect 27020 2420 27060 2490
rect 27130 2420 27170 2490
rect 27240 2420 27280 2490
rect 27350 2420 27380 2490
rect 26900 2370 27380 2420
rect 31100 2610 38500 2630
rect 31100 2540 38190 2610
rect 38260 2540 38280 2610
rect 38350 2540 38370 2610
rect 38440 2540 38500 2610
rect 31100 2520 38500 2540
rect 31100 2450 38190 2520
rect 38260 2450 38280 2520
rect 38350 2450 38370 2520
rect 38440 2450 38500 2520
rect 31100 2430 38500 2450
rect 31100 2360 38190 2430
rect 38260 2360 38280 2430
rect 38350 2360 38370 2430
rect 38440 2360 38500 2430
rect 31100 2340 38500 2360
rect 31100 2270 38190 2340
rect 38260 2270 38280 2340
rect 38350 2270 38370 2340
rect 38440 2270 38500 2340
rect 31100 2250 38500 2270
rect 31100 2180 38190 2250
rect 38260 2180 38280 2250
rect 38350 2180 38370 2250
rect 38440 2180 38500 2250
rect 31100 2160 38500 2180
rect 31100 2090 38190 2160
rect 38260 2090 38280 2160
rect 38350 2090 38370 2160
rect 38440 2090 38500 2160
rect 31100 2070 38500 2090
rect 31100 2000 38190 2070
rect 38260 2000 38280 2070
rect 38350 2000 38370 2070
rect 38440 2000 38500 2070
rect 31100 1980 38500 2000
rect 31100 1910 38190 1980
rect 38260 1910 38280 1980
rect 38350 1910 38370 1980
rect 38440 1910 38500 1980
rect 31100 1890 38500 1910
rect 31100 1820 38190 1890
rect 38260 1820 38280 1890
rect 38350 1820 38370 1890
rect 38440 1820 38500 1890
rect 31100 1800 38500 1820
rect 31100 1730 38190 1800
rect 38260 1730 38280 1800
rect 38350 1730 38370 1800
rect 38440 1730 38500 1800
rect 31100 1710 38500 1730
rect 31100 1640 38190 1710
rect 38260 1640 38280 1710
rect 38350 1640 38370 1710
rect 38440 1640 38500 1710
rect 31100 1620 38500 1640
rect 31100 1550 38190 1620
rect 38260 1550 38280 1620
rect 38350 1550 38370 1620
rect 38440 1550 38500 1620
rect 31100 1530 38500 1550
rect 31100 1460 38190 1530
rect 38260 1460 38280 1530
rect 38350 1460 38370 1530
rect 38440 1460 38500 1530
rect 31100 1440 38500 1460
rect 31100 1370 38190 1440
rect 38260 1370 38280 1440
rect 38350 1370 38370 1440
rect 38440 1370 38500 1440
rect 31100 1350 38500 1370
rect 31100 1280 38190 1350
rect 38260 1280 38280 1350
rect 38350 1280 38370 1350
rect 38440 1280 38500 1350
rect 31100 1260 38500 1280
rect 31100 1190 38190 1260
rect 38260 1190 38280 1260
rect 38350 1190 38370 1260
rect 38440 1190 38500 1260
rect 14590 1160 19085 1180
rect 14590 1090 14600 1160
rect 14670 1090 14700 1160
rect 14770 1090 14810 1160
rect 14880 1090 18995 1160
rect 19065 1090 19085 1160
rect 31100 1150 38500 1190
rect 14590 1050 19085 1090
rect 14590 980 14600 1050
rect 14670 980 14700 1050
rect 14770 980 14810 1050
rect 14880 980 18995 1050
rect 19065 980 19085 1050
rect 14590 940 19085 980
rect 14590 870 14600 940
rect 14670 870 14700 940
rect 14770 870 14810 940
rect 14880 870 18995 940
rect 19065 870 19085 940
rect 14590 850 19085 870
rect 23460 920 23940 970
rect 23460 850 23490 920
rect 23560 850 23600 920
rect 23670 850 23710 920
rect 23780 850 23820 920
rect 23890 850 23940 920
rect 23460 810 23940 850
rect 23460 740 23490 810
rect 23560 740 23600 810
rect 23670 740 23710 810
rect 23780 740 23820 810
rect 23890 740 23940 810
rect 23460 710 23940 740
rect 25860 920 26340 970
rect 25860 850 25890 920
rect 25960 850 26000 920
rect 26070 850 26110 920
rect 26180 850 26220 920
rect 26290 850 26340 920
rect 25860 810 26340 850
rect 25860 740 25890 810
rect 25960 740 26000 810
rect 26070 740 26110 810
rect 26180 740 26220 810
rect 26290 740 26340 810
rect 25860 710 26340 740
rect 31100 220 38500 310
rect 31100 150 38190 220
rect 38260 150 38280 220
rect 38350 150 38370 220
rect 38440 150 38500 220
rect 31100 130 38500 150
rect 31100 60 38190 130
rect 38260 60 38280 130
rect 38350 60 38370 130
rect 38440 60 38500 130
rect 31100 40 38500 60
rect 30720 0 30940 20
rect 30720 -70 30740 0
rect 30810 -70 30850 0
rect 30920 -70 30940 0
rect 8180 -140 15110 -100
rect 8180 -210 14660 -140
rect 14730 -210 14770 -140
rect 14840 -210 14880 -140
rect 14950 -210 14990 -140
rect 15060 -210 15110 -140
rect 8180 -270 15110 -210
rect 8180 -340 14660 -270
rect 14730 -340 14770 -270
rect 14840 -340 14880 -270
rect 14950 -340 14990 -270
rect 15060 -340 15110 -270
rect 8180 -380 15110 -340
rect 30720 -130 30940 -70
rect 30720 -200 30740 -130
rect 30810 -200 30850 -130
rect 30920 -200 30940 -130
rect 30720 -260 30940 -200
rect 30720 -330 30740 -260
rect 30810 -330 30850 -260
rect 30920 -330 30940 -260
rect 30720 -350 30940 -330
rect 31100 -30 38190 40
rect 38260 -30 38280 40
rect 38350 -30 38370 40
rect 38440 -30 38500 40
rect 31100 -50 38500 -30
rect 31100 -120 38190 -50
rect 38260 -120 38280 -50
rect 38350 -120 38370 -50
rect 38440 -120 38500 -50
rect 31100 -140 38500 -120
rect 31100 -210 38190 -140
rect 38260 -210 38280 -140
rect 38350 -210 38370 -140
rect 38440 -210 38500 -140
rect 31100 -230 38500 -210
rect 31100 -300 38190 -230
rect 38260 -300 38280 -230
rect 38350 -300 38370 -230
rect 38440 -300 38500 -230
rect 31100 -320 38500 -300
rect 7290 -3880 7620 -3860
rect 7290 -3950 7310 -3880
rect 7380 -3950 7420 -3880
rect 7490 -3950 7530 -3880
rect 7600 -3950 7620 -3880
rect 7290 -3990 7620 -3950
rect 7290 -4060 7310 -3990
rect 7380 -4060 7420 -3990
rect 7490 -4060 7530 -3990
rect 7600 -4060 7620 -3990
rect 7290 -4100 7620 -4060
rect 7290 -4170 7310 -4100
rect 7380 -4170 7420 -4100
rect 7490 -4170 7530 -4100
rect 7600 -4170 7620 -4100
rect 7290 -4190 7620 -4170
rect -590 -4290 6750 -4270
rect -1350 -4350 -910 -4330
rect -1350 -4420 -1330 -4350
rect -1260 -4420 -1220 -4350
rect -1150 -4420 -1110 -4350
rect -1040 -4420 -1000 -4350
rect -930 -4420 -910 -4350
rect -1350 -4460 -910 -4420
rect -1350 -4530 -1330 -4460
rect -1260 -4530 -1220 -4460
rect -1150 -4530 -1110 -4460
rect -1040 -4530 -1000 -4460
rect -930 -4530 -910 -4460
rect -1350 -4550 -910 -4530
rect -590 -4360 -560 -4290
rect -490 -4360 -450 -4290
rect -380 -4360 -340 -4290
rect -270 -4360 -230 -4290
rect -160 -4360 6750 -4290
rect -590 -4400 6750 -4360
rect -590 -4470 -560 -4400
rect -490 -4470 -450 -4400
rect -380 -4470 -340 -4400
rect -270 -4470 -230 -4400
rect -160 -4470 6750 -4400
rect -590 -4550 6750 -4470
rect -1350 -6330 260 -4630
rect -1350 -6400 -1160 -6330
rect -1090 -6400 -1070 -6330
rect -1000 -6400 -980 -6330
rect -910 -6400 -890 -6330
rect -820 -6400 -800 -6330
rect -730 -6400 -710 -6330
rect -640 -6400 -620 -6330
rect -550 -6400 -530 -6330
rect -460 -6400 -440 -6330
rect -370 -6400 -350 -6330
rect -280 -6400 -260 -6330
rect -190 -6400 -170 -6330
rect -100 -6400 -80 -6330
rect -10 -6400 10 -6330
rect 80 -6400 260 -6330
rect -1350 -6420 260 -6400
rect -1740 -6520 -1600 -6470
rect -1740 -6590 -1710 -6520
rect -1640 -6590 -1600 -6520
rect -1740 -6630 -1600 -6590
rect -1740 -6700 -1710 -6630
rect -1640 -6640 -1600 -6630
rect -1350 -6490 -1160 -6420
rect -1090 -6490 -1070 -6420
rect -1000 -6490 -980 -6420
rect -910 -6490 -890 -6420
rect -820 -6490 -800 -6420
rect -730 -6490 -710 -6420
rect -640 -6490 -620 -6420
rect -550 -6490 -530 -6420
rect -460 -6490 -440 -6420
rect -370 -6490 -350 -6420
rect -280 -6490 -260 -6420
rect -190 -6490 -170 -6420
rect -100 -6490 -80 -6420
rect -10 -6490 10 -6420
rect 80 -6490 260 -6420
rect -1350 -6510 260 -6490
rect -1350 -6580 -1160 -6510
rect -1090 -6580 -1070 -6510
rect -1000 -6580 -980 -6510
rect -910 -6580 -890 -6510
rect -820 -6580 -800 -6510
rect -730 -6580 -710 -6510
rect -640 -6580 -620 -6510
rect -550 -6580 -530 -6510
rect -460 -6580 -440 -6510
rect -370 -6580 -350 -6510
rect -280 -6580 -260 -6510
rect -190 -6580 -170 -6510
rect -100 -6580 -80 -6510
rect -10 -6580 10 -6510
rect 80 -6580 260 -6510
rect -1350 -6640 260 -6580
rect 6440 -6420 6750 -4550
rect 8180 -4270 8490 -380
rect 31100 -390 38190 -320
rect 38260 -390 38280 -320
rect 38350 -390 38370 -320
rect 38440 -390 38500 -320
rect 31100 -450 38500 -390
rect 31100 -520 38190 -450
rect 38260 -520 38280 -450
rect 38350 -520 38370 -450
rect 38440 -520 38500 -450
rect 31100 -540 38500 -520
rect 31100 -610 38190 -540
rect 38260 -610 38280 -540
rect 38350 -610 38370 -540
rect 38440 -610 38500 -540
rect 31100 -630 38500 -610
rect 31100 -700 38190 -630
rect 38260 -700 38280 -630
rect 38350 -700 38370 -630
rect 38440 -700 38500 -630
rect 31100 -720 38500 -700
rect 12220 -790 13820 -760
rect 12220 -860 12250 -790
rect 12320 -860 12360 -790
rect 12430 -860 12470 -790
rect 12540 -860 12580 -790
rect 12650 -860 12690 -790
rect 12760 -860 12800 -790
rect 12870 -860 12910 -790
rect 12980 -860 13020 -790
rect 13090 -860 13130 -790
rect 13200 -860 13240 -790
rect 13310 -860 13350 -790
rect 13420 -860 13460 -790
rect 13530 -860 13570 -790
rect 13640 -860 13680 -790
rect 13750 -860 13820 -790
rect 31100 -790 38190 -720
rect 38260 -790 38280 -720
rect 38350 -790 38370 -720
rect 38440 -790 38500 -720
rect 31100 -810 38500 -790
rect 12220 -900 13820 -860
rect 12220 -970 12250 -900
rect 12320 -970 12360 -900
rect 12430 -970 12470 -900
rect 12540 -970 12580 -900
rect 12650 -970 12690 -900
rect 12760 -970 12800 -900
rect 12870 -970 12910 -900
rect 12980 -970 13020 -900
rect 13090 -970 13130 -900
rect 13200 -970 13240 -900
rect 13310 -970 13350 -900
rect 13420 -970 13460 -900
rect 13530 -970 13570 -900
rect 13640 -970 13680 -900
rect 13750 -970 13820 -900
rect 12220 -1020 13820 -970
rect 21800 -850 22020 -830
rect 21800 -920 21820 -850
rect 21890 -920 21930 -850
rect 22000 -920 22020 -850
rect 21800 -960 22020 -920
rect 21800 -1030 21820 -960
rect 21890 -1030 21930 -960
rect 22000 -1030 22020 -960
rect 21800 -1070 22020 -1030
rect 21800 -1140 21820 -1070
rect 21890 -1140 21930 -1070
rect 22000 -1140 22020 -1070
rect 21800 -1180 22020 -1140
rect 21800 -1250 21820 -1180
rect 21890 -1250 21930 -1180
rect 22000 -1250 22020 -1180
rect 21800 -1290 22020 -1250
rect 21800 -1360 21820 -1290
rect 21890 -1360 21930 -1290
rect 22000 -1360 22020 -1290
rect 21800 -1400 22020 -1360
rect 21800 -1470 21820 -1400
rect 21890 -1470 21930 -1400
rect 22000 -1470 22020 -1400
rect 21800 -1510 22020 -1470
rect 21800 -1580 21820 -1510
rect 21890 -1580 21930 -1510
rect 22000 -1580 22020 -1510
rect 21800 -1620 22020 -1580
rect 21800 -1690 21820 -1620
rect 21890 -1690 21930 -1620
rect 22000 -1690 22020 -1620
rect 21800 -1730 22020 -1690
rect 21800 -1800 21820 -1730
rect 21890 -1800 21930 -1730
rect 22000 -1800 22020 -1730
rect 21800 -1840 22020 -1800
rect 21800 -1910 21820 -1840
rect 21890 -1910 21930 -1840
rect 22000 -1910 22020 -1840
rect 21800 -1950 22020 -1910
rect 21800 -2020 21820 -1950
rect 21890 -2020 21930 -1950
rect 22000 -2020 22020 -1950
rect 21800 -2040 22020 -2020
rect 31100 -880 38190 -810
rect 38260 -880 38280 -810
rect 38350 -880 38370 -810
rect 38440 -880 38500 -810
rect 31100 -900 38500 -880
rect 31100 -970 38190 -900
rect 38260 -970 38280 -900
rect 38350 -970 38370 -900
rect 38440 -970 38500 -900
rect 31100 -990 38500 -970
rect 31100 -1060 38190 -990
rect 38260 -1060 38280 -990
rect 38350 -1060 38370 -990
rect 38440 -1060 38500 -990
rect 31100 -1080 38500 -1060
rect 31100 -1150 38190 -1080
rect 38260 -1150 38280 -1080
rect 38350 -1150 38370 -1080
rect 38440 -1150 38500 -1080
rect 31100 -1170 38500 -1150
rect 31100 -1240 38190 -1170
rect 38260 -1240 38280 -1170
rect 38350 -1240 38370 -1170
rect 38440 -1240 38500 -1170
rect 31100 -1260 38500 -1240
rect 31100 -1330 38190 -1260
rect 38260 -1330 38280 -1260
rect 38350 -1330 38370 -1260
rect 38440 -1330 38500 -1260
rect 31100 -1350 38500 -1330
rect 31100 -1420 38190 -1350
rect 38260 -1420 38280 -1350
rect 38350 -1420 38370 -1350
rect 38440 -1420 38500 -1350
rect 31100 -1440 38500 -1420
rect 31100 -1510 38190 -1440
rect 38260 -1510 38280 -1440
rect 38350 -1510 38370 -1440
rect 38440 -1510 38500 -1440
rect 31100 -1530 38500 -1510
rect 31100 -1600 38190 -1530
rect 38260 -1600 38280 -1530
rect 38350 -1600 38370 -1530
rect 38440 -1600 38500 -1530
rect 31100 -1620 38500 -1600
rect 31100 -1690 38190 -1620
rect 38260 -1690 38280 -1620
rect 38350 -1690 38370 -1620
rect 38440 -1690 38500 -1620
rect 31100 -1710 38500 -1690
rect 31100 -1780 38190 -1710
rect 38260 -1780 38280 -1710
rect 38350 -1780 38370 -1710
rect 38440 -1780 38500 -1710
rect 31100 -1800 38500 -1780
rect 31100 -1870 38190 -1800
rect 38260 -1870 38280 -1800
rect 38350 -1870 38370 -1800
rect 38440 -1870 38500 -1800
rect 31100 -1890 38500 -1870
rect 31100 -1960 38190 -1890
rect 38260 -1960 38280 -1890
rect 38350 -1960 38370 -1890
rect 38440 -1960 38500 -1890
rect 31100 -1980 38500 -1960
rect 31100 -2050 38190 -1980
rect 38260 -2050 38280 -1980
rect 38350 -2050 38370 -1980
rect 38440 -2050 38500 -1980
rect 31100 -2070 38500 -2050
rect 31100 -2140 38190 -2070
rect 38260 -2140 38280 -2070
rect 38350 -2140 38370 -2070
rect 38440 -2140 38500 -2070
rect 31100 -2160 38500 -2140
rect 31100 -2230 38190 -2160
rect 38260 -2230 38280 -2160
rect 38350 -2230 38370 -2160
rect 38440 -2230 38500 -2160
rect 31100 -2250 38500 -2230
rect 31100 -2320 38190 -2250
rect 38260 -2320 38280 -2250
rect 38350 -2320 38370 -2250
rect 38440 -2320 38500 -2250
rect 31100 -2340 38500 -2320
rect 31100 -2410 38190 -2340
rect 38260 -2410 38280 -2340
rect 38350 -2410 38370 -2340
rect 38440 -2410 38500 -2340
rect 31100 -2430 38500 -2410
rect 31100 -2500 38190 -2430
rect 38260 -2500 38280 -2430
rect 38350 -2500 38370 -2430
rect 38440 -2500 38500 -2430
rect 31100 -2520 38500 -2500
rect 31100 -2590 38190 -2520
rect 38260 -2590 38280 -2520
rect 38350 -2590 38370 -2520
rect 38440 -2590 38500 -2520
rect 31100 -2610 38500 -2590
rect 31100 -2680 38190 -2610
rect 38260 -2680 38280 -2610
rect 38350 -2680 38370 -2610
rect 38440 -2680 38500 -2610
rect 31100 -2700 38500 -2680
rect 11760 -2780 13360 -2730
rect 11760 -2850 11790 -2780
rect 11860 -2850 11900 -2780
rect 11970 -2850 12010 -2780
rect 12080 -2850 12120 -2780
rect 12190 -2850 12230 -2780
rect 12300 -2850 12340 -2780
rect 12410 -2850 12450 -2780
rect 12520 -2850 12560 -2780
rect 12630 -2850 12670 -2780
rect 12740 -2850 12780 -2780
rect 12850 -2850 12890 -2780
rect 12960 -2850 13000 -2780
rect 13070 -2850 13110 -2780
rect 13180 -2850 13220 -2780
rect 13290 -2850 13360 -2780
rect 11760 -2890 13360 -2850
rect 11760 -2960 11790 -2890
rect 11860 -2960 11900 -2890
rect 11970 -2960 12010 -2890
rect 12080 -2960 12120 -2890
rect 12190 -2960 12230 -2890
rect 12300 -2960 12340 -2890
rect 12410 -2960 12450 -2890
rect 12520 -2960 12560 -2890
rect 12630 -2960 12670 -2890
rect 12740 -2960 12780 -2890
rect 12850 -2960 12890 -2890
rect 12960 -2960 13000 -2890
rect 13070 -2960 13110 -2890
rect 13180 -2960 13220 -2890
rect 13290 -2960 13360 -2890
rect 11760 -2990 13360 -2960
rect 31100 -2770 38190 -2700
rect 38260 -2770 38280 -2700
rect 38350 -2770 38370 -2700
rect 38440 -2770 38500 -2700
rect 31100 -2790 38500 -2770
rect 31100 -2860 38190 -2790
rect 38260 -2860 38280 -2790
rect 38350 -2860 38370 -2790
rect 38440 -2860 38500 -2790
rect 31100 -2880 38500 -2860
rect 31100 -2950 38190 -2880
rect 38260 -2950 38280 -2880
rect 38350 -2950 38370 -2880
rect 38440 -2950 38500 -2880
rect 31100 -2970 38500 -2950
rect 24720 -3050 25050 -3030
rect 24720 -3120 24740 -3050
rect 24810 -3120 24850 -3050
rect 24920 -3120 24960 -3050
rect 25030 -3120 25050 -3050
rect 24720 -3160 25050 -3120
rect 24720 -3230 24740 -3160
rect 24810 -3230 24850 -3160
rect 24920 -3230 24960 -3160
rect 25030 -3230 25050 -3160
rect 24720 -3270 25050 -3230
rect 24720 -3340 24740 -3270
rect 24810 -3340 24850 -3270
rect 24920 -3340 24960 -3270
rect 25030 -3340 25050 -3270
rect 24720 -3360 25050 -3340
rect 31100 -3040 38190 -2970
rect 38260 -3040 38280 -2970
rect 38350 -3040 38370 -2970
rect 38440 -3040 38500 -2970
rect 31100 -3060 38500 -3040
rect 31100 -3130 38190 -3060
rect 38260 -3130 38280 -3060
rect 38350 -3130 38370 -3060
rect 38440 -3130 38500 -3060
rect 31100 -3150 38500 -3130
rect 31100 -3220 38190 -3150
rect 38260 -3220 38280 -3150
rect 38350 -3220 38370 -3150
rect 38440 -3220 38500 -3150
rect 31100 -3240 38500 -3220
rect 31100 -3310 38190 -3240
rect 38260 -3310 38280 -3240
rect 38350 -3310 38370 -3240
rect 38440 -3310 38500 -3240
rect 31100 -3330 38500 -3310
rect 31100 -3400 38190 -3330
rect 38260 -3400 38280 -3330
rect 38350 -3400 38370 -3330
rect 38440 -3400 38500 -3330
rect 31100 -3460 38500 -3400
rect 31100 -3530 38190 -3460
rect 38260 -3530 38280 -3460
rect 38350 -3530 38370 -3460
rect 38440 -3530 38500 -3460
rect 31100 -3550 38500 -3530
rect 31100 -3620 38190 -3550
rect 38260 -3620 38280 -3550
rect 38350 -3620 38370 -3550
rect 38440 -3620 38500 -3550
rect 31100 -3640 38500 -3620
rect 22420 -3690 22900 -3660
rect 22420 -3760 22470 -3690
rect 22540 -3760 22580 -3690
rect 22650 -3760 22690 -3690
rect 22760 -3760 22800 -3690
rect 22870 -3760 22900 -3690
rect 22420 -3800 22900 -3760
rect 22420 -3870 22470 -3800
rect 22540 -3870 22580 -3800
rect 22650 -3870 22690 -3800
rect 22760 -3870 22800 -3800
rect 22870 -3870 22900 -3800
rect 22420 -3920 22900 -3870
rect 26900 -3690 27380 -3660
rect 26900 -3760 26950 -3690
rect 27020 -3760 27060 -3690
rect 27130 -3760 27170 -3690
rect 27240 -3760 27280 -3690
rect 27350 -3760 27380 -3690
rect 26900 -3800 27380 -3760
rect 26900 -3870 26950 -3800
rect 27020 -3870 27060 -3800
rect 27130 -3870 27170 -3800
rect 27240 -3870 27280 -3800
rect 27350 -3870 27380 -3800
rect 26900 -3920 27380 -3870
rect 31100 -3710 38190 -3640
rect 38260 -3710 38280 -3640
rect 38350 -3710 38370 -3640
rect 38440 -3710 38500 -3640
rect 31100 -3730 38500 -3710
rect 31100 -3800 38190 -3730
rect 38260 -3800 38280 -3730
rect 38350 -3800 38370 -3730
rect 38440 -3800 38500 -3730
rect 31100 -3820 38500 -3800
rect 31100 -3890 38190 -3820
rect 38260 -3890 38280 -3820
rect 38350 -3890 38370 -3820
rect 38440 -3890 38500 -3820
rect 31100 -3910 38500 -3890
rect 31100 -3980 38190 -3910
rect 38260 -3980 38280 -3910
rect 38350 -3980 38370 -3910
rect 38440 -3980 38500 -3910
rect 31100 -4000 38500 -3980
rect 31100 -4070 38190 -4000
rect 38260 -4070 38280 -4000
rect 38350 -4070 38370 -4000
rect 38440 -4070 38500 -4000
rect 31100 -4090 38500 -4070
rect 31100 -4160 38190 -4090
rect 38260 -4160 38280 -4090
rect 38350 -4160 38370 -4090
rect 38440 -4160 38500 -4090
rect 31100 -4180 38500 -4160
rect 31100 -4250 38190 -4180
rect 38260 -4250 38280 -4180
rect 38350 -4250 38370 -4180
rect 38440 -4250 38500 -4180
rect 31100 -4270 38500 -4250
rect 8180 -4290 15370 -4270
rect 8180 -4360 14940 -4290
rect 15010 -4360 15050 -4290
rect 15120 -4360 15160 -4290
rect 15230 -4360 15270 -4290
rect 15340 -4360 15370 -4290
rect 8180 -4400 15370 -4360
rect 8180 -4470 14940 -4400
rect 15010 -4470 15050 -4400
rect 15120 -4470 15160 -4400
rect 15230 -4470 15270 -4400
rect 15340 -4470 15370 -4400
rect 8180 -4550 15370 -4470
rect 15690 -4350 16130 -4330
rect 15690 -4420 15710 -4350
rect 15780 -4420 15820 -4350
rect 15890 -4420 15930 -4350
rect 16000 -4420 16040 -4350
rect 16110 -4420 16130 -4350
rect 15690 -4460 16130 -4420
rect 15690 -4530 15710 -4460
rect 15780 -4530 15820 -4460
rect 15890 -4530 15930 -4460
rect 16000 -4530 16040 -4460
rect 16110 -4530 16130 -4460
rect 15690 -4550 16130 -4530
rect 31100 -4340 38190 -4270
rect 38260 -4340 38280 -4270
rect 38350 -4340 38370 -4270
rect 38440 -4340 38500 -4270
rect 31100 -4360 38500 -4340
rect 31100 -4430 38190 -4360
rect 38260 -4430 38280 -4360
rect 38350 -4430 38370 -4360
rect 38440 -4430 38500 -4360
rect 31100 -4450 38500 -4430
rect 31100 -4520 38190 -4450
rect 38260 -4520 38280 -4450
rect 38350 -4520 38370 -4450
rect 38440 -4520 38500 -4450
rect 31100 -4540 38500 -4520
rect 8180 -6420 8490 -4550
rect 31100 -4610 38190 -4540
rect 38260 -4610 38280 -4540
rect 38350 -4610 38370 -4540
rect 38440 -4610 38500 -4540
rect 31100 -4630 38500 -4610
rect 6440 -6460 7340 -6420
rect 6440 -6520 7050 -6460
rect 7110 -6520 7150 -6460
rect 7210 -6520 7250 -6460
rect 7310 -6520 7340 -6460
rect 6440 -6560 7340 -6520
rect 6440 -6620 7050 -6560
rect 7110 -6620 7150 -6560
rect 7210 -6620 7250 -6560
rect 7310 -6620 7340 -6560
rect -1640 -6670 6190 -6640
rect -1640 -6700 4770 -6670
rect -1740 -6730 4770 -6700
rect 4830 -6730 4870 -6670
rect 4930 -6730 4970 -6670
rect 5030 -6730 6190 -6670
rect -1740 -6740 6190 -6730
rect -1740 -6810 -1710 -6740
rect -1640 -6770 6190 -6740
rect -1640 -6810 4770 -6770
rect -1740 -6830 4770 -6810
rect 4830 -6830 4870 -6770
rect 4930 -6830 4970 -6770
rect 5030 -6830 6190 -6770
rect -1740 -6850 6190 -6830
rect 6440 -6660 7340 -6620
rect 6440 -6720 7050 -6660
rect 7110 -6720 7150 -6660
rect 7210 -6720 7250 -6660
rect 7310 -6720 7340 -6660
rect 6440 -6760 7340 -6720
rect 6440 -6820 7050 -6760
rect 7110 -6820 7150 -6760
rect 7210 -6820 7250 -6760
rect 7310 -6820 7340 -6760
rect 6440 -6850 7340 -6820
rect 7560 -6460 8490 -6420
rect 7560 -6520 7590 -6460
rect 7650 -6520 7690 -6460
rect 7750 -6520 7790 -6460
rect 7850 -6520 8490 -6460
rect 7560 -6560 8490 -6520
rect 7560 -6620 7590 -6560
rect 7650 -6620 7690 -6560
rect 7750 -6620 7790 -6560
rect 7850 -6620 8490 -6560
rect 7560 -6660 8490 -6620
rect 14520 -6330 16130 -4630
rect 14520 -6400 14700 -6330
rect 14770 -6400 14790 -6330
rect 14860 -6400 14880 -6330
rect 14950 -6400 14970 -6330
rect 15040 -6400 15060 -6330
rect 15130 -6400 15150 -6330
rect 15220 -6400 15240 -6330
rect 15310 -6400 15330 -6330
rect 15400 -6400 15420 -6330
rect 15490 -6400 15510 -6330
rect 15580 -6400 15600 -6330
rect 15670 -6400 15690 -6330
rect 15760 -6400 15780 -6330
rect 15850 -6400 15870 -6330
rect 15940 -6400 16130 -6330
rect 14520 -6420 16130 -6400
rect 14520 -6490 14700 -6420
rect 14770 -6490 14790 -6420
rect 14860 -6490 14880 -6420
rect 14950 -6490 14970 -6420
rect 15040 -6490 15060 -6420
rect 15130 -6490 15150 -6420
rect 15220 -6490 15240 -6420
rect 15310 -6490 15330 -6420
rect 15400 -6490 15420 -6420
rect 15490 -6490 15510 -6420
rect 15580 -6490 15600 -6420
rect 15670 -6490 15690 -6420
rect 15760 -6490 15780 -6420
rect 15850 -6490 15870 -6420
rect 15940 -6490 16130 -6420
rect 31100 -4700 38190 -4630
rect 38260 -4700 38280 -4630
rect 38350 -4700 38370 -4630
rect 38440 -4700 38500 -4630
rect 31100 -4720 38500 -4700
rect 31100 -4790 38190 -4720
rect 38260 -4790 38280 -4720
rect 38350 -4790 38370 -4720
rect 38440 -4790 38500 -4720
rect 31100 -4810 38500 -4790
rect 31100 -4880 38190 -4810
rect 38260 -4880 38280 -4810
rect 38350 -4880 38370 -4810
rect 38440 -4880 38500 -4810
rect 31100 -4900 38500 -4880
rect 31100 -4970 38190 -4900
rect 38260 -4970 38280 -4900
rect 38350 -4970 38370 -4900
rect 38440 -4970 38500 -4900
rect 31100 -4990 38500 -4970
rect 31100 -5060 38190 -4990
rect 38260 -5060 38280 -4990
rect 38350 -5060 38370 -4990
rect 38440 -5060 38500 -4990
rect 31100 -5080 38500 -5060
rect 31100 -5150 38190 -5080
rect 38260 -5150 38280 -5080
rect 38350 -5150 38370 -5080
rect 38440 -5150 38500 -5080
rect 31100 -5170 38500 -5150
rect 31100 -5240 38190 -5170
rect 38260 -5240 38280 -5170
rect 38350 -5240 38370 -5170
rect 38440 -5240 38500 -5170
rect 31100 -5260 38500 -5240
rect 31100 -5330 38190 -5260
rect 38260 -5330 38280 -5260
rect 38350 -5330 38370 -5260
rect 38440 -5330 38500 -5260
rect 31100 -5350 38500 -5330
rect 31100 -5420 38190 -5350
rect 38260 -5420 38280 -5350
rect 38350 -5420 38370 -5350
rect 38440 -5420 38500 -5350
rect 31100 -5440 38500 -5420
rect 31100 -5510 38190 -5440
rect 38260 -5510 38280 -5440
rect 38350 -5510 38370 -5440
rect 38440 -5510 38500 -5440
rect 31100 -5530 38500 -5510
rect 31100 -5600 38190 -5530
rect 38260 -5600 38280 -5530
rect 38350 -5600 38370 -5530
rect 38440 -5600 38500 -5530
rect 31100 -5620 38500 -5600
rect 31100 -5690 38190 -5620
rect 38260 -5690 38280 -5620
rect 38350 -5690 38370 -5620
rect 38440 -5690 38500 -5620
rect 31100 -5710 38500 -5690
rect 31100 -5780 38190 -5710
rect 38260 -5780 38280 -5710
rect 38350 -5780 38370 -5710
rect 38440 -5780 38500 -5710
rect 31100 -5800 38500 -5780
rect 31100 -5870 38190 -5800
rect 38260 -5870 38280 -5800
rect 38350 -5870 38370 -5800
rect 38440 -5870 38500 -5800
rect 31100 -5890 38500 -5870
rect 31100 -5960 38190 -5890
rect 38260 -5960 38280 -5890
rect 38350 -5960 38370 -5890
rect 38440 -5960 38500 -5890
rect 31100 -5980 38500 -5960
rect 31100 -6050 38190 -5980
rect 38260 -6050 38280 -5980
rect 38350 -6050 38370 -5980
rect 38440 -6050 38500 -5980
rect 31100 -6070 38500 -6050
rect 31100 -6140 38190 -6070
rect 38260 -6140 38280 -6070
rect 38350 -6140 38370 -6070
rect 38440 -6140 38500 -6070
rect 31100 -6160 38500 -6140
rect 31100 -6230 38190 -6160
rect 38260 -6230 38280 -6160
rect 38350 -6230 38370 -6160
rect 38440 -6230 38500 -6160
rect 31100 -6250 38500 -6230
rect 31100 -6320 38190 -6250
rect 38260 -6320 38280 -6250
rect 38350 -6320 38370 -6250
rect 38440 -6320 38500 -6250
rect 31100 -6340 38500 -6320
rect 31100 -6410 38190 -6340
rect 38260 -6410 38280 -6340
rect 38350 -6410 38370 -6340
rect 38440 -6410 38500 -6340
rect 31100 -6450 38500 -6410
rect 14520 -6510 16130 -6490
rect 14520 -6580 14700 -6510
rect 14770 -6580 14790 -6510
rect 14860 -6580 14880 -6510
rect 14950 -6580 14970 -6510
rect 15040 -6580 15060 -6510
rect 15130 -6580 15150 -6510
rect 15220 -6580 15240 -6510
rect 15310 -6580 15330 -6510
rect 15400 -6580 15420 -6510
rect 15490 -6580 15510 -6510
rect 15580 -6580 15600 -6510
rect 15670 -6580 15690 -6510
rect 15760 -6580 15780 -6510
rect 15850 -6580 15870 -6510
rect 15940 -6580 16130 -6510
rect 14520 -6640 16130 -6580
rect 16380 -6520 16520 -6470
rect 16380 -6590 16420 -6520
rect 16490 -6590 16520 -6520
rect 16380 -6630 16520 -6590
rect 16380 -6640 16420 -6630
rect 7560 -6720 7590 -6660
rect 7650 -6720 7690 -6660
rect 7750 -6720 7790 -6660
rect 7850 -6720 8490 -6660
rect 7560 -6760 8490 -6720
rect 7560 -6820 7590 -6760
rect 7650 -6820 7690 -6760
rect 7750 -6820 7790 -6760
rect 7850 -6820 8490 -6760
rect 7560 -6850 8490 -6820
rect 8710 -6670 16420 -6640
rect 8710 -6730 9870 -6670
rect 9930 -6730 9970 -6670
rect 10030 -6730 10070 -6670
rect 10130 -6700 16420 -6670
rect 16490 -6700 16520 -6630
rect 10130 -6730 16520 -6700
rect 8710 -6740 16520 -6730
rect 8710 -6770 16420 -6740
rect 8710 -6830 9870 -6770
rect 9930 -6830 9970 -6770
rect 10030 -6830 10070 -6770
rect 10130 -6810 16420 -6770
rect 16490 -6810 16520 -6740
rect 10130 -6830 16520 -6810
rect 8710 -6850 16520 -6830
rect -1740 -6920 -1710 -6850
rect -1640 -6870 6190 -6850
rect -1640 -6920 4770 -6870
rect -1740 -6930 4770 -6920
rect 4830 -6930 4870 -6870
rect 4930 -6930 4970 -6870
rect 5030 -6930 6190 -6870
rect -1740 -6950 6190 -6930
rect 0 -8140 310 -8120
rect 0 -8210 20 -8140
rect 90 -8210 130 -8140
rect 200 -8210 230 -8140
rect 300 -8210 310 -8140
rect 0 -8250 310 -8210
rect 0 -8320 20 -8250
rect 90 -8320 130 -8250
rect 200 -8320 230 -8250
rect 300 -8320 310 -8250
rect 0 -8360 310 -8320
rect 0 -8430 20 -8360
rect 90 -8430 130 -8360
rect 200 -8430 230 -8360
rect 300 -8430 310 -8360
rect 0 -8450 310 -8430
rect 5880 -9620 6190 -6950
rect -270 -9660 6190 -9620
rect -270 -9730 -240 -9660
rect -170 -9730 -130 -9660
rect -60 -9730 -20 -9660
rect 50 -9730 90 -9660
rect 160 -9730 6190 -9660
rect -270 -9790 6190 -9730
rect -270 -9860 -240 -9790
rect -170 -9860 -130 -9790
rect -60 -9860 -20 -9790
rect 50 -9860 90 -9790
rect 160 -9860 6190 -9790
rect -270 -9900 6190 -9860
rect 1080 -10340 2680 -10310
rect 1080 -10410 1150 -10340
rect 1220 -10410 1260 -10340
rect 1330 -10410 1370 -10340
rect 1440 -10410 1480 -10340
rect 1550 -10410 1590 -10340
rect 1660 -10410 1700 -10340
rect 1770 -10410 1810 -10340
rect 1880 -10410 1920 -10340
rect 1990 -10410 2030 -10340
rect 2100 -10410 2140 -10340
rect 2210 -10410 2250 -10340
rect 2320 -10410 2360 -10340
rect 2430 -10410 2470 -10340
rect 2540 -10410 2580 -10340
rect 2650 -10410 2680 -10340
rect 1080 -10450 2680 -10410
rect 1080 -10520 1150 -10450
rect 1220 -10520 1260 -10450
rect 1330 -10520 1370 -10450
rect 1440 -10520 1480 -10450
rect 1550 -10520 1590 -10450
rect 1660 -10520 1700 -10450
rect 1770 -10520 1810 -10450
rect 1880 -10520 1920 -10450
rect 1990 -10520 2030 -10450
rect 2100 -10520 2140 -10450
rect 2210 -10520 2250 -10450
rect 2320 -10520 2360 -10450
rect 2430 -10520 2470 -10450
rect 2540 -10520 2580 -10450
rect 2650 -10520 2680 -10450
rect 1080 -10570 2680 -10520
rect 1510 -12300 3110 -12250
rect 1510 -12370 1540 -12300
rect 1610 -12370 1650 -12300
rect 1720 -12370 1760 -12300
rect 1830 -12370 1870 -12300
rect 1940 -12370 1980 -12300
rect 2050 -12370 2090 -12300
rect 2160 -12370 2200 -12300
rect 2270 -12370 2310 -12300
rect 2380 -12370 2420 -12300
rect 2490 -12370 2530 -12300
rect 2600 -12370 2640 -12300
rect 2710 -12370 2750 -12300
rect 2820 -12370 2860 -12300
rect 2930 -12370 2970 -12300
rect 3040 -12370 3110 -12300
rect 1510 -12410 3110 -12370
rect 1510 -12480 1540 -12410
rect 1610 -12480 1650 -12410
rect 1720 -12480 1760 -12410
rect 1830 -12480 1870 -12410
rect 1940 -12480 1980 -12410
rect 2050 -12480 2090 -12410
rect 2160 -12480 2200 -12410
rect 2270 -12480 2310 -12410
rect 2380 -12480 2420 -12410
rect 2490 -12480 2530 -12410
rect 2600 -12480 2640 -12410
rect 2710 -12480 2750 -12410
rect 2820 -12480 2860 -12410
rect 2930 -12480 2970 -12410
rect 3040 -12480 3110 -12410
rect 1510 -12510 3110 -12480
rect 5880 -13220 6190 -9900
rect 8710 -6870 16420 -6850
rect 8710 -6930 9870 -6870
rect 9930 -6930 9970 -6870
rect 10030 -6930 10070 -6870
rect 10130 -6920 16420 -6870
rect 16490 -6920 16520 -6850
rect 10130 -6930 16520 -6920
rect 8710 -6950 16520 -6930
rect 8710 -9620 9020 -6950
rect 14590 -8230 14900 -8210
rect 14590 -8300 14600 -8230
rect 14670 -8300 14700 -8230
rect 14770 -8300 14810 -8230
rect 14880 -8300 14900 -8230
rect 14590 -8340 14900 -8300
rect 14590 -8410 14600 -8340
rect 14670 -8410 14700 -8340
rect 14770 -8410 14810 -8340
rect 14880 -8410 14900 -8340
rect 14590 -8450 14900 -8410
rect 14590 -8520 14600 -8450
rect 14670 -8520 14700 -8450
rect 14770 -8520 14810 -8450
rect 14880 -8520 14900 -8450
rect 14590 -8540 14900 -8520
rect 21610 -8360 21930 -8330
rect 21610 -8430 21630 -8360
rect 21700 -8430 21730 -8360
rect 21800 -8430 21830 -8360
rect 21900 -8430 21930 -8360
rect 21610 -8460 21930 -8430
rect 21610 -8530 21630 -8460
rect 21700 -8530 21730 -8460
rect 21800 -8530 21830 -8460
rect 21900 -8530 21930 -8460
rect 21610 -8560 21930 -8530
rect 21610 -8630 21630 -8560
rect 21700 -8630 21730 -8560
rect 21800 -8630 21830 -8560
rect 21900 -8630 21930 -8560
rect 21610 -8650 21930 -8630
rect 22630 -9010 22950 -8980
rect 22630 -9080 22650 -9010
rect 22720 -9080 22750 -9010
rect 22820 -9080 22850 -9010
rect 22920 -9080 22950 -9010
rect 22630 -9110 22950 -9080
rect 22630 -9180 22650 -9110
rect 22720 -9180 22750 -9110
rect 22820 -9180 22850 -9110
rect 22920 -9180 22950 -9110
rect 22630 -9210 22950 -9180
rect 22630 -9280 22650 -9210
rect 22720 -9280 22750 -9210
rect 22820 -9280 22850 -9210
rect 22920 -9280 22950 -9210
rect 22630 -9300 22950 -9280
rect 8710 -9660 15170 -9620
rect 8710 -9730 14720 -9660
rect 14790 -9730 14830 -9660
rect 14900 -9730 14940 -9660
rect 15010 -9730 15050 -9660
rect 15120 -9730 15170 -9660
rect 8710 -9790 15170 -9730
rect 8710 -9860 14720 -9790
rect 14790 -9860 14830 -9790
rect 14900 -9860 14940 -9790
rect 15010 -9860 15050 -9790
rect 15120 -9860 15170 -9790
rect 8710 -9900 15170 -9860
rect 8710 -13220 9020 -9900
rect 12220 -10370 13820 -10340
rect 12220 -10440 12290 -10370
rect 12360 -10440 12400 -10370
rect 12470 -10440 12510 -10370
rect 12580 -10440 12620 -10370
rect 12690 -10440 12730 -10370
rect 12800 -10440 12840 -10370
rect 12910 -10440 12950 -10370
rect 13020 -10440 13060 -10370
rect 13130 -10440 13170 -10370
rect 13240 -10440 13280 -10370
rect 13350 -10440 13390 -10370
rect 13460 -10440 13500 -10370
rect 13570 -10440 13610 -10370
rect 13680 -10440 13720 -10370
rect 13790 -10440 13820 -10370
rect 12220 -10480 13820 -10440
rect 12220 -10550 12290 -10480
rect 12360 -10550 12400 -10480
rect 12470 -10550 12510 -10480
rect 12580 -10550 12620 -10480
rect 12690 -10550 12730 -10480
rect 12800 -10550 12840 -10480
rect 12910 -10550 12950 -10480
rect 13020 -10550 13060 -10480
rect 13130 -10550 13170 -10480
rect 13240 -10550 13280 -10480
rect 13350 -10550 13390 -10480
rect 13460 -10550 13500 -10480
rect 13570 -10550 13610 -10480
rect 13680 -10550 13720 -10480
rect 13790 -10550 13820 -10480
rect 12220 -10600 13820 -10550
rect 29960 -10520 30790 -10510
rect 29960 -10590 29990 -10520
rect 30060 -10590 30700 -10520
rect 30770 -10590 30790 -10520
rect 29960 -10630 30790 -10590
rect 29960 -10700 29990 -10630
rect 30060 -10700 30700 -10630
rect 30770 -10700 30790 -10630
rect 29960 -10740 30790 -10700
rect 29960 -10810 29990 -10740
rect 30060 -10810 30700 -10740
rect 30770 -10810 30790 -10740
rect 29960 -10830 30790 -10810
rect 11790 -12300 13390 -12250
rect 11790 -12370 11820 -12300
rect 11890 -12370 11930 -12300
rect 12000 -12370 12040 -12300
rect 12110 -12370 12150 -12300
rect 12220 -12370 12260 -12300
rect 12330 -12370 12370 -12300
rect 12440 -12370 12480 -12300
rect 12550 -12370 12590 -12300
rect 12660 -12370 12700 -12300
rect 12770 -12370 12810 -12300
rect 12880 -12370 12920 -12300
rect 12990 -12370 13030 -12300
rect 13100 -12370 13140 -12300
rect 13210 -12370 13250 -12300
rect 13320 -12370 13390 -12300
rect 11790 -12410 13390 -12370
rect 11790 -12480 11820 -12410
rect 11890 -12480 11930 -12410
rect 12000 -12480 12040 -12410
rect 12110 -12480 12150 -12410
rect 12220 -12480 12260 -12410
rect 12330 -12480 12370 -12410
rect 12440 -12480 12480 -12410
rect 12550 -12480 12590 -12410
rect 12660 -12480 12700 -12410
rect 12770 -12480 12810 -12410
rect 12880 -12480 12920 -12410
rect 12990 -12480 13030 -12410
rect 13100 -12480 13140 -12410
rect 13210 -12480 13250 -12410
rect 13320 -12480 13390 -12410
rect 11790 -12510 13390 -12480
rect 5880 -13250 6610 -13220
rect 5880 -13310 6310 -13250
rect 6370 -13310 6410 -13250
rect 6470 -13310 6510 -13250
rect 6570 -13310 6610 -13250
rect 5880 -13340 6610 -13310
rect 5880 -13400 6310 -13340
rect 6370 -13400 6410 -13340
rect 6470 -13400 6510 -13340
rect 6570 -13400 6610 -13340
rect 5880 -13430 6610 -13400
rect 5880 -13490 6310 -13430
rect 6370 -13490 6410 -13430
rect 6470 -13490 6510 -13430
rect 6570 -13490 6610 -13430
rect 5880 -13530 6610 -13490
rect 5880 -13590 6310 -13530
rect 6370 -13590 6410 -13530
rect 6470 -13590 6510 -13530
rect 6570 -13590 6610 -13530
rect 5880 -13620 6610 -13590
rect 5880 -13680 6310 -13620
rect 6370 -13680 6410 -13620
rect 6470 -13680 6510 -13620
rect 6570 -13680 6610 -13620
rect 5880 -13710 6610 -13680
rect 5880 -13770 6310 -13710
rect 6370 -13770 6410 -13710
rect 6470 -13770 6510 -13710
rect 6570 -13770 6610 -13710
rect 5880 -13800 6610 -13770
rect 8290 -13250 9020 -13220
rect 8290 -13310 8330 -13250
rect 8390 -13310 8430 -13250
rect 8490 -13310 8530 -13250
rect 8590 -13310 9020 -13250
rect 8290 -13340 9020 -13310
rect 8290 -13400 8330 -13340
rect 8390 -13400 8430 -13340
rect 8490 -13400 8530 -13340
rect 8590 -13400 9020 -13340
rect 8290 -13430 9020 -13400
rect 8290 -13490 8330 -13430
rect 8390 -13490 8430 -13430
rect 8490 -13490 8530 -13430
rect 8590 -13490 9020 -13430
rect 8290 -13530 9020 -13490
rect 8290 -13590 8330 -13530
rect 8390 -13590 8430 -13530
rect 8490 -13590 8530 -13530
rect 8590 -13590 9020 -13530
rect 8290 -13620 9020 -13590
rect 8290 -13680 8330 -13620
rect 8390 -13680 8430 -13620
rect 8490 -13680 8530 -13620
rect 8590 -13680 9020 -13620
rect 8290 -13710 9020 -13680
rect 8290 -13770 8330 -13710
rect 8390 -13770 8430 -13710
rect 8490 -13770 8530 -13710
rect 8590 -13770 9020 -13710
rect 8290 -13800 9020 -13770
rect 21610 -14020 21930 -13990
rect 21610 -14090 21630 -14020
rect 21700 -14090 21730 -14020
rect 21800 -14090 21830 -14020
rect 21900 -14090 21930 -14020
rect 21610 -14120 21930 -14090
rect 21610 -14190 21630 -14120
rect 21700 -14190 21730 -14120
rect 21800 -14190 21830 -14120
rect 21900 -14190 21930 -14120
rect 21610 -14220 21930 -14190
rect 21610 -14290 21630 -14220
rect 21700 -14290 21730 -14220
rect 21800 -14290 21830 -14220
rect 21900 -14290 21930 -14220
rect 21610 -14310 21930 -14290
rect 22900 -14870 23220 -14840
rect 22900 -14940 22920 -14870
rect 22990 -14940 23020 -14870
rect 23090 -14940 23120 -14870
rect 23190 -14940 23220 -14870
rect 22900 -14970 23220 -14940
rect 22900 -15040 22920 -14970
rect 22990 -15040 23020 -14970
rect 23090 -15040 23120 -14970
rect 23190 -15040 23220 -14970
rect 22900 -15070 23220 -15040
rect 22900 -15140 22920 -15070
rect 22990 -15140 23020 -15070
rect 23090 -15140 23120 -15070
rect 23190 -15140 23220 -15070
rect 22900 -15160 23220 -15140
rect 4950 -17100 5270 -17070
rect 4950 -17160 4980 -17100
rect 5040 -17160 5080 -17100
rect 5140 -17160 5180 -17100
rect 5240 -17160 5270 -17100
rect 4950 -17200 5270 -17160
rect 4950 -17260 4980 -17200
rect 5040 -17260 5080 -17200
rect 5140 -17260 5180 -17200
rect 5240 -17260 5270 -17200
rect 4950 -17300 5270 -17260
rect 4950 -17360 4980 -17300
rect 5040 -17360 5080 -17300
rect 5140 -17360 5180 -17300
rect 5240 -17360 5270 -17300
rect 1550 -22660 3150 -22630
rect 1550 -22730 1620 -22660
rect 1690 -22730 1730 -22660
rect 1800 -22730 1840 -22660
rect 1910 -22730 1950 -22660
rect 2020 -22730 2060 -22660
rect 2130 -22730 2170 -22660
rect 2240 -22730 2280 -22660
rect 2350 -22730 2390 -22660
rect 2460 -22730 2500 -22660
rect 2570 -22730 2610 -22660
rect 2680 -22730 2720 -22660
rect 2790 -22730 2830 -22660
rect 2900 -22730 2940 -22660
rect 3010 -22730 3050 -22660
rect 3120 -22730 3150 -22660
rect 1550 -22770 3150 -22730
rect 1550 -22840 1620 -22770
rect 1690 -22840 1730 -22770
rect 1800 -22840 1840 -22770
rect 1910 -22840 1950 -22770
rect 2020 -22840 2060 -22770
rect 2130 -22840 2170 -22770
rect 2240 -22840 2280 -22770
rect 2350 -22840 2390 -22770
rect 2460 -22840 2500 -22770
rect 2570 -22840 2610 -22770
rect 2680 -22840 2720 -22770
rect 2790 -22840 2830 -22770
rect 2900 -22840 2940 -22770
rect 3010 -22840 3050 -22770
rect 3120 -22840 3150 -22770
rect 1550 -22890 3150 -22840
rect 4950 -24030 5270 -17360
rect 9630 -17100 9950 -17070
rect 9630 -17160 9660 -17100
rect 9720 -17160 9760 -17100
rect 9820 -17160 9860 -17100
rect 9920 -17160 9950 -17100
rect 9630 -17200 9950 -17160
rect 9630 -17260 9660 -17200
rect 9720 -17260 9760 -17200
rect 9820 -17260 9860 -17200
rect 9920 -17260 9950 -17200
rect 9630 -17300 9950 -17260
rect 9630 -17360 9660 -17300
rect 9720 -17360 9760 -17300
rect 9820 -17360 9860 -17300
rect 9920 -17360 9950 -17300
rect 6440 -17750 6750 -17730
rect 6440 -17820 6460 -17750
rect 6530 -17820 6560 -17750
rect 6630 -17820 6660 -17750
rect 6730 -17820 6750 -17750
rect 6440 -17860 6750 -17820
rect 6440 -17930 6460 -17860
rect 6530 -17930 6560 -17860
rect 6630 -17930 6660 -17860
rect 6730 -17930 6750 -17860
rect 6440 -17970 6750 -17930
rect 6440 -18040 6460 -17970
rect 6530 -18040 6560 -17970
rect 6630 -18040 6660 -17970
rect 6730 -18040 6750 -17970
rect 6440 -18080 6750 -18040
rect 6440 -18150 6460 -18080
rect 6530 -18150 6560 -18080
rect 6630 -18150 6660 -18080
rect 6730 -18150 6750 -18080
rect 6440 -18170 6750 -18150
rect 8150 -17750 8460 -17730
rect 8150 -17820 8170 -17750
rect 8240 -17820 8270 -17750
rect 8340 -17820 8370 -17750
rect 8440 -17820 8460 -17750
rect 8150 -17860 8460 -17820
rect 8150 -17930 8170 -17860
rect 8240 -17930 8270 -17860
rect 8340 -17930 8370 -17860
rect 8440 -17930 8460 -17860
rect 8150 -17970 8460 -17930
rect 8150 -18040 8170 -17970
rect 8240 -18040 8270 -17970
rect 8340 -18040 8370 -17970
rect 8440 -18040 8460 -17970
rect 8150 -18080 8460 -18040
rect 8150 -18150 8170 -18080
rect 8240 -18150 8270 -18080
rect 8340 -18150 8370 -18080
rect 8440 -18150 8460 -18080
rect 8150 -18170 8460 -18150
rect 9630 -24030 9950 -17360
rect 21610 -20100 21930 -20070
rect 21610 -20170 21630 -20100
rect 21700 -20170 21730 -20100
rect 21800 -20170 21830 -20100
rect 21900 -20170 21930 -20100
rect 21610 -20200 21930 -20170
rect 21610 -20270 21630 -20200
rect 21700 -20270 21730 -20200
rect 21800 -20270 21830 -20200
rect 21900 -20270 21930 -20200
rect 21610 -20300 21930 -20270
rect 21610 -20370 21630 -20300
rect 21700 -20370 21730 -20300
rect 21800 -20370 21830 -20300
rect 21900 -20370 21930 -20300
rect 21610 -20390 21930 -20370
rect 22680 -20730 23000 -20700
rect 22680 -20800 22700 -20730
rect 22770 -20800 22800 -20730
rect 22870 -20800 22900 -20730
rect 22970 -20800 23000 -20730
rect 22680 -20830 23000 -20800
rect 22680 -20900 22700 -20830
rect 22770 -20900 22800 -20830
rect 22870 -20900 22900 -20830
rect 22970 -20900 23000 -20830
rect 22680 -20930 23000 -20900
rect 22680 -21000 22700 -20930
rect 22770 -21000 22800 -20930
rect 22870 -21000 22900 -20930
rect 22970 -21000 23000 -20930
rect 22680 -21020 23000 -21000
rect 11750 -22660 13350 -22630
rect 11750 -22730 11820 -22660
rect 11890 -22730 11930 -22660
rect 12000 -22730 12040 -22660
rect 12110 -22730 12150 -22660
rect 12220 -22730 12260 -22660
rect 12330 -22730 12370 -22660
rect 12440 -22730 12480 -22660
rect 12550 -22730 12590 -22660
rect 12660 -22730 12700 -22660
rect 12770 -22730 12810 -22660
rect 12880 -22730 12920 -22660
rect 12990 -22730 13030 -22660
rect 13100 -22730 13140 -22660
rect 13210 -22730 13250 -22660
rect 13320 -22730 13350 -22660
rect 11750 -22770 13350 -22730
rect 11750 -22840 11820 -22770
rect 11890 -22840 11930 -22770
rect 12000 -22840 12040 -22770
rect 12110 -22840 12150 -22770
rect 12220 -22840 12260 -22770
rect 12330 -22840 12370 -22770
rect 12440 -22840 12480 -22770
rect 12550 -22840 12590 -22770
rect 12660 -22840 12700 -22770
rect 12770 -22840 12810 -22770
rect 12880 -22840 12920 -22770
rect 12990 -22840 13030 -22770
rect 13100 -22840 13140 -22770
rect 13210 -22840 13250 -22770
rect 13320 -22840 13350 -22770
rect 11750 -22890 13350 -22840
<< via3 >>
rect -5260 21510 -5190 21580
rect -5170 21510 -5100 21580
rect -5080 21510 -5010 21580
rect -4990 21510 -4920 21580
rect -4900 21510 -4830 21580
rect -4810 21510 -4740 21580
rect -4720 21510 -4650 21580
rect -4630 21510 -4560 21580
rect -4540 21510 -4470 21580
rect -4450 21510 -4380 21580
rect -4360 21510 -4290 21580
rect -4270 21510 -4200 21580
rect -4180 21510 -4110 21580
rect -4090 21510 -4020 21580
rect -4000 21510 -3930 21580
rect -3910 21510 -3840 21580
rect -3820 21510 -3750 21580
rect -3730 21510 -3660 21580
rect -3640 21510 -3570 21580
rect -3550 21510 -3480 21580
rect -3460 21510 -3390 21580
rect -3370 21510 -3300 21580
rect -3280 21510 -3210 21580
rect -3190 21510 -3120 21580
rect -3100 21510 -3030 21580
rect -3010 21510 -2940 21580
rect -2920 21510 -2850 21580
rect -2830 21510 -2760 21580
rect -2740 21510 -2670 21580
rect -2650 21510 -2580 21580
rect -2560 21510 -2490 21580
rect -2470 21510 -2400 21580
rect -2380 21510 -2310 21580
rect -2250 21510 -2180 21580
rect -2160 21510 -2090 21580
rect -2070 21510 -2000 21580
rect -1980 21510 -1910 21580
rect -1890 21510 -1820 21580
rect -1800 21510 -1730 21580
rect -1710 21510 -1640 21580
rect -1620 21510 -1550 21580
rect -1530 21510 -1460 21580
rect -1440 21510 -1370 21580
rect -1350 21510 -1280 21580
rect -1260 21510 -1190 21580
rect -1170 21510 -1100 21580
rect -1080 21510 -1010 21580
rect -990 21510 -920 21580
rect -900 21510 -830 21580
rect -810 21510 -740 21580
rect -720 21510 -650 21580
rect -630 21510 -560 21580
rect -540 21510 -470 21580
rect -450 21510 -380 21580
rect -360 21510 -290 21580
rect -270 21510 -200 21580
rect -180 21510 -110 21580
rect -90 21510 -20 21580
rect 0 21510 70 21580
rect 90 21510 160 21580
rect 180 21510 250 21580
rect 270 21510 340 21580
rect 360 21510 430 21580
rect 450 21510 520 21580
rect 540 21510 610 21580
rect 630 21510 700 21580
rect 760 21510 830 21580
rect 850 21510 920 21580
rect 940 21510 1010 21580
rect 1030 21510 1100 21580
rect 1120 21510 1190 21580
rect 1210 21510 1280 21580
rect 1300 21510 1370 21580
rect 1390 21510 1460 21580
rect 1480 21510 1550 21580
rect 1570 21510 1640 21580
rect 1660 21510 1730 21580
rect 1750 21510 1820 21580
rect 1840 21510 1910 21580
rect 1930 21510 2000 21580
rect 2020 21510 2090 21580
rect 2110 21510 2180 21580
rect 2200 21510 2270 21580
rect 2290 21510 2360 21580
rect 2380 21510 2450 21580
rect 2470 21510 2540 21580
rect 2560 21510 2630 21580
rect 2650 21510 2720 21580
rect 2740 21510 2810 21580
rect 2830 21510 2900 21580
rect 2920 21510 2990 21580
rect 3010 21510 3080 21580
rect 3100 21510 3170 21580
rect 3190 21510 3260 21580
rect 3280 21510 3350 21580
rect 3370 21510 3440 21580
rect 3460 21510 3530 21580
rect 3550 21510 3620 21580
rect 3640 21510 3710 21580
rect 3770 21510 3840 21580
rect 3860 21510 3930 21580
rect 3950 21510 4020 21580
rect 4040 21510 4110 21580
rect 4130 21510 4200 21580
rect 4220 21510 4290 21580
rect 4310 21510 4380 21580
rect 4400 21510 4470 21580
rect 4490 21510 4560 21580
rect 4580 21510 4650 21580
rect 4670 21510 4740 21580
rect 4760 21510 4830 21580
rect 4850 21510 4920 21580
rect 4940 21510 5010 21580
rect 5030 21510 5100 21580
rect 5120 21510 5190 21580
rect 5210 21510 5280 21580
rect 5300 21510 5370 21580
rect 5390 21510 5460 21580
rect 5480 21510 5550 21580
rect 5570 21510 5640 21580
rect 5660 21510 5730 21580
rect 5750 21510 5820 21580
rect 5840 21510 5910 21580
rect 5930 21510 6000 21580
rect 6020 21510 6090 21580
rect 6110 21510 6180 21580
rect 6200 21510 6270 21580
rect 6290 21510 6360 21580
rect 6380 21510 6450 21580
rect 6470 21510 6540 21580
rect 6560 21510 6630 21580
rect 6650 21510 6720 21580
rect -5260 21420 -5190 21490
rect -5170 21420 -5100 21490
rect -5080 21420 -5010 21490
rect -4990 21420 -4920 21490
rect -4900 21420 -4830 21490
rect -4810 21420 -4740 21490
rect -4720 21420 -4650 21490
rect -4630 21420 -4560 21490
rect -4540 21420 -4470 21490
rect -4450 21420 -4380 21490
rect -4360 21420 -4290 21490
rect -4270 21420 -4200 21490
rect -4180 21420 -4110 21490
rect -4090 21420 -4020 21490
rect -4000 21420 -3930 21490
rect -3910 21420 -3840 21490
rect -3820 21420 -3750 21490
rect -3730 21420 -3660 21490
rect -3640 21420 -3570 21490
rect -3550 21420 -3480 21490
rect -3460 21420 -3390 21490
rect -3370 21420 -3300 21490
rect -3280 21420 -3210 21490
rect -3190 21420 -3120 21490
rect -3100 21420 -3030 21490
rect -3010 21420 -2940 21490
rect -2920 21420 -2850 21490
rect -2830 21420 -2760 21490
rect -2740 21420 -2670 21490
rect -2650 21420 -2580 21490
rect -2560 21420 -2490 21490
rect -2470 21420 -2400 21490
rect -2380 21420 -2310 21490
rect -2250 21420 -2180 21490
rect -2160 21420 -2090 21490
rect -2070 21420 -2000 21490
rect -1980 21420 -1910 21490
rect -1890 21420 -1820 21490
rect -1800 21420 -1730 21490
rect -1710 21420 -1640 21490
rect -1620 21420 -1550 21490
rect -1530 21420 -1460 21490
rect -1440 21420 -1370 21490
rect -1350 21420 -1280 21490
rect -1260 21420 -1190 21490
rect -1170 21420 -1100 21490
rect -1080 21420 -1010 21490
rect -990 21420 -920 21490
rect -900 21420 -830 21490
rect -810 21420 -740 21490
rect -720 21420 -650 21490
rect -630 21420 -560 21490
rect -540 21420 -470 21490
rect -450 21420 -380 21490
rect -360 21420 -290 21490
rect -270 21420 -200 21490
rect -180 21420 -110 21490
rect -90 21420 -20 21490
rect 0 21420 70 21490
rect 90 21420 160 21490
rect 180 21420 250 21490
rect 270 21420 340 21490
rect 360 21420 430 21490
rect 450 21420 520 21490
rect 540 21420 610 21490
rect 630 21420 700 21490
rect 760 21420 830 21490
rect 850 21420 920 21490
rect 940 21420 1010 21490
rect 1030 21420 1100 21490
rect 1120 21420 1190 21490
rect 1210 21420 1280 21490
rect 1300 21420 1370 21490
rect 1390 21420 1460 21490
rect 1480 21420 1550 21490
rect 1570 21420 1640 21490
rect 1660 21420 1730 21490
rect 1750 21420 1820 21490
rect 1840 21420 1910 21490
rect 1930 21420 2000 21490
rect 2020 21420 2090 21490
rect 2110 21420 2180 21490
rect 2200 21420 2270 21490
rect 2290 21420 2360 21490
rect 2380 21420 2450 21490
rect 2470 21420 2540 21490
rect 2560 21420 2630 21490
rect 2650 21420 2720 21490
rect 2740 21420 2810 21490
rect 2830 21420 2900 21490
rect 2920 21420 2990 21490
rect 3010 21420 3080 21490
rect 3100 21420 3170 21490
rect 3190 21420 3260 21490
rect 3280 21420 3350 21490
rect 3370 21420 3440 21490
rect 3460 21420 3530 21490
rect 3550 21420 3620 21490
rect 3640 21420 3710 21490
rect 3770 21420 3840 21490
rect 3860 21420 3930 21490
rect 3950 21420 4020 21490
rect 4040 21420 4110 21490
rect 4130 21420 4200 21490
rect 4220 21420 4290 21490
rect 4310 21420 4380 21490
rect 4400 21420 4470 21490
rect 4490 21420 4560 21490
rect 4580 21420 4650 21490
rect 4670 21420 4740 21490
rect 4760 21420 4830 21490
rect 4850 21420 4920 21490
rect 4940 21420 5010 21490
rect 5030 21420 5100 21490
rect 5120 21420 5190 21490
rect 5210 21420 5280 21490
rect 5300 21420 5370 21490
rect 5390 21420 5460 21490
rect 5480 21420 5550 21490
rect 5570 21420 5640 21490
rect 5660 21420 5730 21490
rect 5750 21420 5820 21490
rect 5840 21420 5910 21490
rect 5930 21420 6000 21490
rect 6020 21420 6090 21490
rect 6110 21420 6180 21490
rect 6200 21420 6270 21490
rect 6290 21420 6360 21490
rect 6380 21420 6450 21490
rect 6470 21420 6540 21490
rect 6560 21420 6630 21490
rect 6650 21420 6720 21490
rect -5260 21330 -5190 21400
rect -5170 21330 -5100 21400
rect -5080 21330 -5010 21400
rect -4990 21330 -4920 21400
rect -4900 21330 -4830 21400
rect -4810 21330 -4740 21400
rect -4720 21330 -4650 21400
rect -4630 21330 -4560 21400
rect -4540 21330 -4470 21400
rect -4450 21330 -4380 21400
rect -4360 21330 -4290 21400
rect -4270 21330 -4200 21400
rect -4180 21330 -4110 21400
rect -4090 21330 -4020 21400
rect -4000 21330 -3930 21400
rect -3910 21330 -3840 21400
rect -3820 21330 -3750 21400
rect -3730 21330 -3660 21400
rect -3640 21330 -3570 21400
rect -3550 21330 -3480 21400
rect -3460 21330 -3390 21400
rect -3370 21330 -3300 21400
rect -3280 21330 -3210 21400
rect -3190 21330 -3120 21400
rect -3100 21330 -3030 21400
rect -3010 21330 -2940 21400
rect -2920 21330 -2850 21400
rect -2830 21330 -2760 21400
rect -2740 21330 -2670 21400
rect -2650 21330 -2580 21400
rect -2560 21330 -2490 21400
rect -2470 21330 -2400 21400
rect -2380 21330 -2310 21400
rect -2250 21330 -2180 21400
rect -2160 21330 -2090 21400
rect -2070 21330 -2000 21400
rect -1980 21330 -1910 21400
rect -1890 21330 -1820 21400
rect -1800 21330 -1730 21400
rect -1710 21330 -1640 21400
rect -1620 21330 -1550 21400
rect -1530 21330 -1460 21400
rect -1440 21330 -1370 21400
rect -1350 21330 -1280 21400
rect -1260 21330 -1190 21400
rect -1170 21330 -1100 21400
rect -1080 21330 -1010 21400
rect -990 21330 -920 21400
rect -900 21330 -830 21400
rect -810 21330 -740 21400
rect -720 21330 -650 21400
rect -630 21330 -560 21400
rect -540 21330 -470 21400
rect -450 21330 -380 21400
rect -360 21330 -290 21400
rect -270 21330 -200 21400
rect -180 21330 -110 21400
rect -90 21330 -20 21400
rect 0 21330 70 21400
rect 90 21330 160 21400
rect 180 21330 250 21400
rect 270 21330 340 21400
rect 360 21330 430 21400
rect 450 21330 520 21400
rect 540 21330 610 21400
rect 630 21330 700 21400
rect 760 21330 830 21400
rect 850 21330 920 21400
rect 940 21330 1010 21400
rect 1030 21330 1100 21400
rect 1120 21330 1190 21400
rect 1210 21330 1280 21400
rect 1300 21330 1370 21400
rect 1390 21330 1460 21400
rect 1480 21330 1550 21400
rect 1570 21330 1640 21400
rect 1660 21330 1730 21400
rect 1750 21330 1820 21400
rect 1840 21330 1910 21400
rect 1930 21330 2000 21400
rect 2020 21330 2090 21400
rect 2110 21330 2180 21400
rect 2200 21330 2270 21400
rect 2290 21330 2360 21400
rect 2380 21330 2450 21400
rect 2470 21330 2540 21400
rect 2560 21330 2630 21400
rect 2650 21330 2720 21400
rect 2740 21330 2810 21400
rect 2830 21330 2900 21400
rect 2920 21330 2990 21400
rect 3010 21330 3080 21400
rect 3100 21330 3170 21400
rect 3190 21330 3260 21400
rect 3280 21330 3350 21400
rect 3370 21330 3440 21400
rect 3460 21330 3530 21400
rect 3550 21330 3620 21400
rect 3640 21330 3710 21400
rect 3770 21330 3840 21400
rect 3860 21330 3930 21400
rect 3950 21330 4020 21400
rect 4040 21330 4110 21400
rect 4130 21330 4200 21400
rect 4220 21330 4290 21400
rect 4310 21330 4380 21400
rect 4400 21330 4470 21400
rect 4490 21330 4560 21400
rect 4580 21330 4650 21400
rect 4670 21330 4740 21400
rect 4760 21330 4830 21400
rect 4850 21330 4920 21400
rect 4940 21330 5010 21400
rect 5030 21330 5100 21400
rect 5120 21330 5190 21400
rect 5210 21330 5280 21400
rect 5300 21330 5370 21400
rect 5390 21330 5460 21400
rect 5480 21330 5550 21400
rect 5570 21330 5640 21400
rect 5660 21330 5730 21400
rect 5750 21330 5820 21400
rect 5840 21330 5910 21400
rect 5930 21330 6000 21400
rect 6020 21330 6090 21400
rect 6110 21330 6180 21400
rect 6200 21330 6270 21400
rect 6290 21330 6360 21400
rect 6380 21330 6450 21400
rect 6470 21330 6540 21400
rect 6560 21330 6630 21400
rect 6650 21330 6720 21400
rect 8180 21510 8250 21580
rect 8270 21510 8340 21580
rect 8360 21510 8430 21580
rect 8450 21510 8520 21580
rect 8540 21510 8610 21580
rect 8630 21510 8700 21580
rect 8720 21510 8790 21580
rect 8810 21510 8880 21580
rect 8900 21510 8970 21580
rect 8990 21510 9060 21580
rect 9080 21510 9150 21580
rect 9170 21510 9240 21580
rect 9260 21510 9330 21580
rect 9350 21510 9420 21580
rect 9440 21510 9510 21580
rect 9530 21510 9600 21580
rect 9620 21510 9690 21580
rect 9710 21510 9780 21580
rect 9800 21510 9870 21580
rect 9890 21510 9960 21580
rect 9980 21510 10050 21580
rect 10070 21510 10140 21580
rect 10160 21510 10230 21580
rect 10250 21510 10320 21580
rect 10340 21510 10410 21580
rect 10430 21510 10500 21580
rect 10520 21510 10590 21580
rect 10610 21510 10680 21580
rect 10700 21510 10770 21580
rect 10790 21510 10860 21580
rect 10880 21510 10950 21580
rect 10970 21510 11040 21580
rect 11060 21510 11130 21580
rect 11190 21510 11260 21580
rect 11280 21510 11350 21580
rect 11370 21510 11440 21580
rect 11460 21510 11530 21580
rect 11550 21510 11620 21580
rect 11640 21510 11710 21580
rect 11730 21510 11800 21580
rect 11820 21510 11890 21580
rect 11910 21510 11980 21580
rect 12000 21510 12070 21580
rect 12090 21510 12160 21580
rect 12180 21510 12250 21580
rect 12270 21510 12340 21580
rect 12360 21510 12430 21580
rect 12450 21510 12520 21580
rect 12540 21510 12610 21580
rect 12630 21510 12700 21580
rect 12720 21510 12790 21580
rect 12810 21510 12880 21580
rect 12900 21510 12970 21580
rect 12990 21510 13060 21580
rect 13080 21510 13150 21580
rect 13170 21510 13240 21580
rect 13260 21510 13330 21580
rect 13350 21510 13420 21580
rect 13440 21510 13510 21580
rect 13530 21510 13600 21580
rect 13620 21510 13690 21580
rect 13710 21510 13780 21580
rect 13800 21510 13870 21580
rect 13890 21510 13960 21580
rect 13980 21510 14050 21580
rect 14070 21510 14140 21580
rect 14200 21510 14270 21580
rect 14290 21510 14360 21580
rect 14380 21510 14450 21580
rect 14470 21510 14540 21580
rect 14560 21510 14630 21580
rect 14650 21510 14720 21580
rect 14740 21510 14810 21580
rect 14830 21510 14900 21580
rect 14920 21510 14990 21580
rect 15010 21510 15080 21580
rect 15100 21510 15170 21580
rect 15190 21510 15260 21580
rect 15280 21510 15350 21580
rect 15370 21510 15440 21580
rect 15460 21510 15530 21580
rect 15550 21510 15620 21580
rect 15640 21510 15710 21580
rect 15730 21510 15800 21580
rect 15820 21510 15890 21580
rect 15910 21510 15980 21580
rect 16000 21510 16070 21580
rect 16090 21510 16160 21580
rect 16180 21510 16250 21580
rect 16270 21510 16340 21580
rect 16360 21510 16430 21580
rect 16450 21510 16520 21580
rect 16540 21510 16610 21580
rect 16630 21510 16700 21580
rect 16720 21510 16790 21580
rect 16810 21510 16880 21580
rect 16900 21510 16970 21580
rect 16990 21510 17060 21580
rect 17080 21510 17150 21580
rect 17210 21510 17280 21580
rect 17300 21510 17370 21580
rect 17390 21510 17460 21580
rect 17480 21510 17550 21580
rect 17570 21510 17640 21580
rect 17660 21510 17730 21580
rect 17750 21510 17820 21580
rect 17840 21510 17910 21580
rect 17930 21510 18000 21580
rect 18020 21510 18090 21580
rect 18110 21510 18180 21580
rect 18200 21510 18270 21580
rect 18290 21510 18360 21580
rect 18380 21510 18450 21580
rect 18470 21510 18540 21580
rect 18560 21510 18630 21580
rect 18650 21510 18720 21580
rect 18740 21510 18810 21580
rect 18830 21510 18900 21580
rect 18920 21510 18990 21580
rect 19010 21510 19080 21580
rect 19100 21510 19170 21580
rect 19190 21510 19260 21580
rect 19280 21510 19350 21580
rect 19370 21510 19440 21580
rect 19460 21510 19530 21580
rect 19550 21510 19620 21580
rect 19640 21510 19710 21580
rect 19730 21510 19800 21580
rect 19820 21510 19890 21580
rect 19910 21510 19980 21580
rect 20000 21510 20070 21580
rect 20090 21510 20160 21580
rect 8180 21420 8250 21490
rect 8270 21420 8340 21490
rect 8360 21420 8430 21490
rect 8450 21420 8520 21490
rect 8540 21420 8610 21490
rect 8630 21420 8700 21490
rect 8720 21420 8790 21490
rect 8810 21420 8880 21490
rect 8900 21420 8970 21490
rect 8990 21420 9060 21490
rect 9080 21420 9150 21490
rect 9170 21420 9240 21490
rect 9260 21420 9330 21490
rect 9350 21420 9420 21490
rect 9440 21420 9510 21490
rect 9530 21420 9600 21490
rect 9620 21420 9690 21490
rect 9710 21420 9780 21490
rect 9800 21420 9870 21490
rect 9890 21420 9960 21490
rect 9980 21420 10050 21490
rect 10070 21420 10140 21490
rect 10160 21420 10230 21490
rect 10250 21420 10320 21490
rect 10340 21420 10410 21490
rect 10430 21420 10500 21490
rect 10520 21420 10590 21490
rect 10610 21420 10680 21490
rect 10700 21420 10770 21490
rect 10790 21420 10860 21490
rect 10880 21420 10950 21490
rect 10970 21420 11040 21490
rect 11060 21420 11130 21490
rect 11190 21420 11260 21490
rect 11280 21420 11350 21490
rect 11370 21420 11440 21490
rect 11460 21420 11530 21490
rect 11550 21420 11620 21490
rect 11640 21420 11710 21490
rect 11730 21420 11800 21490
rect 11820 21420 11890 21490
rect 11910 21420 11980 21490
rect 12000 21420 12070 21490
rect 12090 21420 12160 21490
rect 12180 21420 12250 21490
rect 12270 21420 12340 21490
rect 12360 21420 12430 21490
rect 12450 21420 12520 21490
rect 12540 21420 12610 21490
rect 12630 21420 12700 21490
rect 12720 21420 12790 21490
rect 12810 21420 12880 21490
rect 12900 21420 12970 21490
rect 12990 21420 13060 21490
rect 13080 21420 13150 21490
rect 13170 21420 13240 21490
rect 13260 21420 13330 21490
rect 13350 21420 13420 21490
rect 13440 21420 13510 21490
rect 13530 21420 13600 21490
rect 13620 21420 13690 21490
rect 13710 21420 13780 21490
rect 13800 21420 13870 21490
rect 13890 21420 13960 21490
rect 13980 21420 14050 21490
rect 14070 21420 14140 21490
rect 14200 21420 14270 21490
rect 14290 21420 14360 21490
rect 14380 21420 14450 21490
rect 14470 21420 14540 21490
rect 14560 21420 14630 21490
rect 14650 21420 14720 21490
rect 14740 21420 14810 21490
rect 14830 21420 14900 21490
rect 14920 21420 14990 21490
rect 15010 21420 15080 21490
rect 15100 21420 15170 21490
rect 15190 21420 15260 21490
rect 15280 21420 15350 21490
rect 15370 21420 15440 21490
rect 15460 21420 15530 21490
rect 15550 21420 15620 21490
rect 15640 21420 15710 21490
rect 15730 21420 15800 21490
rect 15820 21420 15890 21490
rect 15910 21420 15980 21490
rect 16000 21420 16070 21490
rect 16090 21420 16160 21490
rect 16180 21420 16250 21490
rect 16270 21420 16340 21490
rect 16360 21420 16430 21490
rect 16450 21420 16520 21490
rect 16540 21420 16610 21490
rect 16630 21420 16700 21490
rect 16720 21420 16790 21490
rect 16810 21420 16880 21490
rect 16900 21420 16970 21490
rect 16990 21420 17060 21490
rect 17080 21420 17150 21490
rect 17210 21420 17280 21490
rect 17300 21420 17370 21490
rect 17390 21420 17460 21490
rect 17480 21420 17550 21490
rect 17570 21420 17640 21490
rect 17660 21420 17730 21490
rect 17750 21420 17820 21490
rect 17840 21420 17910 21490
rect 17930 21420 18000 21490
rect 18020 21420 18090 21490
rect 18110 21420 18180 21490
rect 18200 21420 18270 21490
rect 18290 21420 18360 21490
rect 18380 21420 18450 21490
rect 18470 21420 18540 21490
rect 18560 21420 18630 21490
rect 18650 21420 18720 21490
rect 18740 21420 18810 21490
rect 18830 21420 18900 21490
rect 18920 21420 18990 21490
rect 19010 21420 19080 21490
rect 19100 21420 19170 21490
rect 19190 21420 19260 21490
rect 19280 21420 19350 21490
rect 19370 21420 19440 21490
rect 19460 21420 19530 21490
rect 19550 21420 19620 21490
rect 19640 21420 19710 21490
rect 19730 21420 19800 21490
rect 19820 21420 19890 21490
rect 19910 21420 19980 21490
rect 20000 21420 20070 21490
rect 20090 21420 20160 21490
rect 8180 21330 8250 21400
rect 8270 21330 8340 21400
rect 8360 21330 8430 21400
rect 8450 21330 8520 21400
rect 8540 21330 8610 21400
rect 8630 21330 8700 21400
rect 8720 21330 8790 21400
rect 8810 21330 8880 21400
rect 8900 21330 8970 21400
rect 8990 21330 9060 21400
rect 9080 21330 9150 21400
rect 9170 21330 9240 21400
rect 9260 21330 9330 21400
rect 9350 21330 9420 21400
rect 9440 21330 9510 21400
rect 9530 21330 9600 21400
rect 9620 21330 9690 21400
rect 9710 21330 9780 21400
rect 9800 21330 9870 21400
rect 9890 21330 9960 21400
rect 9980 21330 10050 21400
rect 10070 21330 10140 21400
rect 10160 21330 10230 21400
rect 10250 21330 10320 21400
rect 10340 21330 10410 21400
rect 10430 21330 10500 21400
rect 10520 21330 10590 21400
rect 10610 21330 10680 21400
rect 10700 21330 10770 21400
rect 10790 21330 10860 21400
rect 10880 21330 10950 21400
rect 10970 21330 11040 21400
rect 11060 21330 11130 21400
rect 11190 21330 11260 21400
rect 11280 21330 11350 21400
rect 11370 21330 11440 21400
rect 11460 21330 11530 21400
rect 11550 21330 11620 21400
rect 11640 21330 11710 21400
rect 11730 21330 11800 21400
rect 11820 21330 11890 21400
rect 11910 21330 11980 21400
rect 12000 21330 12070 21400
rect 12090 21330 12160 21400
rect 12180 21330 12250 21400
rect 12270 21330 12340 21400
rect 12360 21330 12430 21400
rect 12450 21330 12520 21400
rect 12540 21330 12610 21400
rect 12630 21330 12700 21400
rect 12720 21330 12790 21400
rect 12810 21330 12880 21400
rect 12900 21330 12970 21400
rect 12990 21330 13060 21400
rect 13080 21330 13150 21400
rect 13170 21330 13240 21400
rect 13260 21330 13330 21400
rect 13350 21330 13420 21400
rect 13440 21330 13510 21400
rect 13530 21330 13600 21400
rect 13620 21330 13690 21400
rect 13710 21330 13780 21400
rect 13800 21330 13870 21400
rect 13890 21330 13960 21400
rect 13980 21330 14050 21400
rect 14070 21330 14140 21400
rect 14200 21330 14270 21400
rect 14290 21330 14360 21400
rect 14380 21330 14450 21400
rect 14470 21330 14540 21400
rect 14560 21330 14630 21400
rect 14650 21330 14720 21400
rect 14740 21330 14810 21400
rect 14830 21330 14900 21400
rect 14920 21330 14990 21400
rect 15010 21330 15080 21400
rect 15100 21330 15170 21400
rect 15190 21330 15260 21400
rect 15280 21330 15350 21400
rect 15370 21330 15440 21400
rect 15460 21330 15530 21400
rect 15550 21330 15620 21400
rect 15640 21330 15710 21400
rect 15730 21330 15800 21400
rect 15820 21330 15890 21400
rect 15910 21330 15980 21400
rect 16000 21330 16070 21400
rect 16090 21330 16160 21400
rect 16180 21330 16250 21400
rect 16270 21330 16340 21400
rect 16360 21330 16430 21400
rect 16450 21330 16520 21400
rect 16540 21330 16610 21400
rect 16630 21330 16700 21400
rect 16720 21330 16790 21400
rect 16810 21330 16880 21400
rect 16900 21330 16970 21400
rect 16990 21330 17060 21400
rect 17080 21330 17150 21400
rect 17210 21330 17280 21400
rect 17300 21330 17370 21400
rect 17390 21330 17460 21400
rect 17480 21330 17550 21400
rect 17570 21330 17640 21400
rect 17660 21330 17730 21400
rect 17750 21330 17820 21400
rect 17840 21330 17910 21400
rect 17930 21330 18000 21400
rect 18020 21330 18090 21400
rect 18110 21330 18180 21400
rect 18200 21330 18270 21400
rect 18290 21330 18360 21400
rect 18380 21330 18450 21400
rect 18470 21330 18540 21400
rect 18560 21330 18630 21400
rect 18650 21330 18720 21400
rect 18740 21330 18810 21400
rect 18830 21330 18900 21400
rect 18920 21330 18990 21400
rect 19010 21330 19080 21400
rect 19100 21330 19170 21400
rect 19190 21330 19260 21400
rect 19280 21330 19350 21400
rect 19370 21330 19440 21400
rect 19460 21330 19530 21400
rect 19550 21330 19620 21400
rect 19640 21330 19710 21400
rect 19730 21330 19800 21400
rect 19820 21330 19890 21400
rect 19910 21330 19980 21400
rect 20000 21330 20070 21400
rect 20090 21330 20160 21400
rect 6470 8340 6540 8410
rect 6560 8340 6630 8410
rect 6650 8340 6720 8410
rect 6470 8250 6540 8320
rect 6560 8250 6630 8320
rect 6650 8250 6720 8320
rect 1570 6780 1640 6850
rect 1680 6780 1750 6850
rect 1790 6780 1860 6850
rect 1900 6780 1970 6850
rect 2010 6780 2080 6850
rect 2120 6780 2190 6850
rect 2230 6780 2300 6850
rect 2340 6780 2410 6850
rect 2450 6780 2520 6850
rect 2560 6780 2630 6850
rect 2670 6780 2740 6850
rect 2780 6780 2850 6850
rect 2890 6780 2960 6850
rect 3000 6780 3070 6850
rect 1570 6670 1640 6740
rect 1680 6670 1750 6740
rect 1790 6670 1860 6740
rect 1900 6670 1970 6740
rect 2010 6670 2080 6740
rect 2120 6670 2190 6740
rect 2230 6670 2300 6740
rect 2340 6670 2410 6740
rect 2450 6670 2520 6740
rect 2560 6670 2630 6740
rect 2670 6670 2740 6740
rect 2780 6670 2850 6740
rect 2890 6670 2960 6740
rect 3000 6670 3070 6740
rect 8180 8340 8250 8410
rect 8270 8340 8340 8410
rect 8360 8340 8430 8410
rect 8180 8250 8250 8320
rect 8270 8250 8340 8320
rect 8360 8250 8430 8320
rect 7410 5320 7480 5390
rect 7410 5210 7480 5280
rect 7410 5100 7480 5170
rect 7410 4990 7480 5060
rect 7410 4880 7480 4950
rect 38190 7750 38260 7820
rect 38280 7750 38350 7820
rect 38370 7750 38440 7820
rect 38190 7660 38260 7730
rect 38280 7660 38350 7730
rect 38370 7660 38440 7730
rect 38190 7570 38260 7640
rect 38280 7570 38350 7640
rect 38370 7570 38440 7640
rect 38190 7480 38260 7550
rect 38280 7480 38350 7550
rect 38370 7480 38440 7550
rect 38190 7390 38260 7460
rect 38280 7390 38350 7460
rect 38370 7390 38440 7460
rect 38190 7300 38260 7370
rect 38280 7300 38350 7370
rect 38370 7300 38440 7370
rect 23490 7140 23560 7210
rect 23600 7140 23670 7210
rect 23710 7140 23780 7210
rect 23820 7140 23890 7210
rect 23490 7030 23560 7100
rect 23600 7030 23670 7100
rect 23710 7030 23780 7100
rect 23820 7030 23890 7100
rect 25890 7140 25960 7210
rect 26000 7140 26070 7210
rect 26110 7140 26180 7210
rect 26220 7140 26290 7210
rect 25890 7030 25960 7100
rect 26000 7030 26070 7100
rect 26110 7030 26180 7100
rect 26220 7030 26290 7100
rect 38190 7210 38260 7280
rect 38280 7210 38350 7280
rect 38370 7210 38440 7280
rect 38190 7080 38260 7150
rect 38280 7080 38350 7150
rect 38370 7080 38440 7150
rect 38190 6990 38260 7060
rect 38280 6990 38350 7060
rect 38370 6990 38440 7060
rect 11790 6810 11860 6880
rect 11900 6810 11970 6880
rect 12010 6810 12080 6880
rect 12120 6810 12190 6880
rect 12230 6810 12300 6880
rect 12340 6810 12410 6880
rect 12450 6810 12520 6880
rect 12560 6810 12630 6880
rect 12670 6810 12740 6880
rect 12780 6810 12850 6880
rect 12890 6810 12960 6880
rect 13000 6810 13070 6880
rect 13110 6810 13180 6880
rect 13220 6810 13290 6880
rect 11790 6700 11860 6770
rect 11900 6700 11970 6770
rect 12010 6700 12080 6770
rect 12120 6700 12190 6770
rect 12230 6700 12300 6770
rect 12340 6700 12410 6770
rect 12450 6700 12520 6770
rect 12560 6700 12630 6770
rect 12670 6700 12740 6770
rect 12780 6700 12850 6770
rect 12890 6700 12960 6770
rect 13000 6700 13070 6770
rect 13110 6700 13180 6770
rect 13220 6700 13290 6770
rect 38190 6900 38260 6970
rect 38280 6900 38350 6970
rect 38370 6900 38440 6970
rect 38190 6810 38260 6880
rect 38280 6810 38350 6880
rect 38370 6810 38440 6880
rect 38190 6720 38260 6790
rect 38280 6720 38350 6790
rect 38370 6720 38440 6790
rect 38190 6630 38260 6700
rect 38280 6630 38350 6700
rect 38370 6630 38440 6700
rect 38190 6540 38260 6610
rect 38280 6540 38350 6610
rect 38370 6540 38440 6610
rect 38190 6450 38260 6520
rect 38280 6450 38350 6520
rect 38370 6450 38440 6520
rect 38190 6360 38260 6430
rect 38280 6360 38350 6430
rect 38370 6360 38440 6430
rect 30740 6230 30810 6300
rect 30850 6230 30920 6300
rect 30740 6100 30810 6170
rect 30850 6100 30920 6170
rect 30740 5970 30810 6040
rect 30850 5970 30920 6040
rect 38190 6270 38260 6340
rect 38280 6270 38350 6340
rect 38370 6270 38440 6340
rect 38190 6180 38260 6250
rect 38280 6180 38350 6250
rect 38370 6180 38440 6250
rect 38190 6090 38260 6160
rect 38280 6090 38350 6160
rect 38370 6090 38440 6160
rect 38190 6000 38260 6070
rect 38280 6000 38350 6070
rect 38370 6000 38440 6070
rect 38190 5910 38260 5980
rect 38280 5910 38350 5980
rect 38370 5910 38440 5980
rect 38190 5820 38260 5890
rect 38280 5820 38350 5890
rect 38370 5820 38440 5890
rect 38190 5730 38260 5800
rect 38280 5730 38350 5800
rect 38370 5730 38440 5800
rect 21820 5600 21890 5670
rect 21930 5600 22000 5670
rect 21820 5490 21890 5560
rect 21930 5490 22000 5560
rect 21820 5380 21890 5450
rect 21930 5380 22000 5450
rect 21820 5270 21890 5340
rect 21930 5270 22000 5340
rect 21820 5160 21890 5230
rect 21930 5160 22000 5230
rect 21820 5050 21890 5120
rect 21930 5050 22000 5120
rect 21820 4940 21890 5010
rect 21930 4940 22000 5010
rect 21820 4830 21890 4900
rect 21930 4830 22000 4900
rect 21820 4720 21890 4790
rect 21930 4720 22000 4790
rect 21820 4610 21890 4680
rect 21930 4610 22000 4680
rect 21820 4500 21890 4570
rect 21930 4500 22000 4570
rect 38190 5640 38260 5710
rect 38280 5640 38350 5710
rect 38370 5640 38440 5710
rect 38190 5550 38260 5620
rect 38280 5550 38350 5620
rect 38370 5550 38440 5620
rect 38190 5460 38260 5530
rect 38280 5460 38350 5530
rect 38370 5460 38440 5530
rect 38190 5370 38260 5440
rect 38280 5370 38350 5440
rect 38370 5370 38440 5440
rect 38190 5280 38260 5350
rect 38280 5280 38350 5350
rect 38370 5280 38440 5350
rect 38190 5190 38260 5260
rect 38280 5190 38350 5260
rect 38370 5190 38440 5260
rect 38190 5100 38260 5170
rect 38280 5100 38350 5170
rect 38370 5100 38440 5170
rect 38190 5010 38260 5080
rect 38280 5010 38350 5080
rect 38370 5010 38440 5080
rect 38190 4920 38260 4990
rect 38280 4920 38350 4990
rect 38370 4920 38440 4990
rect 38190 4830 38260 4900
rect 38280 4830 38350 4900
rect 38370 4830 38440 4900
rect 38190 4740 38260 4810
rect 38280 4740 38350 4810
rect 38370 4740 38440 4810
rect 38190 4650 38260 4720
rect 38280 4650 38350 4720
rect 38370 4650 38440 4720
rect 38190 4560 38260 4630
rect 38280 4560 38350 4630
rect 38370 4560 38440 4630
rect 38190 4470 38260 4540
rect 38280 4470 38350 4540
rect 38370 4470 38440 4540
rect 38190 4380 38260 4450
rect 38280 4380 38350 4450
rect 38370 4380 38440 4450
rect 38190 4290 38260 4360
rect 38280 4290 38350 4360
rect 38370 4290 38440 4360
rect 38190 4200 38260 4270
rect 38280 4200 38350 4270
rect 38370 4200 38440 4270
rect 38190 4070 38260 4140
rect 38280 4070 38350 4140
rect 38370 4070 38440 4140
rect 38190 3980 38260 4050
rect 38280 3980 38350 4050
rect 38370 3980 38440 4050
rect 38190 3890 38260 3960
rect 38280 3890 38350 3960
rect 38370 3890 38440 3960
rect 38190 3800 38260 3870
rect 38280 3800 38350 3870
rect 38370 3800 38440 3870
rect 38190 3710 38260 3780
rect 38280 3710 38350 3780
rect 38370 3710 38440 3780
rect 38190 3620 38260 3690
rect 38280 3620 38350 3690
rect 38370 3620 38440 3690
rect 38190 3530 38260 3600
rect 38280 3530 38350 3600
rect 38370 3530 38440 3600
rect 38190 3440 38260 3510
rect 38280 3440 38350 3510
rect 38370 3440 38440 3510
rect 24720 3290 24790 3360
rect 24830 3290 24900 3360
rect 24940 3290 25010 3360
rect 24720 3180 24790 3250
rect 24830 3180 24900 3250
rect 24940 3180 25010 3250
rect 24720 3070 24790 3140
rect 24830 3070 24900 3140
rect 24940 3070 25010 3140
rect 38190 3350 38260 3420
rect 38280 3350 38350 3420
rect 38370 3350 38440 3420
rect 38190 3260 38260 3330
rect 38280 3260 38350 3330
rect 38370 3260 38440 3330
rect 38190 3170 38260 3240
rect 38280 3170 38350 3240
rect 38370 3170 38440 3240
rect 38190 3080 38260 3150
rect 38280 3080 38350 3150
rect 38370 3080 38440 3150
rect 38190 2990 38260 3060
rect 38280 2990 38350 3060
rect 38370 2990 38440 3060
rect 1150 -860 1220 -790
rect 1260 -860 1330 -790
rect 1370 -860 1440 -790
rect 1480 -860 1550 -790
rect 1590 -860 1660 -790
rect 1700 -860 1770 -790
rect 1810 -860 1880 -790
rect 1920 -860 1990 -790
rect 2030 -860 2100 -790
rect 2140 -860 2210 -790
rect 2250 -860 2320 -790
rect 2360 -860 2430 -790
rect 2470 -860 2540 -790
rect 2580 -860 2650 -790
rect 1150 -970 1220 -900
rect 1260 -970 1330 -900
rect 1370 -970 1440 -900
rect 1480 -970 1550 -900
rect 1590 -970 1660 -900
rect 1700 -970 1770 -900
rect 1810 -970 1880 -900
rect 1920 -970 1990 -900
rect 2030 -970 2100 -900
rect 2140 -970 2210 -900
rect 2250 -970 2320 -900
rect 2360 -970 2430 -900
rect 2470 -970 2540 -900
rect 2580 -970 2650 -900
rect 1570 -2850 1640 -2780
rect 1680 -2850 1750 -2780
rect 1790 -2850 1860 -2780
rect 1900 -2850 1970 -2780
rect 2010 -2850 2080 -2780
rect 2120 -2850 2190 -2780
rect 2230 -2850 2300 -2780
rect 2340 -2850 2410 -2780
rect 2450 -2850 2520 -2780
rect 2560 -2850 2630 -2780
rect 2670 -2850 2740 -2780
rect 2780 -2850 2850 -2780
rect 2890 -2850 2960 -2780
rect 3000 -2850 3070 -2780
rect 1570 -2960 1640 -2890
rect 1680 -2960 1750 -2890
rect 1790 -2960 1860 -2890
rect 1900 -2960 1970 -2890
rect 2010 -2960 2080 -2890
rect 2120 -2960 2190 -2890
rect 2230 -2960 2300 -2890
rect 2340 -2960 2410 -2890
rect 2450 -2960 2520 -2890
rect 2560 -2960 2630 -2890
rect 2670 -2960 2740 -2890
rect 2780 -2960 2850 -2890
rect 2890 -2960 2960 -2890
rect 3000 -2960 3070 -2890
rect 38190 2900 38260 2970
rect 38280 2900 38350 2970
rect 38370 2900 38440 2970
rect 38190 2810 38260 2880
rect 38280 2810 38350 2880
rect 38370 2810 38440 2880
rect 38190 2720 38260 2790
rect 38280 2720 38350 2790
rect 38370 2720 38440 2790
rect 38190 2630 38260 2700
rect 38280 2630 38350 2700
rect 38370 2630 38440 2700
rect 22470 2530 22540 2600
rect 22580 2530 22650 2600
rect 22690 2530 22760 2600
rect 22800 2530 22870 2600
rect 22470 2420 22540 2490
rect 22580 2420 22650 2490
rect 22690 2420 22760 2490
rect 22800 2420 22870 2490
rect 26950 2530 27020 2600
rect 27060 2530 27130 2600
rect 27170 2530 27240 2600
rect 27280 2530 27350 2600
rect 26950 2420 27020 2490
rect 27060 2420 27130 2490
rect 27170 2420 27240 2490
rect 27280 2420 27350 2490
rect 38190 2540 38260 2610
rect 38280 2540 38350 2610
rect 38370 2540 38440 2610
rect 38190 2450 38260 2520
rect 38280 2450 38350 2520
rect 38370 2450 38440 2520
rect 38190 2360 38260 2430
rect 38280 2360 38350 2430
rect 38370 2360 38440 2430
rect 38190 2270 38260 2340
rect 38280 2270 38350 2340
rect 38370 2270 38440 2340
rect 38190 2180 38260 2250
rect 38280 2180 38350 2250
rect 38370 2180 38440 2250
rect 38190 2090 38260 2160
rect 38280 2090 38350 2160
rect 38370 2090 38440 2160
rect 38190 2000 38260 2070
rect 38280 2000 38350 2070
rect 38370 2000 38440 2070
rect 38190 1910 38260 1980
rect 38280 1910 38350 1980
rect 38370 1910 38440 1980
rect 38190 1820 38260 1890
rect 38280 1820 38350 1890
rect 38370 1820 38440 1890
rect 38190 1730 38260 1800
rect 38280 1730 38350 1800
rect 38370 1730 38440 1800
rect 38190 1640 38260 1710
rect 38280 1640 38350 1710
rect 38370 1640 38440 1710
rect 38190 1550 38260 1620
rect 38280 1550 38350 1620
rect 38370 1550 38440 1620
rect 38190 1460 38260 1530
rect 38280 1460 38350 1530
rect 38370 1460 38440 1530
rect 38190 1370 38260 1440
rect 38280 1370 38350 1440
rect 38370 1370 38440 1440
rect 38190 1280 38260 1350
rect 38280 1280 38350 1350
rect 38370 1280 38440 1350
rect 38190 1190 38260 1260
rect 38280 1190 38350 1260
rect 38370 1190 38440 1260
rect 18995 1090 19065 1160
rect 18995 980 19065 1050
rect 18995 870 19065 940
rect 23490 850 23560 920
rect 23600 850 23670 920
rect 23710 850 23780 920
rect 23820 850 23890 920
rect 23490 740 23560 810
rect 23600 740 23670 810
rect 23710 740 23780 810
rect 23820 740 23890 810
rect 25890 850 25960 920
rect 26000 850 26070 920
rect 26110 850 26180 920
rect 26220 850 26290 920
rect 25890 740 25960 810
rect 26000 740 26070 810
rect 26110 740 26180 810
rect 26220 740 26290 810
rect 38190 150 38260 220
rect 38280 150 38350 220
rect 38370 150 38440 220
rect 38190 60 38260 130
rect 38280 60 38350 130
rect 38370 60 38440 130
rect 30740 -70 30810 0
rect 30850 -70 30920 0
rect 30740 -200 30810 -130
rect 30850 -200 30920 -130
rect 30740 -330 30810 -260
rect 30850 -330 30920 -260
rect 38190 -30 38260 40
rect 38280 -30 38350 40
rect 38370 -30 38440 40
rect 38190 -120 38260 -50
rect 38280 -120 38350 -50
rect 38370 -120 38440 -50
rect 38190 -210 38260 -140
rect 38280 -210 38350 -140
rect 38370 -210 38440 -140
rect 38190 -300 38260 -230
rect 38280 -300 38350 -230
rect 38370 -300 38440 -230
rect 7310 -3950 7380 -3880
rect 7420 -3950 7490 -3880
rect 7530 -3950 7600 -3880
rect 7310 -4060 7380 -3990
rect 7420 -4060 7490 -3990
rect 7530 -4060 7600 -3990
rect 7310 -4170 7380 -4100
rect 7420 -4170 7490 -4100
rect 7530 -4170 7600 -4100
rect -1330 -4420 -1260 -4350
rect -1220 -4420 -1150 -4350
rect -1110 -4420 -1040 -4350
rect -1000 -4420 -930 -4350
rect -1330 -4530 -1260 -4460
rect -1220 -4530 -1150 -4460
rect -1110 -4530 -1040 -4460
rect -1000 -4530 -930 -4460
rect -1160 -6400 -1090 -6330
rect -1070 -6400 -1000 -6330
rect -980 -6400 -910 -6330
rect -890 -6400 -820 -6330
rect -800 -6400 -730 -6330
rect -710 -6400 -640 -6330
rect -620 -6400 -550 -6330
rect -530 -6400 -460 -6330
rect -440 -6400 -370 -6330
rect -350 -6400 -280 -6330
rect -260 -6400 -190 -6330
rect -170 -6400 -100 -6330
rect -80 -6400 -10 -6330
rect 10 -6400 80 -6330
rect -1160 -6490 -1090 -6420
rect -1070 -6490 -1000 -6420
rect -980 -6490 -910 -6420
rect -890 -6490 -820 -6420
rect -800 -6490 -730 -6420
rect -710 -6490 -640 -6420
rect -620 -6490 -550 -6420
rect -530 -6490 -460 -6420
rect -440 -6490 -370 -6420
rect -350 -6490 -280 -6420
rect -260 -6490 -190 -6420
rect -170 -6490 -100 -6420
rect -80 -6490 -10 -6420
rect 10 -6490 80 -6420
rect -1160 -6580 -1090 -6510
rect -1070 -6580 -1000 -6510
rect -980 -6580 -910 -6510
rect -890 -6580 -820 -6510
rect -800 -6580 -730 -6510
rect -710 -6580 -640 -6510
rect -620 -6580 -550 -6510
rect -530 -6580 -460 -6510
rect -440 -6580 -370 -6510
rect -350 -6580 -280 -6510
rect -260 -6580 -190 -6510
rect -170 -6580 -100 -6510
rect -80 -6580 -10 -6510
rect 10 -6580 80 -6510
rect 38190 -390 38260 -320
rect 38280 -390 38350 -320
rect 38370 -390 38440 -320
rect 38190 -520 38260 -450
rect 38280 -520 38350 -450
rect 38370 -520 38440 -450
rect 38190 -610 38260 -540
rect 38280 -610 38350 -540
rect 38370 -610 38440 -540
rect 38190 -700 38260 -630
rect 38280 -700 38350 -630
rect 38370 -700 38440 -630
rect 12250 -860 12320 -790
rect 12360 -860 12430 -790
rect 12470 -860 12540 -790
rect 12580 -860 12650 -790
rect 12690 -860 12760 -790
rect 12800 -860 12870 -790
rect 12910 -860 12980 -790
rect 13020 -860 13090 -790
rect 13130 -860 13200 -790
rect 13240 -860 13310 -790
rect 13350 -860 13420 -790
rect 13460 -860 13530 -790
rect 13570 -860 13640 -790
rect 13680 -860 13750 -790
rect 38190 -790 38260 -720
rect 38280 -790 38350 -720
rect 38370 -790 38440 -720
rect 12250 -970 12320 -900
rect 12360 -970 12430 -900
rect 12470 -970 12540 -900
rect 12580 -970 12650 -900
rect 12690 -970 12760 -900
rect 12800 -970 12870 -900
rect 12910 -970 12980 -900
rect 13020 -970 13090 -900
rect 13130 -970 13200 -900
rect 13240 -970 13310 -900
rect 13350 -970 13420 -900
rect 13460 -970 13530 -900
rect 13570 -970 13640 -900
rect 13680 -970 13750 -900
rect 21820 -920 21890 -850
rect 21930 -920 22000 -850
rect 21820 -1030 21890 -960
rect 21930 -1030 22000 -960
rect 21820 -1140 21890 -1070
rect 21930 -1140 22000 -1070
rect 21820 -1250 21890 -1180
rect 21930 -1250 22000 -1180
rect 21820 -1360 21890 -1290
rect 21930 -1360 22000 -1290
rect 21820 -1470 21890 -1400
rect 21930 -1470 22000 -1400
rect 21820 -1580 21890 -1510
rect 21930 -1580 22000 -1510
rect 21820 -1690 21890 -1620
rect 21930 -1690 22000 -1620
rect 21820 -1800 21890 -1730
rect 21930 -1800 22000 -1730
rect 21820 -1910 21890 -1840
rect 21930 -1910 22000 -1840
rect 21820 -2020 21890 -1950
rect 21930 -2020 22000 -1950
rect 38190 -880 38260 -810
rect 38280 -880 38350 -810
rect 38370 -880 38440 -810
rect 38190 -970 38260 -900
rect 38280 -970 38350 -900
rect 38370 -970 38440 -900
rect 38190 -1060 38260 -990
rect 38280 -1060 38350 -990
rect 38370 -1060 38440 -990
rect 38190 -1150 38260 -1080
rect 38280 -1150 38350 -1080
rect 38370 -1150 38440 -1080
rect 38190 -1240 38260 -1170
rect 38280 -1240 38350 -1170
rect 38370 -1240 38440 -1170
rect 38190 -1330 38260 -1260
rect 38280 -1330 38350 -1260
rect 38370 -1330 38440 -1260
rect 38190 -1420 38260 -1350
rect 38280 -1420 38350 -1350
rect 38370 -1420 38440 -1350
rect 38190 -1510 38260 -1440
rect 38280 -1510 38350 -1440
rect 38370 -1510 38440 -1440
rect 38190 -1600 38260 -1530
rect 38280 -1600 38350 -1530
rect 38370 -1600 38440 -1530
rect 38190 -1690 38260 -1620
rect 38280 -1690 38350 -1620
rect 38370 -1690 38440 -1620
rect 38190 -1780 38260 -1710
rect 38280 -1780 38350 -1710
rect 38370 -1780 38440 -1710
rect 38190 -1870 38260 -1800
rect 38280 -1870 38350 -1800
rect 38370 -1870 38440 -1800
rect 38190 -1960 38260 -1890
rect 38280 -1960 38350 -1890
rect 38370 -1960 38440 -1890
rect 38190 -2050 38260 -1980
rect 38280 -2050 38350 -1980
rect 38370 -2050 38440 -1980
rect 38190 -2140 38260 -2070
rect 38280 -2140 38350 -2070
rect 38370 -2140 38440 -2070
rect 38190 -2230 38260 -2160
rect 38280 -2230 38350 -2160
rect 38370 -2230 38440 -2160
rect 38190 -2320 38260 -2250
rect 38280 -2320 38350 -2250
rect 38370 -2320 38440 -2250
rect 38190 -2410 38260 -2340
rect 38280 -2410 38350 -2340
rect 38370 -2410 38440 -2340
rect 38190 -2500 38260 -2430
rect 38280 -2500 38350 -2430
rect 38370 -2500 38440 -2430
rect 38190 -2590 38260 -2520
rect 38280 -2590 38350 -2520
rect 38370 -2590 38440 -2520
rect 38190 -2680 38260 -2610
rect 38280 -2680 38350 -2610
rect 38370 -2680 38440 -2610
rect 11790 -2850 11860 -2780
rect 11900 -2850 11970 -2780
rect 12010 -2850 12080 -2780
rect 12120 -2850 12190 -2780
rect 12230 -2850 12300 -2780
rect 12340 -2850 12410 -2780
rect 12450 -2850 12520 -2780
rect 12560 -2850 12630 -2780
rect 12670 -2850 12740 -2780
rect 12780 -2850 12850 -2780
rect 12890 -2850 12960 -2780
rect 13000 -2850 13070 -2780
rect 13110 -2850 13180 -2780
rect 13220 -2850 13290 -2780
rect 11790 -2960 11860 -2890
rect 11900 -2960 11970 -2890
rect 12010 -2960 12080 -2890
rect 12120 -2960 12190 -2890
rect 12230 -2960 12300 -2890
rect 12340 -2960 12410 -2890
rect 12450 -2960 12520 -2890
rect 12560 -2960 12630 -2890
rect 12670 -2960 12740 -2890
rect 12780 -2960 12850 -2890
rect 12890 -2960 12960 -2890
rect 13000 -2960 13070 -2890
rect 13110 -2960 13180 -2890
rect 13220 -2960 13290 -2890
rect 38190 -2770 38260 -2700
rect 38280 -2770 38350 -2700
rect 38370 -2770 38440 -2700
rect 38190 -2860 38260 -2790
rect 38280 -2860 38350 -2790
rect 38370 -2860 38440 -2790
rect 38190 -2950 38260 -2880
rect 38280 -2950 38350 -2880
rect 38370 -2950 38440 -2880
rect 24740 -3120 24810 -3050
rect 24850 -3120 24920 -3050
rect 24960 -3120 25030 -3050
rect 24740 -3230 24810 -3160
rect 24850 -3230 24920 -3160
rect 24960 -3230 25030 -3160
rect 24740 -3340 24810 -3270
rect 24850 -3340 24920 -3270
rect 24960 -3340 25030 -3270
rect 38190 -3040 38260 -2970
rect 38280 -3040 38350 -2970
rect 38370 -3040 38440 -2970
rect 38190 -3130 38260 -3060
rect 38280 -3130 38350 -3060
rect 38370 -3130 38440 -3060
rect 38190 -3220 38260 -3150
rect 38280 -3220 38350 -3150
rect 38370 -3220 38440 -3150
rect 38190 -3310 38260 -3240
rect 38280 -3310 38350 -3240
rect 38370 -3310 38440 -3240
rect 38190 -3400 38260 -3330
rect 38280 -3400 38350 -3330
rect 38370 -3400 38440 -3330
rect 38190 -3530 38260 -3460
rect 38280 -3530 38350 -3460
rect 38370 -3530 38440 -3460
rect 38190 -3620 38260 -3550
rect 38280 -3620 38350 -3550
rect 38370 -3620 38440 -3550
rect 22470 -3760 22540 -3690
rect 22580 -3760 22650 -3690
rect 22690 -3760 22760 -3690
rect 22800 -3760 22870 -3690
rect 22470 -3870 22540 -3800
rect 22580 -3870 22650 -3800
rect 22690 -3870 22760 -3800
rect 22800 -3870 22870 -3800
rect 26950 -3760 27020 -3690
rect 27060 -3760 27130 -3690
rect 27170 -3760 27240 -3690
rect 27280 -3760 27350 -3690
rect 26950 -3870 27020 -3800
rect 27060 -3870 27130 -3800
rect 27170 -3870 27240 -3800
rect 27280 -3870 27350 -3800
rect 38190 -3710 38260 -3640
rect 38280 -3710 38350 -3640
rect 38370 -3710 38440 -3640
rect 38190 -3800 38260 -3730
rect 38280 -3800 38350 -3730
rect 38370 -3800 38440 -3730
rect 38190 -3890 38260 -3820
rect 38280 -3890 38350 -3820
rect 38370 -3890 38440 -3820
rect 38190 -3980 38260 -3910
rect 38280 -3980 38350 -3910
rect 38370 -3980 38440 -3910
rect 38190 -4070 38260 -4000
rect 38280 -4070 38350 -4000
rect 38370 -4070 38440 -4000
rect 38190 -4160 38260 -4090
rect 38280 -4160 38350 -4090
rect 38370 -4160 38440 -4090
rect 38190 -4250 38260 -4180
rect 38280 -4250 38350 -4180
rect 38370 -4250 38440 -4180
rect 15710 -4420 15780 -4350
rect 15820 -4420 15890 -4350
rect 15930 -4420 16000 -4350
rect 16040 -4420 16110 -4350
rect 15710 -4530 15780 -4460
rect 15820 -4530 15890 -4460
rect 15930 -4530 16000 -4460
rect 16040 -4530 16110 -4460
rect 38190 -4340 38260 -4270
rect 38280 -4340 38350 -4270
rect 38370 -4340 38440 -4270
rect 38190 -4430 38260 -4360
rect 38280 -4430 38350 -4360
rect 38370 -4430 38440 -4360
rect 38190 -4520 38260 -4450
rect 38280 -4520 38350 -4450
rect 38370 -4520 38440 -4450
rect 38190 -4610 38260 -4540
rect 38280 -4610 38350 -4540
rect 38370 -4610 38440 -4540
rect 14700 -6400 14770 -6330
rect 14790 -6400 14860 -6330
rect 14880 -6400 14950 -6330
rect 14970 -6400 15040 -6330
rect 15060 -6400 15130 -6330
rect 15150 -6400 15220 -6330
rect 15240 -6400 15310 -6330
rect 15330 -6400 15400 -6330
rect 15420 -6400 15490 -6330
rect 15510 -6400 15580 -6330
rect 15600 -6400 15670 -6330
rect 15690 -6400 15760 -6330
rect 15780 -6400 15850 -6330
rect 15870 -6400 15940 -6330
rect 14700 -6490 14770 -6420
rect 14790 -6490 14860 -6420
rect 14880 -6490 14950 -6420
rect 14970 -6490 15040 -6420
rect 15060 -6490 15130 -6420
rect 15150 -6490 15220 -6420
rect 15240 -6490 15310 -6420
rect 15330 -6490 15400 -6420
rect 15420 -6490 15490 -6420
rect 15510 -6490 15580 -6420
rect 15600 -6490 15670 -6420
rect 15690 -6490 15760 -6420
rect 15780 -6490 15850 -6420
rect 15870 -6490 15940 -6420
rect 38190 -4700 38260 -4630
rect 38280 -4700 38350 -4630
rect 38370 -4700 38440 -4630
rect 38190 -4790 38260 -4720
rect 38280 -4790 38350 -4720
rect 38370 -4790 38440 -4720
rect 38190 -4880 38260 -4810
rect 38280 -4880 38350 -4810
rect 38370 -4880 38440 -4810
rect 38190 -4970 38260 -4900
rect 38280 -4970 38350 -4900
rect 38370 -4970 38440 -4900
rect 38190 -5060 38260 -4990
rect 38280 -5060 38350 -4990
rect 38370 -5060 38440 -4990
rect 38190 -5150 38260 -5080
rect 38280 -5150 38350 -5080
rect 38370 -5150 38440 -5080
rect 38190 -5240 38260 -5170
rect 38280 -5240 38350 -5170
rect 38370 -5240 38440 -5170
rect 38190 -5330 38260 -5260
rect 38280 -5330 38350 -5260
rect 38370 -5330 38440 -5260
rect 38190 -5420 38260 -5350
rect 38280 -5420 38350 -5350
rect 38370 -5420 38440 -5350
rect 38190 -5510 38260 -5440
rect 38280 -5510 38350 -5440
rect 38370 -5510 38440 -5440
rect 38190 -5600 38260 -5530
rect 38280 -5600 38350 -5530
rect 38370 -5600 38440 -5530
rect 38190 -5690 38260 -5620
rect 38280 -5690 38350 -5620
rect 38370 -5690 38440 -5620
rect 38190 -5780 38260 -5710
rect 38280 -5780 38350 -5710
rect 38370 -5780 38440 -5710
rect 38190 -5870 38260 -5800
rect 38280 -5870 38350 -5800
rect 38370 -5870 38440 -5800
rect 38190 -5960 38260 -5890
rect 38280 -5960 38350 -5890
rect 38370 -5960 38440 -5890
rect 38190 -6050 38260 -5980
rect 38280 -6050 38350 -5980
rect 38370 -6050 38440 -5980
rect 38190 -6140 38260 -6070
rect 38280 -6140 38350 -6070
rect 38370 -6140 38440 -6070
rect 38190 -6230 38260 -6160
rect 38280 -6230 38350 -6160
rect 38370 -6230 38440 -6160
rect 38190 -6320 38260 -6250
rect 38280 -6320 38350 -6250
rect 38370 -6320 38440 -6250
rect 38190 -6410 38260 -6340
rect 38280 -6410 38350 -6340
rect 38370 -6410 38440 -6340
rect 14700 -6580 14770 -6510
rect 14790 -6580 14860 -6510
rect 14880 -6580 14950 -6510
rect 14970 -6580 15040 -6510
rect 15060 -6580 15130 -6510
rect 15150 -6580 15220 -6510
rect 15240 -6580 15310 -6510
rect 15330 -6580 15400 -6510
rect 15420 -6580 15490 -6510
rect 15510 -6580 15580 -6510
rect 15600 -6580 15670 -6510
rect 15690 -6580 15760 -6510
rect 15780 -6580 15850 -6510
rect 15870 -6580 15940 -6510
rect 20 -8210 90 -8140
rect 130 -8210 200 -8140
rect 230 -8210 300 -8140
rect 20 -8320 90 -8250
rect 130 -8320 200 -8250
rect 230 -8320 300 -8250
rect 20 -8430 90 -8360
rect 130 -8430 200 -8360
rect 230 -8430 300 -8360
rect 1150 -10410 1220 -10340
rect 1260 -10410 1330 -10340
rect 1370 -10410 1440 -10340
rect 1480 -10410 1550 -10340
rect 1590 -10410 1660 -10340
rect 1700 -10410 1770 -10340
rect 1810 -10410 1880 -10340
rect 1920 -10410 1990 -10340
rect 2030 -10410 2100 -10340
rect 2140 -10410 2210 -10340
rect 2250 -10410 2320 -10340
rect 2360 -10410 2430 -10340
rect 2470 -10410 2540 -10340
rect 2580 -10410 2650 -10340
rect 1150 -10520 1220 -10450
rect 1260 -10520 1330 -10450
rect 1370 -10520 1440 -10450
rect 1480 -10520 1550 -10450
rect 1590 -10520 1660 -10450
rect 1700 -10520 1770 -10450
rect 1810 -10520 1880 -10450
rect 1920 -10520 1990 -10450
rect 2030 -10520 2100 -10450
rect 2140 -10520 2210 -10450
rect 2250 -10520 2320 -10450
rect 2360 -10520 2430 -10450
rect 2470 -10520 2540 -10450
rect 2580 -10520 2650 -10450
rect 1540 -12370 1610 -12300
rect 1650 -12370 1720 -12300
rect 1760 -12370 1830 -12300
rect 1870 -12370 1940 -12300
rect 1980 -12370 2050 -12300
rect 2090 -12370 2160 -12300
rect 2200 -12370 2270 -12300
rect 2310 -12370 2380 -12300
rect 2420 -12370 2490 -12300
rect 2530 -12370 2600 -12300
rect 2640 -12370 2710 -12300
rect 2750 -12370 2820 -12300
rect 2860 -12370 2930 -12300
rect 2970 -12370 3040 -12300
rect 1540 -12480 1610 -12410
rect 1650 -12480 1720 -12410
rect 1760 -12480 1830 -12410
rect 1870 -12480 1940 -12410
rect 1980 -12480 2050 -12410
rect 2090 -12480 2160 -12410
rect 2200 -12480 2270 -12410
rect 2310 -12480 2380 -12410
rect 2420 -12480 2490 -12410
rect 2530 -12480 2600 -12410
rect 2640 -12480 2710 -12410
rect 2750 -12480 2820 -12410
rect 2860 -12480 2930 -12410
rect 2970 -12480 3040 -12410
rect 14600 -8300 14670 -8230
rect 14700 -8300 14770 -8230
rect 14810 -8300 14880 -8230
rect 14600 -8410 14670 -8340
rect 14700 -8410 14770 -8340
rect 14810 -8410 14880 -8340
rect 14600 -8520 14670 -8450
rect 14700 -8520 14770 -8450
rect 14810 -8520 14880 -8450
rect 21630 -8430 21700 -8360
rect 21730 -8430 21800 -8360
rect 21830 -8430 21900 -8360
rect 21630 -8530 21700 -8460
rect 21730 -8530 21800 -8460
rect 21830 -8530 21900 -8460
rect 21630 -8630 21700 -8560
rect 21730 -8630 21800 -8560
rect 21830 -8630 21900 -8560
rect 22650 -9080 22720 -9010
rect 22750 -9080 22820 -9010
rect 22850 -9080 22920 -9010
rect 22650 -9180 22720 -9110
rect 22750 -9180 22820 -9110
rect 22850 -9180 22920 -9110
rect 22650 -9280 22720 -9210
rect 22750 -9280 22820 -9210
rect 22850 -9280 22920 -9210
rect 12290 -10440 12360 -10370
rect 12400 -10440 12470 -10370
rect 12510 -10440 12580 -10370
rect 12620 -10440 12690 -10370
rect 12730 -10440 12800 -10370
rect 12840 -10440 12910 -10370
rect 12950 -10440 13020 -10370
rect 13060 -10440 13130 -10370
rect 13170 -10440 13240 -10370
rect 13280 -10440 13350 -10370
rect 13390 -10440 13460 -10370
rect 13500 -10440 13570 -10370
rect 13610 -10440 13680 -10370
rect 13720 -10440 13790 -10370
rect 12290 -10550 12360 -10480
rect 12400 -10550 12470 -10480
rect 12510 -10550 12580 -10480
rect 12620 -10550 12690 -10480
rect 12730 -10550 12800 -10480
rect 12840 -10550 12910 -10480
rect 12950 -10550 13020 -10480
rect 13060 -10550 13130 -10480
rect 13170 -10550 13240 -10480
rect 13280 -10550 13350 -10480
rect 13390 -10550 13460 -10480
rect 13500 -10550 13570 -10480
rect 13610 -10550 13680 -10480
rect 13720 -10550 13790 -10480
rect 29990 -10590 30060 -10520
rect 30700 -10590 30770 -10520
rect 29990 -10700 30060 -10630
rect 30700 -10700 30770 -10630
rect 29990 -10810 30060 -10740
rect 30700 -10810 30770 -10740
rect 11820 -12370 11890 -12300
rect 11930 -12370 12000 -12300
rect 12040 -12370 12110 -12300
rect 12150 -12370 12220 -12300
rect 12260 -12370 12330 -12300
rect 12370 -12370 12440 -12300
rect 12480 -12370 12550 -12300
rect 12590 -12370 12660 -12300
rect 12700 -12370 12770 -12300
rect 12810 -12370 12880 -12300
rect 12920 -12370 12990 -12300
rect 13030 -12370 13100 -12300
rect 13140 -12370 13210 -12300
rect 13250 -12370 13320 -12300
rect 11820 -12480 11890 -12410
rect 11930 -12480 12000 -12410
rect 12040 -12480 12110 -12410
rect 12150 -12480 12220 -12410
rect 12260 -12480 12330 -12410
rect 12370 -12480 12440 -12410
rect 12480 -12480 12550 -12410
rect 12590 -12480 12660 -12410
rect 12700 -12480 12770 -12410
rect 12810 -12480 12880 -12410
rect 12920 -12480 12990 -12410
rect 13030 -12480 13100 -12410
rect 13140 -12480 13210 -12410
rect 13250 -12480 13320 -12410
rect 21630 -14090 21700 -14020
rect 21730 -14090 21800 -14020
rect 21830 -14090 21900 -14020
rect 21630 -14190 21700 -14120
rect 21730 -14190 21800 -14120
rect 21830 -14190 21900 -14120
rect 21630 -14290 21700 -14220
rect 21730 -14290 21800 -14220
rect 21830 -14290 21900 -14220
rect 22920 -14940 22990 -14870
rect 23020 -14940 23090 -14870
rect 23120 -14940 23190 -14870
rect 22920 -15040 22990 -14970
rect 23020 -15040 23090 -14970
rect 23120 -15040 23190 -14970
rect 22920 -15140 22990 -15070
rect 23020 -15140 23090 -15070
rect 23120 -15140 23190 -15070
rect 1620 -22730 1690 -22660
rect 1730 -22730 1800 -22660
rect 1840 -22730 1910 -22660
rect 1950 -22730 2020 -22660
rect 2060 -22730 2130 -22660
rect 2170 -22730 2240 -22660
rect 2280 -22730 2350 -22660
rect 2390 -22730 2460 -22660
rect 2500 -22730 2570 -22660
rect 2610 -22730 2680 -22660
rect 2720 -22730 2790 -22660
rect 2830 -22730 2900 -22660
rect 2940 -22730 3010 -22660
rect 3050 -22730 3120 -22660
rect 1620 -22840 1690 -22770
rect 1730 -22840 1800 -22770
rect 1840 -22840 1910 -22770
rect 1950 -22840 2020 -22770
rect 2060 -22840 2130 -22770
rect 2170 -22840 2240 -22770
rect 2280 -22840 2350 -22770
rect 2390 -22840 2460 -22770
rect 2500 -22840 2570 -22770
rect 2610 -22840 2680 -22770
rect 2720 -22840 2790 -22770
rect 2830 -22840 2900 -22770
rect 2940 -22840 3010 -22770
rect 3050 -22840 3120 -22770
rect 6460 -17820 6530 -17750
rect 6560 -17820 6630 -17750
rect 6660 -17820 6730 -17750
rect 6460 -17930 6530 -17860
rect 6560 -17930 6630 -17860
rect 6660 -17930 6730 -17860
rect 6460 -18040 6530 -17970
rect 6560 -18040 6630 -17970
rect 6660 -18040 6730 -17970
rect 6460 -18150 6530 -18080
rect 6560 -18150 6630 -18080
rect 6660 -18150 6730 -18080
rect 8170 -17820 8240 -17750
rect 8270 -17820 8340 -17750
rect 8370 -17820 8440 -17750
rect 8170 -17930 8240 -17860
rect 8270 -17930 8340 -17860
rect 8370 -17930 8440 -17860
rect 8170 -18040 8240 -17970
rect 8270 -18040 8340 -17970
rect 8370 -18040 8440 -17970
rect 8170 -18150 8240 -18080
rect 8270 -18150 8340 -18080
rect 8370 -18150 8440 -18080
rect 21630 -20170 21700 -20100
rect 21730 -20170 21800 -20100
rect 21830 -20170 21900 -20100
rect 21630 -20270 21700 -20200
rect 21730 -20270 21800 -20200
rect 21830 -20270 21900 -20200
rect 21630 -20370 21700 -20300
rect 21730 -20370 21800 -20300
rect 21830 -20370 21900 -20300
rect 22700 -20800 22770 -20730
rect 22800 -20800 22870 -20730
rect 22900 -20800 22970 -20730
rect 22700 -20900 22770 -20830
rect 22800 -20900 22870 -20830
rect 22900 -20900 22970 -20830
rect 22700 -21000 22770 -20930
rect 22800 -21000 22870 -20930
rect 22900 -21000 22970 -20930
rect 11820 -22730 11890 -22660
rect 11930 -22730 12000 -22660
rect 12040 -22730 12110 -22660
rect 12150 -22730 12220 -22660
rect 12260 -22730 12330 -22660
rect 12370 -22730 12440 -22660
rect 12480 -22730 12550 -22660
rect 12590 -22730 12660 -22660
rect 12700 -22730 12770 -22660
rect 12810 -22730 12880 -22660
rect 12920 -22730 12990 -22660
rect 13030 -22730 13100 -22660
rect 13140 -22730 13210 -22660
rect 13250 -22730 13320 -22660
rect 11820 -22840 11890 -22770
rect 11930 -22840 12000 -22770
rect 12040 -22840 12110 -22770
rect 12150 -22840 12220 -22770
rect 12260 -22840 12330 -22770
rect 12370 -22840 12440 -22770
rect 12480 -22840 12550 -22770
rect 12590 -22840 12660 -22770
rect 12700 -22840 12770 -22770
rect 12810 -22840 12880 -22770
rect 12920 -22840 12990 -22770
rect 13030 -22840 13100 -22770
rect 13140 -22840 13210 -22770
rect 13250 -22840 13320 -22770
<< mimcap >>
rect -5510 20830 6730 20960
rect -5510 20590 -5200 20830
rect -4960 20590 -4870 20830
rect -4630 20590 -4540 20830
rect -4300 20590 -4210 20830
rect -3970 20590 -3880 20830
rect -3640 20590 -3550 20830
rect -3310 20590 -3220 20830
rect -2980 20590 -2890 20830
rect -2650 20590 -2560 20830
rect -2320 20590 -2230 20830
rect -1990 20590 -1900 20830
rect -1660 20590 -1570 20830
rect -1330 20590 -1240 20830
rect -1000 20590 -910 20830
rect -670 20590 -580 20830
rect -340 20590 -250 20830
rect -10 20590 80 20830
rect 320 20590 410 20830
rect 650 20590 740 20830
rect 980 20590 1070 20830
rect 1310 20590 1400 20830
rect 1640 20590 1730 20830
rect 1970 20590 2060 20830
rect 2300 20590 2390 20830
rect 2630 20590 2720 20830
rect 2960 20590 3050 20830
rect 3290 20590 3380 20830
rect 3620 20590 3710 20830
rect 3950 20590 4040 20830
rect 4280 20590 4370 20830
rect 4610 20590 4700 20830
rect 4940 20590 5030 20830
rect 5270 20590 5360 20830
rect 5600 20590 5690 20830
rect 5930 20590 6020 20830
rect 6260 20590 6350 20830
rect 6590 20590 6730 20830
rect -5510 20500 6730 20590
rect -5510 20260 -5200 20500
rect -4960 20260 -4870 20500
rect -4630 20260 -4540 20500
rect -4300 20260 -4210 20500
rect -3970 20260 -3880 20500
rect -3640 20260 -3550 20500
rect -3310 20260 -3220 20500
rect -2980 20260 -2890 20500
rect -2650 20260 -2560 20500
rect -2320 20260 -2230 20500
rect -1990 20260 -1900 20500
rect -1660 20260 -1570 20500
rect -1330 20260 -1240 20500
rect -1000 20260 -910 20500
rect -670 20260 -580 20500
rect -340 20260 -250 20500
rect -10 20260 80 20500
rect 320 20260 410 20500
rect 650 20260 740 20500
rect 980 20260 1070 20500
rect 1310 20260 1400 20500
rect 1640 20260 1730 20500
rect 1970 20260 2060 20500
rect 2300 20260 2390 20500
rect 2630 20260 2720 20500
rect 2960 20260 3050 20500
rect 3290 20260 3380 20500
rect 3620 20260 3710 20500
rect 3950 20260 4040 20500
rect 4280 20260 4370 20500
rect 4610 20260 4700 20500
rect 4940 20260 5030 20500
rect 5270 20260 5360 20500
rect 5600 20260 5690 20500
rect 5930 20260 6020 20500
rect 6260 20260 6350 20500
rect 6590 20260 6730 20500
rect -5510 20170 6730 20260
rect -5510 19930 -5200 20170
rect -4960 19930 -4870 20170
rect -4630 19930 -4540 20170
rect -4300 19930 -4210 20170
rect -3970 19930 -3880 20170
rect -3640 19930 -3550 20170
rect -3310 19930 -3220 20170
rect -2980 19930 -2890 20170
rect -2650 19930 -2560 20170
rect -2320 19930 -2230 20170
rect -1990 19930 -1900 20170
rect -1660 19930 -1570 20170
rect -1330 19930 -1240 20170
rect -1000 19930 -910 20170
rect -670 19930 -580 20170
rect -340 19930 -250 20170
rect -10 19930 80 20170
rect 320 19930 410 20170
rect 650 19930 740 20170
rect 980 19930 1070 20170
rect 1310 19930 1400 20170
rect 1640 19930 1730 20170
rect 1970 19930 2060 20170
rect 2300 19930 2390 20170
rect 2630 19930 2720 20170
rect 2960 19930 3050 20170
rect 3290 19930 3380 20170
rect 3620 19930 3710 20170
rect 3950 19930 4040 20170
rect 4280 19930 4370 20170
rect 4610 19930 4700 20170
rect 4940 19930 5030 20170
rect 5270 19930 5360 20170
rect 5600 19930 5690 20170
rect 5930 19930 6020 20170
rect 6260 19930 6350 20170
rect 6590 19930 6730 20170
rect -5510 19840 6730 19930
rect -5510 19600 -5200 19840
rect -4960 19600 -4870 19840
rect -4630 19600 -4540 19840
rect -4300 19600 -4210 19840
rect -3970 19600 -3880 19840
rect -3640 19600 -3550 19840
rect -3310 19600 -3220 19840
rect -2980 19600 -2890 19840
rect -2650 19600 -2560 19840
rect -2320 19600 -2230 19840
rect -1990 19600 -1900 19840
rect -1660 19600 -1570 19840
rect -1330 19600 -1240 19840
rect -1000 19600 -910 19840
rect -670 19600 -580 19840
rect -340 19600 -250 19840
rect -10 19600 80 19840
rect 320 19600 410 19840
rect 650 19600 740 19840
rect 980 19600 1070 19840
rect 1310 19600 1400 19840
rect 1640 19600 1730 19840
rect 1970 19600 2060 19840
rect 2300 19600 2390 19840
rect 2630 19600 2720 19840
rect 2960 19600 3050 19840
rect 3290 19600 3380 19840
rect 3620 19600 3710 19840
rect 3950 19600 4040 19840
rect 4280 19600 4370 19840
rect 4610 19600 4700 19840
rect 4940 19600 5030 19840
rect 5270 19600 5360 19840
rect 5600 19600 5690 19840
rect 5930 19600 6020 19840
rect 6260 19600 6350 19840
rect 6590 19600 6730 19840
rect -5510 19510 6730 19600
rect -5510 19270 -5200 19510
rect -4960 19270 -4870 19510
rect -4630 19270 -4540 19510
rect -4300 19270 -4210 19510
rect -3970 19270 -3880 19510
rect -3640 19270 -3550 19510
rect -3310 19270 -3220 19510
rect -2980 19270 -2890 19510
rect -2650 19270 -2560 19510
rect -2320 19270 -2230 19510
rect -1990 19270 -1900 19510
rect -1660 19270 -1570 19510
rect -1330 19270 -1240 19510
rect -1000 19270 -910 19510
rect -670 19270 -580 19510
rect -340 19270 -250 19510
rect -10 19270 80 19510
rect 320 19270 410 19510
rect 650 19270 740 19510
rect 980 19270 1070 19510
rect 1310 19270 1400 19510
rect 1640 19270 1730 19510
rect 1970 19270 2060 19510
rect 2300 19270 2390 19510
rect 2630 19270 2720 19510
rect 2960 19270 3050 19510
rect 3290 19270 3380 19510
rect 3620 19270 3710 19510
rect 3950 19270 4040 19510
rect 4280 19270 4370 19510
rect 4610 19270 4700 19510
rect 4940 19270 5030 19510
rect 5270 19270 5360 19510
rect 5600 19270 5690 19510
rect 5930 19270 6020 19510
rect 6260 19270 6350 19510
rect 6590 19270 6730 19510
rect -5510 19180 6730 19270
rect -5510 18940 -5200 19180
rect -4960 18940 -4870 19180
rect -4630 18940 -4540 19180
rect -4300 18940 -4210 19180
rect -3970 18940 -3880 19180
rect -3640 18940 -3550 19180
rect -3310 18940 -3220 19180
rect -2980 18940 -2890 19180
rect -2650 18940 -2560 19180
rect -2320 18940 -2230 19180
rect -1990 18940 -1900 19180
rect -1660 18940 -1570 19180
rect -1330 18940 -1240 19180
rect -1000 18940 -910 19180
rect -670 18940 -580 19180
rect -340 18940 -250 19180
rect -10 18940 80 19180
rect 320 18940 410 19180
rect 650 18940 740 19180
rect 980 18940 1070 19180
rect 1310 18940 1400 19180
rect 1640 18940 1730 19180
rect 1970 18940 2060 19180
rect 2300 18940 2390 19180
rect 2630 18940 2720 19180
rect 2960 18940 3050 19180
rect 3290 18940 3380 19180
rect 3620 18940 3710 19180
rect 3950 18940 4040 19180
rect 4280 18940 4370 19180
rect 4610 18940 4700 19180
rect 4940 18940 5030 19180
rect 5270 18940 5360 19180
rect 5600 18940 5690 19180
rect 5930 18940 6020 19180
rect 6260 18940 6350 19180
rect 6590 18940 6730 19180
rect -5510 18850 6730 18940
rect -5510 18610 -5200 18850
rect -4960 18610 -4870 18850
rect -4630 18610 -4540 18850
rect -4300 18610 -4210 18850
rect -3970 18610 -3880 18850
rect -3640 18610 -3550 18850
rect -3310 18610 -3220 18850
rect -2980 18610 -2890 18850
rect -2650 18610 -2560 18850
rect -2320 18610 -2230 18850
rect -1990 18610 -1900 18850
rect -1660 18610 -1570 18850
rect -1330 18610 -1240 18850
rect -1000 18610 -910 18850
rect -670 18610 -580 18850
rect -340 18610 -250 18850
rect -10 18610 80 18850
rect 320 18610 410 18850
rect 650 18610 740 18850
rect 980 18610 1070 18850
rect 1310 18610 1400 18850
rect 1640 18610 1730 18850
rect 1970 18610 2060 18850
rect 2300 18610 2390 18850
rect 2630 18610 2720 18850
rect 2960 18610 3050 18850
rect 3290 18610 3380 18850
rect 3620 18610 3710 18850
rect 3950 18610 4040 18850
rect 4280 18610 4370 18850
rect 4610 18610 4700 18850
rect 4940 18610 5030 18850
rect 5270 18610 5360 18850
rect 5600 18610 5690 18850
rect 5930 18610 6020 18850
rect 6260 18610 6350 18850
rect 6590 18610 6730 18850
rect -5510 18520 6730 18610
rect -5510 18280 -5200 18520
rect -4960 18280 -4870 18520
rect -4630 18280 -4540 18520
rect -4300 18280 -4210 18520
rect -3970 18280 -3880 18520
rect -3640 18280 -3550 18520
rect -3310 18280 -3220 18520
rect -2980 18280 -2890 18520
rect -2650 18280 -2560 18520
rect -2320 18280 -2230 18520
rect -1990 18280 -1900 18520
rect -1660 18280 -1570 18520
rect -1330 18280 -1240 18520
rect -1000 18280 -910 18520
rect -670 18280 -580 18520
rect -340 18280 -250 18520
rect -10 18280 80 18520
rect 320 18280 410 18520
rect 650 18280 740 18520
rect 980 18280 1070 18520
rect 1310 18280 1400 18520
rect 1640 18280 1730 18520
rect 1970 18280 2060 18520
rect 2300 18280 2390 18520
rect 2630 18280 2720 18520
rect 2960 18280 3050 18520
rect 3290 18280 3380 18520
rect 3620 18280 3710 18520
rect 3950 18280 4040 18520
rect 4280 18280 4370 18520
rect 4610 18280 4700 18520
rect 4940 18280 5030 18520
rect 5270 18280 5360 18520
rect 5600 18280 5690 18520
rect 5930 18280 6020 18520
rect 6260 18280 6350 18520
rect 6590 18280 6730 18520
rect -5510 18190 6730 18280
rect -5510 17950 -5200 18190
rect -4960 17950 -4870 18190
rect -4630 17950 -4540 18190
rect -4300 17950 -4210 18190
rect -3970 17950 -3880 18190
rect -3640 17950 -3550 18190
rect -3310 17950 -3220 18190
rect -2980 17950 -2890 18190
rect -2650 17950 -2560 18190
rect -2320 17950 -2230 18190
rect -1990 17950 -1900 18190
rect -1660 17950 -1570 18190
rect -1330 17950 -1240 18190
rect -1000 17950 -910 18190
rect -670 17950 -580 18190
rect -340 17950 -250 18190
rect -10 17950 80 18190
rect 320 17950 410 18190
rect 650 17950 740 18190
rect 980 17950 1070 18190
rect 1310 17950 1400 18190
rect 1640 17950 1730 18190
rect 1970 17950 2060 18190
rect 2300 17950 2390 18190
rect 2630 17950 2720 18190
rect 2960 17950 3050 18190
rect 3290 17950 3380 18190
rect 3620 17950 3710 18190
rect 3950 17950 4040 18190
rect 4280 17950 4370 18190
rect 4610 17950 4700 18190
rect 4940 17950 5030 18190
rect 5270 17950 5360 18190
rect 5600 17950 5690 18190
rect 5930 17950 6020 18190
rect 6260 17950 6350 18190
rect 6590 17950 6730 18190
rect -5510 17860 6730 17950
rect -5510 17620 -5200 17860
rect -4960 17620 -4870 17860
rect -4630 17620 -4540 17860
rect -4300 17620 -4210 17860
rect -3970 17620 -3880 17860
rect -3640 17620 -3550 17860
rect -3310 17620 -3220 17860
rect -2980 17620 -2890 17860
rect -2650 17620 -2560 17860
rect -2320 17620 -2230 17860
rect -1990 17620 -1900 17860
rect -1660 17620 -1570 17860
rect -1330 17620 -1240 17860
rect -1000 17620 -910 17860
rect -670 17620 -580 17860
rect -340 17620 -250 17860
rect -10 17620 80 17860
rect 320 17620 410 17860
rect 650 17620 740 17860
rect 980 17620 1070 17860
rect 1310 17620 1400 17860
rect 1640 17620 1730 17860
rect 1970 17620 2060 17860
rect 2300 17620 2390 17860
rect 2630 17620 2720 17860
rect 2960 17620 3050 17860
rect 3290 17620 3380 17860
rect 3620 17620 3710 17860
rect 3950 17620 4040 17860
rect 4280 17620 4370 17860
rect 4610 17620 4700 17860
rect 4940 17620 5030 17860
rect 5270 17620 5360 17860
rect 5600 17620 5690 17860
rect 5930 17620 6020 17860
rect 6260 17620 6350 17860
rect 6590 17620 6730 17860
rect -5510 17530 6730 17620
rect -5510 17290 -5200 17530
rect -4960 17290 -4870 17530
rect -4630 17290 -4540 17530
rect -4300 17290 -4210 17530
rect -3970 17290 -3880 17530
rect -3640 17290 -3550 17530
rect -3310 17290 -3220 17530
rect -2980 17290 -2890 17530
rect -2650 17290 -2560 17530
rect -2320 17290 -2230 17530
rect -1990 17290 -1900 17530
rect -1660 17290 -1570 17530
rect -1330 17290 -1240 17530
rect -1000 17290 -910 17530
rect -670 17290 -580 17530
rect -340 17290 -250 17530
rect -10 17290 80 17530
rect 320 17290 410 17530
rect 650 17290 740 17530
rect 980 17290 1070 17530
rect 1310 17290 1400 17530
rect 1640 17290 1730 17530
rect 1970 17290 2060 17530
rect 2300 17290 2390 17530
rect 2630 17290 2720 17530
rect 2960 17290 3050 17530
rect 3290 17290 3380 17530
rect 3620 17290 3710 17530
rect 3950 17290 4040 17530
rect 4280 17290 4370 17530
rect 4610 17290 4700 17530
rect 4940 17290 5030 17530
rect 5270 17290 5360 17530
rect 5600 17290 5690 17530
rect 5930 17290 6020 17530
rect 6260 17290 6350 17530
rect 6590 17290 6730 17530
rect -5510 17200 6730 17290
rect -5510 16960 -5200 17200
rect -4960 16960 -4870 17200
rect -4630 16960 -4540 17200
rect -4300 16960 -4210 17200
rect -3970 16960 -3880 17200
rect -3640 16960 -3550 17200
rect -3310 16960 -3220 17200
rect -2980 16960 -2890 17200
rect -2650 16960 -2560 17200
rect -2320 16960 -2230 17200
rect -1990 16960 -1900 17200
rect -1660 16960 -1570 17200
rect -1330 16960 -1240 17200
rect -1000 16960 -910 17200
rect -670 16960 -580 17200
rect -340 16960 -250 17200
rect -10 16960 80 17200
rect 320 16960 410 17200
rect 650 16960 740 17200
rect 980 16960 1070 17200
rect 1310 16960 1400 17200
rect 1640 16960 1730 17200
rect 1970 16960 2060 17200
rect 2300 16960 2390 17200
rect 2630 16960 2720 17200
rect 2960 16960 3050 17200
rect 3290 16960 3380 17200
rect 3620 16960 3710 17200
rect 3950 16960 4040 17200
rect 4280 16960 4370 17200
rect 4610 16960 4700 17200
rect 4940 16960 5030 17200
rect 5270 16960 5360 17200
rect 5600 16960 5690 17200
rect 5930 16960 6020 17200
rect 6260 16960 6350 17200
rect 6590 16960 6730 17200
rect -5510 16870 6730 16960
rect -5510 16630 -5200 16870
rect -4960 16630 -4870 16870
rect -4630 16630 -4540 16870
rect -4300 16630 -4210 16870
rect -3970 16630 -3880 16870
rect -3640 16630 -3550 16870
rect -3310 16630 -3220 16870
rect -2980 16630 -2890 16870
rect -2650 16630 -2560 16870
rect -2320 16630 -2230 16870
rect -1990 16630 -1900 16870
rect -1660 16630 -1570 16870
rect -1330 16630 -1240 16870
rect -1000 16630 -910 16870
rect -670 16630 -580 16870
rect -340 16630 -250 16870
rect -10 16630 80 16870
rect 320 16630 410 16870
rect 650 16630 740 16870
rect 980 16630 1070 16870
rect 1310 16630 1400 16870
rect 1640 16630 1730 16870
rect 1970 16630 2060 16870
rect 2300 16630 2390 16870
rect 2630 16630 2720 16870
rect 2960 16630 3050 16870
rect 3290 16630 3380 16870
rect 3620 16630 3710 16870
rect 3950 16630 4040 16870
rect 4280 16630 4370 16870
rect 4610 16630 4700 16870
rect 4940 16630 5030 16870
rect 5270 16630 5360 16870
rect 5600 16630 5690 16870
rect 5930 16630 6020 16870
rect 6260 16630 6350 16870
rect 6590 16630 6730 16870
rect -5510 16540 6730 16630
rect -5510 16300 -5200 16540
rect -4960 16300 -4870 16540
rect -4630 16300 -4540 16540
rect -4300 16300 -4210 16540
rect -3970 16300 -3880 16540
rect -3640 16300 -3550 16540
rect -3310 16300 -3220 16540
rect -2980 16300 -2890 16540
rect -2650 16300 -2560 16540
rect -2320 16300 -2230 16540
rect -1990 16300 -1900 16540
rect -1660 16300 -1570 16540
rect -1330 16300 -1240 16540
rect -1000 16300 -910 16540
rect -670 16300 -580 16540
rect -340 16300 -250 16540
rect -10 16300 80 16540
rect 320 16300 410 16540
rect 650 16300 740 16540
rect 980 16300 1070 16540
rect 1310 16300 1400 16540
rect 1640 16300 1730 16540
rect 1970 16300 2060 16540
rect 2300 16300 2390 16540
rect 2630 16300 2720 16540
rect 2960 16300 3050 16540
rect 3290 16300 3380 16540
rect 3620 16300 3710 16540
rect 3950 16300 4040 16540
rect 4280 16300 4370 16540
rect 4610 16300 4700 16540
rect 4940 16300 5030 16540
rect 5270 16300 5360 16540
rect 5600 16300 5690 16540
rect 5930 16300 6020 16540
rect 6260 16300 6350 16540
rect 6590 16300 6730 16540
rect -5510 16210 6730 16300
rect -5510 15970 -5200 16210
rect -4960 15970 -4870 16210
rect -4630 15970 -4540 16210
rect -4300 15970 -4210 16210
rect -3970 15970 -3880 16210
rect -3640 15970 -3550 16210
rect -3310 15970 -3220 16210
rect -2980 15970 -2890 16210
rect -2650 15970 -2560 16210
rect -2320 15970 -2230 16210
rect -1990 15970 -1900 16210
rect -1660 15970 -1570 16210
rect -1330 15970 -1240 16210
rect -1000 15970 -910 16210
rect -670 15970 -580 16210
rect -340 15970 -250 16210
rect -10 15970 80 16210
rect 320 15970 410 16210
rect 650 15970 740 16210
rect 980 15970 1070 16210
rect 1310 15970 1400 16210
rect 1640 15970 1730 16210
rect 1970 15970 2060 16210
rect 2300 15970 2390 16210
rect 2630 15970 2720 16210
rect 2960 15970 3050 16210
rect 3290 15970 3380 16210
rect 3620 15970 3710 16210
rect 3950 15970 4040 16210
rect 4280 15970 4370 16210
rect 4610 15970 4700 16210
rect 4940 15970 5030 16210
rect 5270 15970 5360 16210
rect 5600 15970 5690 16210
rect 5930 15970 6020 16210
rect 6260 15970 6350 16210
rect 6590 15970 6730 16210
rect -5510 15880 6730 15970
rect -5510 15640 -5200 15880
rect -4960 15640 -4870 15880
rect -4630 15640 -4540 15880
rect -4300 15640 -4210 15880
rect -3970 15640 -3880 15880
rect -3640 15640 -3550 15880
rect -3310 15640 -3220 15880
rect -2980 15640 -2890 15880
rect -2650 15640 -2560 15880
rect -2320 15640 -2230 15880
rect -1990 15640 -1900 15880
rect -1660 15640 -1570 15880
rect -1330 15640 -1240 15880
rect -1000 15640 -910 15880
rect -670 15640 -580 15880
rect -340 15640 -250 15880
rect -10 15640 80 15880
rect 320 15640 410 15880
rect 650 15640 740 15880
rect 980 15640 1070 15880
rect 1310 15640 1400 15880
rect 1640 15640 1730 15880
rect 1970 15640 2060 15880
rect 2300 15640 2390 15880
rect 2630 15640 2720 15880
rect 2960 15640 3050 15880
rect 3290 15640 3380 15880
rect 3620 15640 3710 15880
rect 3950 15640 4040 15880
rect 4280 15640 4370 15880
rect 4610 15640 4700 15880
rect 4940 15640 5030 15880
rect 5270 15640 5360 15880
rect 5600 15640 5690 15880
rect 5930 15640 6020 15880
rect 6260 15640 6350 15880
rect 6590 15640 6730 15880
rect -5510 15550 6730 15640
rect -5510 15310 -5200 15550
rect -4960 15310 -4870 15550
rect -4630 15310 -4540 15550
rect -4300 15310 -4210 15550
rect -3970 15310 -3880 15550
rect -3640 15310 -3550 15550
rect -3310 15310 -3220 15550
rect -2980 15310 -2890 15550
rect -2650 15310 -2560 15550
rect -2320 15310 -2230 15550
rect -1990 15310 -1900 15550
rect -1660 15310 -1570 15550
rect -1330 15310 -1240 15550
rect -1000 15310 -910 15550
rect -670 15310 -580 15550
rect -340 15310 -250 15550
rect -10 15310 80 15550
rect 320 15310 410 15550
rect 650 15310 740 15550
rect 980 15310 1070 15550
rect 1310 15310 1400 15550
rect 1640 15310 1730 15550
rect 1970 15310 2060 15550
rect 2300 15310 2390 15550
rect 2630 15310 2720 15550
rect 2960 15310 3050 15550
rect 3290 15310 3380 15550
rect 3620 15310 3710 15550
rect 3950 15310 4040 15550
rect 4280 15310 4370 15550
rect 4610 15310 4700 15550
rect 4940 15310 5030 15550
rect 5270 15310 5360 15550
rect 5600 15310 5690 15550
rect 5930 15310 6020 15550
rect 6260 15310 6350 15550
rect 6590 15310 6730 15550
rect -5510 15220 6730 15310
rect -5510 14980 -5200 15220
rect -4960 14980 -4870 15220
rect -4630 14980 -4540 15220
rect -4300 14980 -4210 15220
rect -3970 14980 -3880 15220
rect -3640 14980 -3550 15220
rect -3310 14980 -3220 15220
rect -2980 14980 -2890 15220
rect -2650 14980 -2560 15220
rect -2320 14980 -2230 15220
rect -1990 14980 -1900 15220
rect -1660 14980 -1570 15220
rect -1330 14980 -1240 15220
rect -1000 14980 -910 15220
rect -670 14980 -580 15220
rect -340 14980 -250 15220
rect -10 14980 80 15220
rect 320 14980 410 15220
rect 650 14980 740 15220
rect 980 14980 1070 15220
rect 1310 14980 1400 15220
rect 1640 14980 1730 15220
rect 1970 14980 2060 15220
rect 2300 14980 2390 15220
rect 2630 14980 2720 15220
rect 2960 14980 3050 15220
rect 3290 14980 3380 15220
rect 3620 14980 3710 15220
rect 3950 14980 4040 15220
rect 4280 14980 4370 15220
rect 4610 14980 4700 15220
rect 4940 14980 5030 15220
rect 5270 14980 5360 15220
rect 5600 14980 5690 15220
rect 5930 14980 6020 15220
rect 6260 14980 6350 15220
rect 6590 14980 6730 15220
rect -5510 14890 6730 14980
rect -5510 14650 -5200 14890
rect -4960 14650 -4870 14890
rect -4630 14650 -4540 14890
rect -4300 14650 -4210 14890
rect -3970 14650 -3880 14890
rect -3640 14650 -3550 14890
rect -3310 14650 -3220 14890
rect -2980 14650 -2890 14890
rect -2650 14650 -2560 14890
rect -2320 14650 -2230 14890
rect -1990 14650 -1900 14890
rect -1660 14650 -1570 14890
rect -1330 14650 -1240 14890
rect -1000 14650 -910 14890
rect -670 14650 -580 14890
rect -340 14650 -250 14890
rect -10 14650 80 14890
rect 320 14650 410 14890
rect 650 14650 740 14890
rect 980 14650 1070 14890
rect 1310 14650 1400 14890
rect 1640 14650 1730 14890
rect 1970 14650 2060 14890
rect 2300 14650 2390 14890
rect 2630 14650 2720 14890
rect 2960 14650 3050 14890
rect 3290 14650 3380 14890
rect 3620 14650 3710 14890
rect 3950 14650 4040 14890
rect 4280 14650 4370 14890
rect 4610 14650 4700 14890
rect 4940 14650 5030 14890
rect 5270 14650 5360 14890
rect 5600 14650 5690 14890
rect 5930 14650 6020 14890
rect 6260 14650 6350 14890
rect 6590 14650 6730 14890
rect -5510 14560 6730 14650
rect -5510 14320 -5200 14560
rect -4960 14320 -4870 14560
rect -4630 14320 -4540 14560
rect -4300 14320 -4210 14560
rect -3970 14320 -3880 14560
rect -3640 14320 -3550 14560
rect -3310 14320 -3220 14560
rect -2980 14320 -2890 14560
rect -2650 14320 -2560 14560
rect -2320 14320 -2230 14560
rect -1990 14320 -1900 14560
rect -1660 14320 -1570 14560
rect -1330 14320 -1240 14560
rect -1000 14320 -910 14560
rect -670 14320 -580 14560
rect -340 14320 -250 14560
rect -10 14320 80 14560
rect 320 14320 410 14560
rect 650 14320 740 14560
rect 980 14320 1070 14560
rect 1310 14320 1400 14560
rect 1640 14320 1730 14560
rect 1970 14320 2060 14560
rect 2300 14320 2390 14560
rect 2630 14320 2720 14560
rect 2960 14320 3050 14560
rect 3290 14320 3380 14560
rect 3620 14320 3710 14560
rect 3950 14320 4040 14560
rect 4280 14320 4370 14560
rect 4610 14320 4700 14560
rect 4940 14320 5030 14560
rect 5270 14320 5360 14560
rect 5600 14320 5690 14560
rect 5930 14320 6020 14560
rect 6260 14320 6350 14560
rect 6590 14320 6730 14560
rect -5510 14230 6730 14320
rect -5510 13990 -5200 14230
rect -4960 13990 -4870 14230
rect -4630 13990 -4540 14230
rect -4300 13990 -4210 14230
rect -3970 13990 -3880 14230
rect -3640 13990 -3550 14230
rect -3310 13990 -3220 14230
rect -2980 13990 -2890 14230
rect -2650 13990 -2560 14230
rect -2320 13990 -2230 14230
rect -1990 13990 -1900 14230
rect -1660 13990 -1570 14230
rect -1330 13990 -1240 14230
rect -1000 13990 -910 14230
rect -670 13990 -580 14230
rect -340 13990 -250 14230
rect -10 13990 80 14230
rect 320 13990 410 14230
rect 650 13990 740 14230
rect 980 13990 1070 14230
rect 1310 13990 1400 14230
rect 1640 13990 1730 14230
rect 1970 13990 2060 14230
rect 2300 13990 2390 14230
rect 2630 13990 2720 14230
rect 2960 13990 3050 14230
rect 3290 13990 3380 14230
rect 3620 13990 3710 14230
rect 3950 13990 4040 14230
rect 4280 13990 4370 14230
rect 4610 13990 4700 14230
rect 4940 13990 5030 14230
rect 5270 13990 5360 14230
rect 5600 13990 5690 14230
rect 5930 13990 6020 14230
rect 6260 13990 6350 14230
rect 6590 13990 6730 14230
rect -5510 13900 6730 13990
rect -5510 13660 -5200 13900
rect -4960 13660 -4870 13900
rect -4630 13660 -4540 13900
rect -4300 13660 -4210 13900
rect -3970 13660 -3880 13900
rect -3640 13660 -3550 13900
rect -3310 13660 -3220 13900
rect -2980 13660 -2890 13900
rect -2650 13660 -2560 13900
rect -2320 13660 -2230 13900
rect -1990 13660 -1900 13900
rect -1660 13660 -1570 13900
rect -1330 13660 -1240 13900
rect -1000 13660 -910 13900
rect -670 13660 -580 13900
rect -340 13660 -250 13900
rect -10 13660 80 13900
rect 320 13660 410 13900
rect 650 13660 740 13900
rect 980 13660 1070 13900
rect 1310 13660 1400 13900
rect 1640 13660 1730 13900
rect 1970 13660 2060 13900
rect 2300 13660 2390 13900
rect 2630 13660 2720 13900
rect 2960 13660 3050 13900
rect 3290 13660 3380 13900
rect 3620 13660 3710 13900
rect 3950 13660 4040 13900
rect 4280 13660 4370 13900
rect 4610 13660 4700 13900
rect 4940 13660 5030 13900
rect 5270 13660 5360 13900
rect 5600 13660 5690 13900
rect 5930 13660 6020 13900
rect 6260 13660 6350 13900
rect 6590 13660 6730 13900
rect -5510 13570 6730 13660
rect -5510 13330 -5200 13570
rect -4960 13330 -4870 13570
rect -4630 13330 -4540 13570
rect -4300 13330 -4210 13570
rect -3970 13330 -3880 13570
rect -3640 13330 -3550 13570
rect -3310 13330 -3220 13570
rect -2980 13330 -2890 13570
rect -2650 13330 -2560 13570
rect -2320 13330 -2230 13570
rect -1990 13330 -1900 13570
rect -1660 13330 -1570 13570
rect -1330 13330 -1240 13570
rect -1000 13330 -910 13570
rect -670 13330 -580 13570
rect -340 13330 -250 13570
rect -10 13330 80 13570
rect 320 13330 410 13570
rect 650 13330 740 13570
rect 980 13330 1070 13570
rect 1310 13330 1400 13570
rect 1640 13330 1730 13570
rect 1970 13330 2060 13570
rect 2300 13330 2390 13570
rect 2630 13330 2720 13570
rect 2960 13330 3050 13570
rect 3290 13330 3380 13570
rect 3620 13330 3710 13570
rect 3950 13330 4040 13570
rect 4280 13330 4370 13570
rect 4610 13330 4700 13570
rect 4940 13330 5030 13570
rect 5270 13330 5360 13570
rect 5600 13330 5690 13570
rect 5930 13330 6020 13570
rect 6260 13330 6350 13570
rect 6590 13330 6730 13570
rect -5510 13240 6730 13330
rect -5510 13000 -5200 13240
rect -4960 13000 -4870 13240
rect -4630 13000 -4540 13240
rect -4300 13000 -4210 13240
rect -3970 13000 -3880 13240
rect -3640 13000 -3550 13240
rect -3310 13000 -3220 13240
rect -2980 13000 -2890 13240
rect -2650 13000 -2560 13240
rect -2320 13000 -2230 13240
rect -1990 13000 -1900 13240
rect -1660 13000 -1570 13240
rect -1330 13000 -1240 13240
rect -1000 13000 -910 13240
rect -670 13000 -580 13240
rect -340 13000 -250 13240
rect -10 13000 80 13240
rect 320 13000 410 13240
rect 650 13000 740 13240
rect 980 13000 1070 13240
rect 1310 13000 1400 13240
rect 1640 13000 1730 13240
rect 1970 13000 2060 13240
rect 2300 13000 2390 13240
rect 2630 13000 2720 13240
rect 2960 13000 3050 13240
rect 3290 13000 3380 13240
rect 3620 13000 3710 13240
rect 3950 13000 4040 13240
rect 4280 13000 4370 13240
rect 4610 13000 4700 13240
rect 4940 13000 5030 13240
rect 5270 13000 5360 13240
rect 5600 13000 5690 13240
rect 5930 13000 6020 13240
rect 6260 13000 6350 13240
rect 6590 13000 6730 13240
rect -5510 12910 6730 13000
rect -5510 12670 -5200 12910
rect -4960 12670 -4870 12910
rect -4630 12670 -4540 12910
rect -4300 12670 -4210 12910
rect -3970 12670 -3880 12910
rect -3640 12670 -3550 12910
rect -3310 12670 -3220 12910
rect -2980 12670 -2890 12910
rect -2650 12670 -2560 12910
rect -2320 12670 -2230 12910
rect -1990 12670 -1900 12910
rect -1660 12670 -1570 12910
rect -1330 12670 -1240 12910
rect -1000 12670 -910 12910
rect -670 12670 -580 12910
rect -340 12670 -250 12910
rect -10 12670 80 12910
rect 320 12670 410 12910
rect 650 12670 740 12910
rect 980 12670 1070 12910
rect 1310 12670 1400 12910
rect 1640 12670 1730 12910
rect 1970 12670 2060 12910
rect 2300 12670 2390 12910
rect 2630 12670 2720 12910
rect 2960 12670 3050 12910
rect 3290 12670 3380 12910
rect 3620 12670 3710 12910
rect 3950 12670 4040 12910
rect 4280 12670 4370 12910
rect 4610 12670 4700 12910
rect 4940 12670 5030 12910
rect 5270 12670 5360 12910
rect 5600 12670 5690 12910
rect 5930 12670 6020 12910
rect 6260 12670 6350 12910
rect 6590 12670 6730 12910
rect -5510 12580 6730 12670
rect -5510 12340 -5200 12580
rect -4960 12340 -4870 12580
rect -4630 12340 -4540 12580
rect -4300 12340 -4210 12580
rect -3970 12340 -3880 12580
rect -3640 12340 -3550 12580
rect -3310 12340 -3220 12580
rect -2980 12340 -2890 12580
rect -2650 12340 -2560 12580
rect -2320 12340 -2230 12580
rect -1990 12340 -1900 12580
rect -1660 12340 -1570 12580
rect -1330 12340 -1240 12580
rect -1000 12340 -910 12580
rect -670 12340 -580 12580
rect -340 12340 -250 12580
rect -10 12340 80 12580
rect 320 12340 410 12580
rect 650 12340 740 12580
rect 980 12340 1070 12580
rect 1310 12340 1400 12580
rect 1640 12340 1730 12580
rect 1970 12340 2060 12580
rect 2300 12340 2390 12580
rect 2630 12340 2720 12580
rect 2960 12340 3050 12580
rect 3290 12340 3380 12580
rect 3620 12340 3710 12580
rect 3950 12340 4040 12580
rect 4280 12340 4370 12580
rect 4610 12340 4700 12580
rect 4940 12340 5030 12580
rect 5270 12340 5360 12580
rect 5600 12340 5690 12580
rect 5930 12340 6020 12580
rect 6260 12340 6350 12580
rect 6590 12340 6730 12580
rect -5510 12250 6730 12340
rect -5510 12010 -5200 12250
rect -4960 12010 -4870 12250
rect -4630 12010 -4540 12250
rect -4300 12010 -4210 12250
rect -3970 12010 -3880 12250
rect -3640 12010 -3550 12250
rect -3310 12010 -3220 12250
rect -2980 12010 -2890 12250
rect -2650 12010 -2560 12250
rect -2320 12010 -2230 12250
rect -1990 12010 -1900 12250
rect -1660 12010 -1570 12250
rect -1330 12010 -1240 12250
rect -1000 12010 -910 12250
rect -670 12010 -580 12250
rect -340 12010 -250 12250
rect -10 12010 80 12250
rect 320 12010 410 12250
rect 650 12010 740 12250
rect 980 12010 1070 12250
rect 1310 12010 1400 12250
rect 1640 12010 1730 12250
rect 1970 12010 2060 12250
rect 2300 12010 2390 12250
rect 2630 12010 2720 12250
rect 2960 12010 3050 12250
rect 3290 12010 3380 12250
rect 3620 12010 3710 12250
rect 3950 12010 4040 12250
rect 4280 12010 4370 12250
rect 4610 12010 4700 12250
rect 4940 12010 5030 12250
rect 5270 12010 5360 12250
rect 5600 12010 5690 12250
rect 5930 12010 6020 12250
rect 6260 12010 6350 12250
rect 6590 12010 6730 12250
rect -5510 11920 6730 12010
rect -5510 11680 -5200 11920
rect -4960 11680 -4870 11920
rect -4630 11680 -4540 11920
rect -4300 11680 -4210 11920
rect -3970 11680 -3880 11920
rect -3640 11680 -3550 11920
rect -3310 11680 -3220 11920
rect -2980 11680 -2890 11920
rect -2650 11680 -2560 11920
rect -2320 11680 -2230 11920
rect -1990 11680 -1900 11920
rect -1660 11680 -1570 11920
rect -1330 11680 -1240 11920
rect -1000 11680 -910 11920
rect -670 11680 -580 11920
rect -340 11680 -250 11920
rect -10 11680 80 11920
rect 320 11680 410 11920
rect 650 11680 740 11920
rect 980 11680 1070 11920
rect 1310 11680 1400 11920
rect 1640 11680 1730 11920
rect 1970 11680 2060 11920
rect 2300 11680 2390 11920
rect 2630 11680 2720 11920
rect 2960 11680 3050 11920
rect 3290 11680 3380 11920
rect 3620 11680 3710 11920
rect 3950 11680 4040 11920
rect 4280 11680 4370 11920
rect 4610 11680 4700 11920
rect 4940 11680 5030 11920
rect 5270 11680 5360 11920
rect 5600 11680 5690 11920
rect 5930 11680 6020 11920
rect 6260 11680 6350 11920
rect 6590 11680 6730 11920
rect -5510 11590 6730 11680
rect -5510 11350 -5200 11590
rect -4960 11350 -4870 11590
rect -4630 11350 -4540 11590
rect -4300 11350 -4210 11590
rect -3970 11350 -3880 11590
rect -3640 11350 -3550 11590
rect -3310 11350 -3220 11590
rect -2980 11350 -2890 11590
rect -2650 11350 -2560 11590
rect -2320 11350 -2230 11590
rect -1990 11350 -1900 11590
rect -1660 11350 -1570 11590
rect -1330 11350 -1240 11590
rect -1000 11350 -910 11590
rect -670 11350 -580 11590
rect -340 11350 -250 11590
rect -10 11350 80 11590
rect 320 11350 410 11590
rect 650 11350 740 11590
rect 980 11350 1070 11590
rect 1310 11350 1400 11590
rect 1640 11350 1730 11590
rect 1970 11350 2060 11590
rect 2300 11350 2390 11590
rect 2630 11350 2720 11590
rect 2960 11350 3050 11590
rect 3290 11350 3380 11590
rect 3620 11350 3710 11590
rect 3950 11350 4040 11590
rect 4280 11350 4370 11590
rect 4610 11350 4700 11590
rect 4940 11350 5030 11590
rect 5270 11350 5360 11590
rect 5600 11350 5690 11590
rect 5930 11350 6020 11590
rect 6260 11350 6350 11590
rect 6590 11350 6730 11590
rect -5510 11260 6730 11350
rect -5510 11020 -5200 11260
rect -4960 11020 -4870 11260
rect -4630 11020 -4540 11260
rect -4300 11020 -4210 11260
rect -3970 11020 -3880 11260
rect -3640 11020 -3550 11260
rect -3310 11020 -3220 11260
rect -2980 11020 -2890 11260
rect -2650 11020 -2560 11260
rect -2320 11020 -2230 11260
rect -1990 11020 -1900 11260
rect -1660 11020 -1570 11260
rect -1330 11020 -1240 11260
rect -1000 11020 -910 11260
rect -670 11020 -580 11260
rect -340 11020 -250 11260
rect -10 11020 80 11260
rect 320 11020 410 11260
rect 650 11020 740 11260
rect 980 11020 1070 11260
rect 1310 11020 1400 11260
rect 1640 11020 1730 11260
rect 1970 11020 2060 11260
rect 2300 11020 2390 11260
rect 2630 11020 2720 11260
rect 2960 11020 3050 11260
rect 3290 11020 3380 11260
rect 3620 11020 3710 11260
rect 3950 11020 4040 11260
rect 4280 11020 4370 11260
rect 4610 11020 4700 11260
rect 4940 11020 5030 11260
rect 5270 11020 5360 11260
rect 5600 11020 5690 11260
rect 5930 11020 6020 11260
rect 6260 11020 6350 11260
rect 6590 11020 6730 11260
rect -5510 10930 6730 11020
rect -5510 10690 -5200 10930
rect -4960 10690 -4870 10930
rect -4630 10690 -4540 10930
rect -4300 10690 -4210 10930
rect -3970 10690 -3880 10930
rect -3640 10690 -3550 10930
rect -3310 10690 -3220 10930
rect -2980 10690 -2890 10930
rect -2650 10690 -2560 10930
rect -2320 10690 -2230 10930
rect -1990 10690 -1900 10930
rect -1660 10690 -1570 10930
rect -1330 10690 -1240 10930
rect -1000 10690 -910 10930
rect -670 10690 -580 10930
rect -340 10690 -250 10930
rect -10 10690 80 10930
rect 320 10690 410 10930
rect 650 10690 740 10930
rect 980 10690 1070 10930
rect 1310 10690 1400 10930
rect 1640 10690 1730 10930
rect 1970 10690 2060 10930
rect 2300 10690 2390 10930
rect 2630 10690 2720 10930
rect 2960 10690 3050 10930
rect 3290 10690 3380 10930
rect 3620 10690 3710 10930
rect 3950 10690 4040 10930
rect 4280 10690 4370 10930
rect 4610 10690 4700 10930
rect 4940 10690 5030 10930
rect 5270 10690 5360 10930
rect 5600 10690 5690 10930
rect 5930 10690 6020 10930
rect 6260 10690 6350 10930
rect 6590 10690 6730 10930
rect -5510 10600 6730 10690
rect -5510 10360 -5200 10600
rect -4960 10360 -4870 10600
rect -4630 10360 -4540 10600
rect -4300 10360 -4210 10600
rect -3970 10360 -3880 10600
rect -3640 10360 -3550 10600
rect -3310 10360 -3220 10600
rect -2980 10360 -2890 10600
rect -2650 10360 -2560 10600
rect -2320 10360 -2230 10600
rect -1990 10360 -1900 10600
rect -1660 10360 -1570 10600
rect -1330 10360 -1240 10600
rect -1000 10360 -910 10600
rect -670 10360 -580 10600
rect -340 10360 -250 10600
rect -10 10360 80 10600
rect 320 10360 410 10600
rect 650 10360 740 10600
rect 980 10360 1070 10600
rect 1310 10360 1400 10600
rect 1640 10360 1730 10600
rect 1970 10360 2060 10600
rect 2300 10360 2390 10600
rect 2630 10360 2720 10600
rect 2960 10360 3050 10600
rect 3290 10360 3380 10600
rect 3620 10360 3710 10600
rect 3950 10360 4040 10600
rect 4280 10360 4370 10600
rect 4610 10360 4700 10600
rect 4940 10360 5030 10600
rect 5270 10360 5360 10600
rect 5600 10360 5690 10600
rect 5930 10360 6020 10600
rect 6260 10360 6350 10600
rect 6590 10360 6730 10600
rect -5510 10270 6730 10360
rect -5510 10030 -5200 10270
rect -4960 10030 -4870 10270
rect -4630 10030 -4540 10270
rect -4300 10030 -4210 10270
rect -3970 10030 -3880 10270
rect -3640 10030 -3550 10270
rect -3310 10030 -3220 10270
rect -2980 10030 -2890 10270
rect -2650 10030 -2560 10270
rect -2320 10030 -2230 10270
rect -1990 10030 -1900 10270
rect -1660 10030 -1570 10270
rect -1330 10030 -1240 10270
rect -1000 10030 -910 10270
rect -670 10030 -580 10270
rect -340 10030 -250 10270
rect -10 10030 80 10270
rect 320 10030 410 10270
rect 650 10030 740 10270
rect 980 10030 1070 10270
rect 1310 10030 1400 10270
rect 1640 10030 1730 10270
rect 1970 10030 2060 10270
rect 2300 10030 2390 10270
rect 2630 10030 2720 10270
rect 2960 10030 3050 10270
rect 3290 10030 3380 10270
rect 3620 10030 3710 10270
rect 3950 10030 4040 10270
rect 4280 10030 4370 10270
rect 4610 10030 4700 10270
rect 4940 10030 5030 10270
rect 5270 10030 5360 10270
rect 5600 10030 5690 10270
rect 5930 10030 6020 10270
rect 6260 10030 6350 10270
rect 6590 10030 6730 10270
rect -5510 9940 6730 10030
rect -5510 9700 -5200 9940
rect -4960 9700 -4870 9940
rect -4630 9700 -4540 9940
rect -4300 9700 -4210 9940
rect -3970 9700 -3880 9940
rect -3640 9700 -3550 9940
rect -3310 9700 -3220 9940
rect -2980 9700 -2890 9940
rect -2650 9700 -2560 9940
rect -2320 9700 -2230 9940
rect -1990 9700 -1900 9940
rect -1660 9700 -1570 9940
rect -1330 9700 -1240 9940
rect -1000 9700 -910 9940
rect -670 9700 -580 9940
rect -340 9700 -250 9940
rect -10 9700 80 9940
rect 320 9700 410 9940
rect 650 9700 740 9940
rect 980 9700 1070 9940
rect 1310 9700 1400 9940
rect 1640 9700 1730 9940
rect 1970 9700 2060 9940
rect 2300 9700 2390 9940
rect 2630 9700 2720 9940
rect 2960 9700 3050 9940
rect 3290 9700 3380 9940
rect 3620 9700 3710 9940
rect 3950 9700 4040 9940
rect 4280 9700 4370 9940
rect 4610 9700 4700 9940
rect 4940 9700 5030 9940
rect 5270 9700 5360 9940
rect 5600 9700 5690 9940
rect 5930 9700 6020 9940
rect 6260 9700 6350 9940
rect 6590 9700 6730 9940
rect -5510 9610 6730 9700
rect -5510 9370 -5200 9610
rect -4960 9370 -4870 9610
rect -4630 9370 -4540 9610
rect -4300 9370 -4210 9610
rect -3970 9370 -3880 9610
rect -3640 9370 -3550 9610
rect -3310 9370 -3220 9610
rect -2980 9370 -2890 9610
rect -2650 9370 -2560 9610
rect -2320 9370 -2230 9610
rect -1990 9370 -1900 9610
rect -1660 9370 -1570 9610
rect -1330 9370 -1240 9610
rect -1000 9370 -910 9610
rect -670 9370 -580 9610
rect -340 9370 -250 9610
rect -10 9370 80 9610
rect 320 9370 410 9610
rect 650 9370 740 9610
rect 980 9370 1070 9610
rect 1310 9370 1400 9610
rect 1640 9370 1730 9610
rect 1970 9370 2060 9610
rect 2300 9370 2390 9610
rect 2630 9370 2720 9610
rect 2960 9370 3050 9610
rect 3290 9370 3380 9610
rect 3620 9370 3710 9610
rect 3950 9370 4040 9610
rect 4280 9370 4370 9610
rect 4610 9370 4700 9610
rect 4940 9370 5030 9610
rect 5270 9370 5360 9610
rect 5600 9370 5690 9610
rect 5930 9370 6020 9610
rect 6260 9370 6350 9610
rect 6590 9370 6730 9610
rect -5510 9280 6730 9370
rect -5510 9040 -5200 9280
rect -4960 9040 -4870 9280
rect -4630 9040 -4540 9280
rect -4300 9040 -4210 9280
rect -3970 9040 -3880 9280
rect -3640 9040 -3550 9280
rect -3310 9040 -3220 9280
rect -2980 9040 -2890 9280
rect -2650 9040 -2560 9280
rect -2320 9040 -2230 9280
rect -1990 9040 -1900 9280
rect -1660 9040 -1570 9280
rect -1330 9040 -1240 9280
rect -1000 9040 -910 9280
rect -670 9040 -580 9280
rect -340 9040 -250 9280
rect -10 9040 80 9280
rect 320 9040 410 9280
rect 650 9040 740 9280
rect 980 9040 1070 9280
rect 1310 9040 1400 9280
rect 1640 9040 1730 9280
rect 1970 9040 2060 9280
rect 2300 9040 2390 9280
rect 2630 9040 2720 9280
rect 2960 9040 3050 9280
rect 3290 9040 3380 9280
rect 3620 9040 3710 9280
rect 3950 9040 4040 9280
rect 4280 9040 4370 9280
rect 4610 9040 4700 9280
rect 4940 9040 5030 9280
rect 5270 9040 5360 9280
rect 5600 9040 5690 9280
rect 5930 9040 6020 9280
rect 6260 9040 6350 9280
rect 6590 9040 6730 9280
rect -5510 8720 6730 9040
rect 8170 20830 20410 20960
rect 8170 20590 8310 20830
rect 8550 20590 8640 20830
rect 8880 20590 8970 20830
rect 9210 20590 9300 20830
rect 9540 20590 9630 20830
rect 9870 20590 9960 20830
rect 10200 20590 10290 20830
rect 10530 20590 10620 20830
rect 10860 20590 10950 20830
rect 11190 20590 11280 20830
rect 11520 20590 11610 20830
rect 11850 20590 11940 20830
rect 12180 20590 12270 20830
rect 12510 20590 12600 20830
rect 12840 20590 12930 20830
rect 13170 20590 13260 20830
rect 13500 20590 13590 20830
rect 13830 20590 13920 20830
rect 14160 20590 14250 20830
rect 14490 20590 14580 20830
rect 14820 20590 14910 20830
rect 15150 20590 15240 20830
rect 15480 20590 15570 20830
rect 15810 20590 15900 20830
rect 16140 20590 16230 20830
rect 16470 20590 16560 20830
rect 16800 20590 16890 20830
rect 17130 20590 17220 20830
rect 17460 20590 17550 20830
rect 17790 20590 17880 20830
rect 18120 20590 18210 20830
rect 18450 20590 18540 20830
rect 18780 20590 18870 20830
rect 19110 20590 19200 20830
rect 19440 20590 19530 20830
rect 19770 20590 19860 20830
rect 20100 20590 20410 20830
rect 8170 20500 20410 20590
rect 8170 20260 8310 20500
rect 8550 20260 8640 20500
rect 8880 20260 8970 20500
rect 9210 20260 9300 20500
rect 9540 20260 9630 20500
rect 9870 20260 9960 20500
rect 10200 20260 10290 20500
rect 10530 20260 10620 20500
rect 10860 20260 10950 20500
rect 11190 20260 11280 20500
rect 11520 20260 11610 20500
rect 11850 20260 11940 20500
rect 12180 20260 12270 20500
rect 12510 20260 12600 20500
rect 12840 20260 12930 20500
rect 13170 20260 13260 20500
rect 13500 20260 13590 20500
rect 13830 20260 13920 20500
rect 14160 20260 14250 20500
rect 14490 20260 14580 20500
rect 14820 20260 14910 20500
rect 15150 20260 15240 20500
rect 15480 20260 15570 20500
rect 15810 20260 15900 20500
rect 16140 20260 16230 20500
rect 16470 20260 16560 20500
rect 16800 20260 16890 20500
rect 17130 20260 17220 20500
rect 17460 20260 17550 20500
rect 17790 20260 17880 20500
rect 18120 20260 18210 20500
rect 18450 20260 18540 20500
rect 18780 20260 18870 20500
rect 19110 20260 19200 20500
rect 19440 20260 19530 20500
rect 19770 20260 19860 20500
rect 20100 20260 20410 20500
rect 8170 20170 20410 20260
rect 8170 19930 8310 20170
rect 8550 19930 8640 20170
rect 8880 19930 8970 20170
rect 9210 19930 9300 20170
rect 9540 19930 9630 20170
rect 9870 19930 9960 20170
rect 10200 19930 10290 20170
rect 10530 19930 10620 20170
rect 10860 19930 10950 20170
rect 11190 19930 11280 20170
rect 11520 19930 11610 20170
rect 11850 19930 11940 20170
rect 12180 19930 12270 20170
rect 12510 19930 12600 20170
rect 12840 19930 12930 20170
rect 13170 19930 13260 20170
rect 13500 19930 13590 20170
rect 13830 19930 13920 20170
rect 14160 19930 14250 20170
rect 14490 19930 14580 20170
rect 14820 19930 14910 20170
rect 15150 19930 15240 20170
rect 15480 19930 15570 20170
rect 15810 19930 15900 20170
rect 16140 19930 16230 20170
rect 16470 19930 16560 20170
rect 16800 19930 16890 20170
rect 17130 19930 17220 20170
rect 17460 19930 17550 20170
rect 17790 19930 17880 20170
rect 18120 19930 18210 20170
rect 18450 19930 18540 20170
rect 18780 19930 18870 20170
rect 19110 19930 19200 20170
rect 19440 19930 19530 20170
rect 19770 19930 19860 20170
rect 20100 19930 20410 20170
rect 8170 19840 20410 19930
rect 8170 19600 8310 19840
rect 8550 19600 8640 19840
rect 8880 19600 8970 19840
rect 9210 19600 9300 19840
rect 9540 19600 9630 19840
rect 9870 19600 9960 19840
rect 10200 19600 10290 19840
rect 10530 19600 10620 19840
rect 10860 19600 10950 19840
rect 11190 19600 11280 19840
rect 11520 19600 11610 19840
rect 11850 19600 11940 19840
rect 12180 19600 12270 19840
rect 12510 19600 12600 19840
rect 12840 19600 12930 19840
rect 13170 19600 13260 19840
rect 13500 19600 13590 19840
rect 13830 19600 13920 19840
rect 14160 19600 14250 19840
rect 14490 19600 14580 19840
rect 14820 19600 14910 19840
rect 15150 19600 15240 19840
rect 15480 19600 15570 19840
rect 15810 19600 15900 19840
rect 16140 19600 16230 19840
rect 16470 19600 16560 19840
rect 16800 19600 16890 19840
rect 17130 19600 17220 19840
rect 17460 19600 17550 19840
rect 17790 19600 17880 19840
rect 18120 19600 18210 19840
rect 18450 19600 18540 19840
rect 18780 19600 18870 19840
rect 19110 19600 19200 19840
rect 19440 19600 19530 19840
rect 19770 19600 19860 19840
rect 20100 19600 20410 19840
rect 8170 19510 20410 19600
rect 8170 19270 8310 19510
rect 8550 19270 8640 19510
rect 8880 19270 8970 19510
rect 9210 19270 9300 19510
rect 9540 19270 9630 19510
rect 9870 19270 9960 19510
rect 10200 19270 10290 19510
rect 10530 19270 10620 19510
rect 10860 19270 10950 19510
rect 11190 19270 11280 19510
rect 11520 19270 11610 19510
rect 11850 19270 11940 19510
rect 12180 19270 12270 19510
rect 12510 19270 12600 19510
rect 12840 19270 12930 19510
rect 13170 19270 13260 19510
rect 13500 19270 13590 19510
rect 13830 19270 13920 19510
rect 14160 19270 14250 19510
rect 14490 19270 14580 19510
rect 14820 19270 14910 19510
rect 15150 19270 15240 19510
rect 15480 19270 15570 19510
rect 15810 19270 15900 19510
rect 16140 19270 16230 19510
rect 16470 19270 16560 19510
rect 16800 19270 16890 19510
rect 17130 19270 17220 19510
rect 17460 19270 17550 19510
rect 17790 19270 17880 19510
rect 18120 19270 18210 19510
rect 18450 19270 18540 19510
rect 18780 19270 18870 19510
rect 19110 19270 19200 19510
rect 19440 19270 19530 19510
rect 19770 19270 19860 19510
rect 20100 19270 20410 19510
rect 8170 19180 20410 19270
rect 8170 18940 8310 19180
rect 8550 18940 8640 19180
rect 8880 18940 8970 19180
rect 9210 18940 9300 19180
rect 9540 18940 9630 19180
rect 9870 18940 9960 19180
rect 10200 18940 10290 19180
rect 10530 18940 10620 19180
rect 10860 18940 10950 19180
rect 11190 18940 11280 19180
rect 11520 18940 11610 19180
rect 11850 18940 11940 19180
rect 12180 18940 12270 19180
rect 12510 18940 12600 19180
rect 12840 18940 12930 19180
rect 13170 18940 13260 19180
rect 13500 18940 13590 19180
rect 13830 18940 13920 19180
rect 14160 18940 14250 19180
rect 14490 18940 14580 19180
rect 14820 18940 14910 19180
rect 15150 18940 15240 19180
rect 15480 18940 15570 19180
rect 15810 18940 15900 19180
rect 16140 18940 16230 19180
rect 16470 18940 16560 19180
rect 16800 18940 16890 19180
rect 17130 18940 17220 19180
rect 17460 18940 17550 19180
rect 17790 18940 17880 19180
rect 18120 18940 18210 19180
rect 18450 18940 18540 19180
rect 18780 18940 18870 19180
rect 19110 18940 19200 19180
rect 19440 18940 19530 19180
rect 19770 18940 19860 19180
rect 20100 18940 20410 19180
rect 8170 18850 20410 18940
rect 8170 18610 8310 18850
rect 8550 18610 8640 18850
rect 8880 18610 8970 18850
rect 9210 18610 9300 18850
rect 9540 18610 9630 18850
rect 9870 18610 9960 18850
rect 10200 18610 10290 18850
rect 10530 18610 10620 18850
rect 10860 18610 10950 18850
rect 11190 18610 11280 18850
rect 11520 18610 11610 18850
rect 11850 18610 11940 18850
rect 12180 18610 12270 18850
rect 12510 18610 12600 18850
rect 12840 18610 12930 18850
rect 13170 18610 13260 18850
rect 13500 18610 13590 18850
rect 13830 18610 13920 18850
rect 14160 18610 14250 18850
rect 14490 18610 14580 18850
rect 14820 18610 14910 18850
rect 15150 18610 15240 18850
rect 15480 18610 15570 18850
rect 15810 18610 15900 18850
rect 16140 18610 16230 18850
rect 16470 18610 16560 18850
rect 16800 18610 16890 18850
rect 17130 18610 17220 18850
rect 17460 18610 17550 18850
rect 17790 18610 17880 18850
rect 18120 18610 18210 18850
rect 18450 18610 18540 18850
rect 18780 18610 18870 18850
rect 19110 18610 19200 18850
rect 19440 18610 19530 18850
rect 19770 18610 19860 18850
rect 20100 18610 20410 18850
rect 8170 18520 20410 18610
rect 8170 18280 8310 18520
rect 8550 18280 8640 18520
rect 8880 18280 8970 18520
rect 9210 18280 9300 18520
rect 9540 18280 9630 18520
rect 9870 18280 9960 18520
rect 10200 18280 10290 18520
rect 10530 18280 10620 18520
rect 10860 18280 10950 18520
rect 11190 18280 11280 18520
rect 11520 18280 11610 18520
rect 11850 18280 11940 18520
rect 12180 18280 12270 18520
rect 12510 18280 12600 18520
rect 12840 18280 12930 18520
rect 13170 18280 13260 18520
rect 13500 18280 13590 18520
rect 13830 18280 13920 18520
rect 14160 18280 14250 18520
rect 14490 18280 14580 18520
rect 14820 18280 14910 18520
rect 15150 18280 15240 18520
rect 15480 18280 15570 18520
rect 15810 18280 15900 18520
rect 16140 18280 16230 18520
rect 16470 18280 16560 18520
rect 16800 18280 16890 18520
rect 17130 18280 17220 18520
rect 17460 18280 17550 18520
rect 17790 18280 17880 18520
rect 18120 18280 18210 18520
rect 18450 18280 18540 18520
rect 18780 18280 18870 18520
rect 19110 18280 19200 18520
rect 19440 18280 19530 18520
rect 19770 18280 19860 18520
rect 20100 18280 20410 18520
rect 8170 18190 20410 18280
rect 8170 17950 8310 18190
rect 8550 17950 8640 18190
rect 8880 17950 8970 18190
rect 9210 17950 9300 18190
rect 9540 17950 9630 18190
rect 9870 17950 9960 18190
rect 10200 17950 10290 18190
rect 10530 17950 10620 18190
rect 10860 17950 10950 18190
rect 11190 17950 11280 18190
rect 11520 17950 11610 18190
rect 11850 17950 11940 18190
rect 12180 17950 12270 18190
rect 12510 17950 12600 18190
rect 12840 17950 12930 18190
rect 13170 17950 13260 18190
rect 13500 17950 13590 18190
rect 13830 17950 13920 18190
rect 14160 17950 14250 18190
rect 14490 17950 14580 18190
rect 14820 17950 14910 18190
rect 15150 17950 15240 18190
rect 15480 17950 15570 18190
rect 15810 17950 15900 18190
rect 16140 17950 16230 18190
rect 16470 17950 16560 18190
rect 16800 17950 16890 18190
rect 17130 17950 17220 18190
rect 17460 17950 17550 18190
rect 17790 17950 17880 18190
rect 18120 17950 18210 18190
rect 18450 17950 18540 18190
rect 18780 17950 18870 18190
rect 19110 17950 19200 18190
rect 19440 17950 19530 18190
rect 19770 17950 19860 18190
rect 20100 17950 20410 18190
rect 8170 17860 20410 17950
rect 8170 17620 8310 17860
rect 8550 17620 8640 17860
rect 8880 17620 8970 17860
rect 9210 17620 9300 17860
rect 9540 17620 9630 17860
rect 9870 17620 9960 17860
rect 10200 17620 10290 17860
rect 10530 17620 10620 17860
rect 10860 17620 10950 17860
rect 11190 17620 11280 17860
rect 11520 17620 11610 17860
rect 11850 17620 11940 17860
rect 12180 17620 12270 17860
rect 12510 17620 12600 17860
rect 12840 17620 12930 17860
rect 13170 17620 13260 17860
rect 13500 17620 13590 17860
rect 13830 17620 13920 17860
rect 14160 17620 14250 17860
rect 14490 17620 14580 17860
rect 14820 17620 14910 17860
rect 15150 17620 15240 17860
rect 15480 17620 15570 17860
rect 15810 17620 15900 17860
rect 16140 17620 16230 17860
rect 16470 17620 16560 17860
rect 16800 17620 16890 17860
rect 17130 17620 17220 17860
rect 17460 17620 17550 17860
rect 17790 17620 17880 17860
rect 18120 17620 18210 17860
rect 18450 17620 18540 17860
rect 18780 17620 18870 17860
rect 19110 17620 19200 17860
rect 19440 17620 19530 17860
rect 19770 17620 19860 17860
rect 20100 17620 20410 17860
rect 8170 17530 20410 17620
rect 8170 17290 8310 17530
rect 8550 17290 8640 17530
rect 8880 17290 8970 17530
rect 9210 17290 9300 17530
rect 9540 17290 9630 17530
rect 9870 17290 9960 17530
rect 10200 17290 10290 17530
rect 10530 17290 10620 17530
rect 10860 17290 10950 17530
rect 11190 17290 11280 17530
rect 11520 17290 11610 17530
rect 11850 17290 11940 17530
rect 12180 17290 12270 17530
rect 12510 17290 12600 17530
rect 12840 17290 12930 17530
rect 13170 17290 13260 17530
rect 13500 17290 13590 17530
rect 13830 17290 13920 17530
rect 14160 17290 14250 17530
rect 14490 17290 14580 17530
rect 14820 17290 14910 17530
rect 15150 17290 15240 17530
rect 15480 17290 15570 17530
rect 15810 17290 15900 17530
rect 16140 17290 16230 17530
rect 16470 17290 16560 17530
rect 16800 17290 16890 17530
rect 17130 17290 17220 17530
rect 17460 17290 17550 17530
rect 17790 17290 17880 17530
rect 18120 17290 18210 17530
rect 18450 17290 18540 17530
rect 18780 17290 18870 17530
rect 19110 17290 19200 17530
rect 19440 17290 19530 17530
rect 19770 17290 19860 17530
rect 20100 17290 20410 17530
rect 8170 17200 20410 17290
rect 8170 16960 8310 17200
rect 8550 16960 8640 17200
rect 8880 16960 8970 17200
rect 9210 16960 9300 17200
rect 9540 16960 9630 17200
rect 9870 16960 9960 17200
rect 10200 16960 10290 17200
rect 10530 16960 10620 17200
rect 10860 16960 10950 17200
rect 11190 16960 11280 17200
rect 11520 16960 11610 17200
rect 11850 16960 11940 17200
rect 12180 16960 12270 17200
rect 12510 16960 12600 17200
rect 12840 16960 12930 17200
rect 13170 16960 13260 17200
rect 13500 16960 13590 17200
rect 13830 16960 13920 17200
rect 14160 16960 14250 17200
rect 14490 16960 14580 17200
rect 14820 16960 14910 17200
rect 15150 16960 15240 17200
rect 15480 16960 15570 17200
rect 15810 16960 15900 17200
rect 16140 16960 16230 17200
rect 16470 16960 16560 17200
rect 16800 16960 16890 17200
rect 17130 16960 17220 17200
rect 17460 16960 17550 17200
rect 17790 16960 17880 17200
rect 18120 16960 18210 17200
rect 18450 16960 18540 17200
rect 18780 16960 18870 17200
rect 19110 16960 19200 17200
rect 19440 16960 19530 17200
rect 19770 16960 19860 17200
rect 20100 16960 20410 17200
rect 8170 16870 20410 16960
rect 8170 16630 8310 16870
rect 8550 16630 8640 16870
rect 8880 16630 8970 16870
rect 9210 16630 9300 16870
rect 9540 16630 9630 16870
rect 9870 16630 9960 16870
rect 10200 16630 10290 16870
rect 10530 16630 10620 16870
rect 10860 16630 10950 16870
rect 11190 16630 11280 16870
rect 11520 16630 11610 16870
rect 11850 16630 11940 16870
rect 12180 16630 12270 16870
rect 12510 16630 12600 16870
rect 12840 16630 12930 16870
rect 13170 16630 13260 16870
rect 13500 16630 13590 16870
rect 13830 16630 13920 16870
rect 14160 16630 14250 16870
rect 14490 16630 14580 16870
rect 14820 16630 14910 16870
rect 15150 16630 15240 16870
rect 15480 16630 15570 16870
rect 15810 16630 15900 16870
rect 16140 16630 16230 16870
rect 16470 16630 16560 16870
rect 16800 16630 16890 16870
rect 17130 16630 17220 16870
rect 17460 16630 17550 16870
rect 17790 16630 17880 16870
rect 18120 16630 18210 16870
rect 18450 16630 18540 16870
rect 18780 16630 18870 16870
rect 19110 16630 19200 16870
rect 19440 16630 19530 16870
rect 19770 16630 19860 16870
rect 20100 16630 20410 16870
rect 8170 16540 20410 16630
rect 8170 16300 8310 16540
rect 8550 16300 8640 16540
rect 8880 16300 8970 16540
rect 9210 16300 9300 16540
rect 9540 16300 9630 16540
rect 9870 16300 9960 16540
rect 10200 16300 10290 16540
rect 10530 16300 10620 16540
rect 10860 16300 10950 16540
rect 11190 16300 11280 16540
rect 11520 16300 11610 16540
rect 11850 16300 11940 16540
rect 12180 16300 12270 16540
rect 12510 16300 12600 16540
rect 12840 16300 12930 16540
rect 13170 16300 13260 16540
rect 13500 16300 13590 16540
rect 13830 16300 13920 16540
rect 14160 16300 14250 16540
rect 14490 16300 14580 16540
rect 14820 16300 14910 16540
rect 15150 16300 15240 16540
rect 15480 16300 15570 16540
rect 15810 16300 15900 16540
rect 16140 16300 16230 16540
rect 16470 16300 16560 16540
rect 16800 16300 16890 16540
rect 17130 16300 17220 16540
rect 17460 16300 17550 16540
rect 17790 16300 17880 16540
rect 18120 16300 18210 16540
rect 18450 16300 18540 16540
rect 18780 16300 18870 16540
rect 19110 16300 19200 16540
rect 19440 16300 19530 16540
rect 19770 16300 19860 16540
rect 20100 16300 20410 16540
rect 8170 16210 20410 16300
rect 8170 15970 8310 16210
rect 8550 15970 8640 16210
rect 8880 15970 8970 16210
rect 9210 15970 9300 16210
rect 9540 15970 9630 16210
rect 9870 15970 9960 16210
rect 10200 15970 10290 16210
rect 10530 15970 10620 16210
rect 10860 15970 10950 16210
rect 11190 15970 11280 16210
rect 11520 15970 11610 16210
rect 11850 15970 11940 16210
rect 12180 15970 12270 16210
rect 12510 15970 12600 16210
rect 12840 15970 12930 16210
rect 13170 15970 13260 16210
rect 13500 15970 13590 16210
rect 13830 15970 13920 16210
rect 14160 15970 14250 16210
rect 14490 15970 14580 16210
rect 14820 15970 14910 16210
rect 15150 15970 15240 16210
rect 15480 15970 15570 16210
rect 15810 15970 15900 16210
rect 16140 15970 16230 16210
rect 16470 15970 16560 16210
rect 16800 15970 16890 16210
rect 17130 15970 17220 16210
rect 17460 15970 17550 16210
rect 17790 15970 17880 16210
rect 18120 15970 18210 16210
rect 18450 15970 18540 16210
rect 18780 15970 18870 16210
rect 19110 15970 19200 16210
rect 19440 15970 19530 16210
rect 19770 15970 19860 16210
rect 20100 15970 20410 16210
rect 8170 15880 20410 15970
rect 8170 15640 8310 15880
rect 8550 15640 8640 15880
rect 8880 15640 8970 15880
rect 9210 15640 9300 15880
rect 9540 15640 9630 15880
rect 9870 15640 9960 15880
rect 10200 15640 10290 15880
rect 10530 15640 10620 15880
rect 10860 15640 10950 15880
rect 11190 15640 11280 15880
rect 11520 15640 11610 15880
rect 11850 15640 11940 15880
rect 12180 15640 12270 15880
rect 12510 15640 12600 15880
rect 12840 15640 12930 15880
rect 13170 15640 13260 15880
rect 13500 15640 13590 15880
rect 13830 15640 13920 15880
rect 14160 15640 14250 15880
rect 14490 15640 14580 15880
rect 14820 15640 14910 15880
rect 15150 15640 15240 15880
rect 15480 15640 15570 15880
rect 15810 15640 15900 15880
rect 16140 15640 16230 15880
rect 16470 15640 16560 15880
rect 16800 15640 16890 15880
rect 17130 15640 17220 15880
rect 17460 15640 17550 15880
rect 17790 15640 17880 15880
rect 18120 15640 18210 15880
rect 18450 15640 18540 15880
rect 18780 15640 18870 15880
rect 19110 15640 19200 15880
rect 19440 15640 19530 15880
rect 19770 15640 19860 15880
rect 20100 15640 20410 15880
rect 8170 15550 20410 15640
rect 8170 15310 8310 15550
rect 8550 15310 8640 15550
rect 8880 15310 8970 15550
rect 9210 15310 9300 15550
rect 9540 15310 9630 15550
rect 9870 15310 9960 15550
rect 10200 15310 10290 15550
rect 10530 15310 10620 15550
rect 10860 15310 10950 15550
rect 11190 15310 11280 15550
rect 11520 15310 11610 15550
rect 11850 15310 11940 15550
rect 12180 15310 12270 15550
rect 12510 15310 12600 15550
rect 12840 15310 12930 15550
rect 13170 15310 13260 15550
rect 13500 15310 13590 15550
rect 13830 15310 13920 15550
rect 14160 15310 14250 15550
rect 14490 15310 14580 15550
rect 14820 15310 14910 15550
rect 15150 15310 15240 15550
rect 15480 15310 15570 15550
rect 15810 15310 15900 15550
rect 16140 15310 16230 15550
rect 16470 15310 16560 15550
rect 16800 15310 16890 15550
rect 17130 15310 17220 15550
rect 17460 15310 17550 15550
rect 17790 15310 17880 15550
rect 18120 15310 18210 15550
rect 18450 15310 18540 15550
rect 18780 15310 18870 15550
rect 19110 15310 19200 15550
rect 19440 15310 19530 15550
rect 19770 15310 19860 15550
rect 20100 15310 20410 15550
rect 8170 15220 20410 15310
rect 8170 14980 8310 15220
rect 8550 14980 8640 15220
rect 8880 14980 8970 15220
rect 9210 14980 9300 15220
rect 9540 14980 9630 15220
rect 9870 14980 9960 15220
rect 10200 14980 10290 15220
rect 10530 14980 10620 15220
rect 10860 14980 10950 15220
rect 11190 14980 11280 15220
rect 11520 14980 11610 15220
rect 11850 14980 11940 15220
rect 12180 14980 12270 15220
rect 12510 14980 12600 15220
rect 12840 14980 12930 15220
rect 13170 14980 13260 15220
rect 13500 14980 13590 15220
rect 13830 14980 13920 15220
rect 14160 14980 14250 15220
rect 14490 14980 14580 15220
rect 14820 14980 14910 15220
rect 15150 14980 15240 15220
rect 15480 14980 15570 15220
rect 15810 14980 15900 15220
rect 16140 14980 16230 15220
rect 16470 14980 16560 15220
rect 16800 14980 16890 15220
rect 17130 14980 17220 15220
rect 17460 14980 17550 15220
rect 17790 14980 17880 15220
rect 18120 14980 18210 15220
rect 18450 14980 18540 15220
rect 18780 14980 18870 15220
rect 19110 14980 19200 15220
rect 19440 14980 19530 15220
rect 19770 14980 19860 15220
rect 20100 14980 20410 15220
rect 8170 14890 20410 14980
rect 8170 14650 8310 14890
rect 8550 14650 8640 14890
rect 8880 14650 8970 14890
rect 9210 14650 9300 14890
rect 9540 14650 9630 14890
rect 9870 14650 9960 14890
rect 10200 14650 10290 14890
rect 10530 14650 10620 14890
rect 10860 14650 10950 14890
rect 11190 14650 11280 14890
rect 11520 14650 11610 14890
rect 11850 14650 11940 14890
rect 12180 14650 12270 14890
rect 12510 14650 12600 14890
rect 12840 14650 12930 14890
rect 13170 14650 13260 14890
rect 13500 14650 13590 14890
rect 13830 14650 13920 14890
rect 14160 14650 14250 14890
rect 14490 14650 14580 14890
rect 14820 14650 14910 14890
rect 15150 14650 15240 14890
rect 15480 14650 15570 14890
rect 15810 14650 15900 14890
rect 16140 14650 16230 14890
rect 16470 14650 16560 14890
rect 16800 14650 16890 14890
rect 17130 14650 17220 14890
rect 17460 14650 17550 14890
rect 17790 14650 17880 14890
rect 18120 14650 18210 14890
rect 18450 14650 18540 14890
rect 18780 14650 18870 14890
rect 19110 14650 19200 14890
rect 19440 14650 19530 14890
rect 19770 14650 19860 14890
rect 20100 14650 20410 14890
rect 8170 14560 20410 14650
rect 8170 14320 8310 14560
rect 8550 14320 8640 14560
rect 8880 14320 8970 14560
rect 9210 14320 9300 14560
rect 9540 14320 9630 14560
rect 9870 14320 9960 14560
rect 10200 14320 10290 14560
rect 10530 14320 10620 14560
rect 10860 14320 10950 14560
rect 11190 14320 11280 14560
rect 11520 14320 11610 14560
rect 11850 14320 11940 14560
rect 12180 14320 12270 14560
rect 12510 14320 12600 14560
rect 12840 14320 12930 14560
rect 13170 14320 13260 14560
rect 13500 14320 13590 14560
rect 13830 14320 13920 14560
rect 14160 14320 14250 14560
rect 14490 14320 14580 14560
rect 14820 14320 14910 14560
rect 15150 14320 15240 14560
rect 15480 14320 15570 14560
rect 15810 14320 15900 14560
rect 16140 14320 16230 14560
rect 16470 14320 16560 14560
rect 16800 14320 16890 14560
rect 17130 14320 17220 14560
rect 17460 14320 17550 14560
rect 17790 14320 17880 14560
rect 18120 14320 18210 14560
rect 18450 14320 18540 14560
rect 18780 14320 18870 14560
rect 19110 14320 19200 14560
rect 19440 14320 19530 14560
rect 19770 14320 19860 14560
rect 20100 14320 20410 14560
rect 8170 14230 20410 14320
rect 8170 13990 8310 14230
rect 8550 13990 8640 14230
rect 8880 13990 8970 14230
rect 9210 13990 9300 14230
rect 9540 13990 9630 14230
rect 9870 13990 9960 14230
rect 10200 13990 10290 14230
rect 10530 13990 10620 14230
rect 10860 13990 10950 14230
rect 11190 13990 11280 14230
rect 11520 13990 11610 14230
rect 11850 13990 11940 14230
rect 12180 13990 12270 14230
rect 12510 13990 12600 14230
rect 12840 13990 12930 14230
rect 13170 13990 13260 14230
rect 13500 13990 13590 14230
rect 13830 13990 13920 14230
rect 14160 13990 14250 14230
rect 14490 13990 14580 14230
rect 14820 13990 14910 14230
rect 15150 13990 15240 14230
rect 15480 13990 15570 14230
rect 15810 13990 15900 14230
rect 16140 13990 16230 14230
rect 16470 13990 16560 14230
rect 16800 13990 16890 14230
rect 17130 13990 17220 14230
rect 17460 13990 17550 14230
rect 17790 13990 17880 14230
rect 18120 13990 18210 14230
rect 18450 13990 18540 14230
rect 18780 13990 18870 14230
rect 19110 13990 19200 14230
rect 19440 13990 19530 14230
rect 19770 13990 19860 14230
rect 20100 13990 20410 14230
rect 8170 13900 20410 13990
rect 8170 13660 8310 13900
rect 8550 13660 8640 13900
rect 8880 13660 8970 13900
rect 9210 13660 9300 13900
rect 9540 13660 9630 13900
rect 9870 13660 9960 13900
rect 10200 13660 10290 13900
rect 10530 13660 10620 13900
rect 10860 13660 10950 13900
rect 11190 13660 11280 13900
rect 11520 13660 11610 13900
rect 11850 13660 11940 13900
rect 12180 13660 12270 13900
rect 12510 13660 12600 13900
rect 12840 13660 12930 13900
rect 13170 13660 13260 13900
rect 13500 13660 13590 13900
rect 13830 13660 13920 13900
rect 14160 13660 14250 13900
rect 14490 13660 14580 13900
rect 14820 13660 14910 13900
rect 15150 13660 15240 13900
rect 15480 13660 15570 13900
rect 15810 13660 15900 13900
rect 16140 13660 16230 13900
rect 16470 13660 16560 13900
rect 16800 13660 16890 13900
rect 17130 13660 17220 13900
rect 17460 13660 17550 13900
rect 17790 13660 17880 13900
rect 18120 13660 18210 13900
rect 18450 13660 18540 13900
rect 18780 13660 18870 13900
rect 19110 13660 19200 13900
rect 19440 13660 19530 13900
rect 19770 13660 19860 13900
rect 20100 13660 20410 13900
rect 8170 13570 20410 13660
rect 8170 13330 8310 13570
rect 8550 13330 8640 13570
rect 8880 13330 8970 13570
rect 9210 13330 9300 13570
rect 9540 13330 9630 13570
rect 9870 13330 9960 13570
rect 10200 13330 10290 13570
rect 10530 13330 10620 13570
rect 10860 13330 10950 13570
rect 11190 13330 11280 13570
rect 11520 13330 11610 13570
rect 11850 13330 11940 13570
rect 12180 13330 12270 13570
rect 12510 13330 12600 13570
rect 12840 13330 12930 13570
rect 13170 13330 13260 13570
rect 13500 13330 13590 13570
rect 13830 13330 13920 13570
rect 14160 13330 14250 13570
rect 14490 13330 14580 13570
rect 14820 13330 14910 13570
rect 15150 13330 15240 13570
rect 15480 13330 15570 13570
rect 15810 13330 15900 13570
rect 16140 13330 16230 13570
rect 16470 13330 16560 13570
rect 16800 13330 16890 13570
rect 17130 13330 17220 13570
rect 17460 13330 17550 13570
rect 17790 13330 17880 13570
rect 18120 13330 18210 13570
rect 18450 13330 18540 13570
rect 18780 13330 18870 13570
rect 19110 13330 19200 13570
rect 19440 13330 19530 13570
rect 19770 13330 19860 13570
rect 20100 13330 20410 13570
rect 8170 13240 20410 13330
rect 8170 13000 8310 13240
rect 8550 13000 8640 13240
rect 8880 13000 8970 13240
rect 9210 13000 9300 13240
rect 9540 13000 9630 13240
rect 9870 13000 9960 13240
rect 10200 13000 10290 13240
rect 10530 13000 10620 13240
rect 10860 13000 10950 13240
rect 11190 13000 11280 13240
rect 11520 13000 11610 13240
rect 11850 13000 11940 13240
rect 12180 13000 12270 13240
rect 12510 13000 12600 13240
rect 12840 13000 12930 13240
rect 13170 13000 13260 13240
rect 13500 13000 13590 13240
rect 13830 13000 13920 13240
rect 14160 13000 14250 13240
rect 14490 13000 14580 13240
rect 14820 13000 14910 13240
rect 15150 13000 15240 13240
rect 15480 13000 15570 13240
rect 15810 13000 15900 13240
rect 16140 13000 16230 13240
rect 16470 13000 16560 13240
rect 16800 13000 16890 13240
rect 17130 13000 17220 13240
rect 17460 13000 17550 13240
rect 17790 13000 17880 13240
rect 18120 13000 18210 13240
rect 18450 13000 18540 13240
rect 18780 13000 18870 13240
rect 19110 13000 19200 13240
rect 19440 13000 19530 13240
rect 19770 13000 19860 13240
rect 20100 13000 20410 13240
rect 8170 12910 20410 13000
rect 8170 12670 8310 12910
rect 8550 12670 8640 12910
rect 8880 12670 8970 12910
rect 9210 12670 9300 12910
rect 9540 12670 9630 12910
rect 9870 12670 9960 12910
rect 10200 12670 10290 12910
rect 10530 12670 10620 12910
rect 10860 12670 10950 12910
rect 11190 12670 11280 12910
rect 11520 12670 11610 12910
rect 11850 12670 11940 12910
rect 12180 12670 12270 12910
rect 12510 12670 12600 12910
rect 12840 12670 12930 12910
rect 13170 12670 13260 12910
rect 13500 12670 13590 12910
rect 13830 12670 13920 12910
rect 14160 12670 14250 12910
rect 14490 12670 14580 12910
rect 14820 12670 14910 12910
rect 15150 12670 15240 12910
rect 15480 12670 15570 12910
rect 15810 12670 15900 12910
rect 16140 12670 16230 12910
rect 16470 12670 16560 12910
rect 16800 12670 16890 12910
rect 17130 12670 17220 12910
rect 17460 12670 17550 12910
rect 17790 12670 17880 12910
rect 18120 12670 18210 12910
rect 18450 12670 18540 12910
rect 18780 12670 18870 12910
rect 19110 12670 19200 12910
rect 19440 12670 19530 12910
rect 19770 12670 19860 12910
rect 20100 12670 20410 12910
rect 8170 12580 20410 12670
rect 8170 12340 8310 12580
rect 8550 12340 8640 12580
rect 8880 12340 8970 12580
rect 9210 12340 9300 12580
rect 9540 12340 9630 12580
rect 9870 12340 9960 12580
rect 10200 12340 10290 12580
rect 10530 12340 10620 12580
rect 10860 12340 10950 12580
rect 11190 12340 11280 12580
rect 11520 12340 11610 12580
rect 11850 12340 11940 12580
rect 12180 12340 12270 12580
rect 12510 12340 12600 12580
rect 12840 12340 12930 12580
rect 13170 12340 13260 12580
rect 13500 12340 13590 12580
rect 13830 12340 13920 12580
rect 14160 12340 14250 12580
rect 14490 12340 14580 12580
rect 14820 12340 14910 12580
rect 15150 12340 15240 12580
rect 15480 12340 15570 12580
rect 15810 12340 15900 12580
rect 16140 12340 16230 12580
rect 16470 12340 16560 12580
rect 16800 12340 16890 12580
rect 17130 12340 17220 12580
rect 17460 12340 17550 12580
rect 17790 12340 17880 12580
rect 18120 12340 18210 12580
rect 18450 12340 18540 12580
rect 18780 12340 18870 12580
rect 19110 12340 19200 12580
rect 19440 12340 19530 12580
rect 19770 12340 19860 12580
rect 20100 12340 20410 12580
rect 8170 12250 20410 12340
rect 8170 12010 8310 12250
rect 8550 12010 8640 12250
rect 8880 12010 8970 12250
rect 9210 12010 9300 12250
rect 9540 12010 9630 12250
rect 9870 12010 9960 12250
rect 10200 12010 10290 12250
rect 10530 12010 10620 12250
rect 10860 12010 10950 12250
rect 11190 12010 11280 12250
rect 11520 12010 11610 12250
rect 11850 12010 11940 12250
rect 12180 12010 12270 12250
rect 12510 12010 12600 12250
rect 12840 12010 12930 12250
rect 13170 12010 13260 12250
rect 13500 12010 13590 12250
rect 13830 12010 13920 12250
rect 14160 12010 14250 12250
rect 14490 12010 14580 12250
rect 14820 12010 14910 12250
rect 15150 12010 15240 12250
rect 15480 12010 15570 12250
rect 15810 12010 15900 12250
rect 16140 12010 16230 12250
rect 16470 12010 16560 12250
rect 16800 12010 16890 12250
rect 17130 12010 17220 12250
rect 17460 12010 17550 12250
rect 17790 12010 17880 12250
rect 18120 12010 18210 12250
rect 18450 12010 18540 12250
rect 18780 12010 18870 12250
rect 19110 12010 19200 12250
rect 19440 12010 19530 12250
rect 19770 12010 19860 12250
rect 20100 12010 20410 12250
rect 8170 11920 20410 12010
rect 8170 11680 8310 11920
rect 8550 11680 8640 11920
rect 8880 11680 8970 11920
rect 9210 11680 9300 11920
rect 9540 11680 9630 11920
rect 9870 11680 9960 11920
rect 10200 11680 10290 11920
rect 10530 11680 10620 11920
rect 10860 11680 10950 11920
rect 11190 11680 11280 11920
rect 11520 11680 11610 11920
rect 11850 11680 11940 11920
rect 12180 11680 12270 11920
rect 12510 11680 12600 11920
rect 12840 11680 12930 11920
rect 13170 11680 13260 11920
rect 13500 11680 13590 11920
rect 13830 11680 13920 11920
rect 14160 11680 14250 11920
rect 14490 11680 14580 11920
rect 14820 11680 14910 11920
rect 15150 11680 15240 11920
rect 15480 11680 15570 11920
rect 15810 11680 15900 11920
rect 16140 11680 16230 11920
rect 16470 11680 16560 11920
rect 16800 11680 16890 11920
rect 17130 11680 17220 11920
rect 17460 11680 17550 11920
rect 17790 11680 17880 11920
rect 18120 11680 18210 11920
rect 18450 11680 18540 11920
rect 18780 11680 18870 11920
rect 19110 11680 19200 11920
rect 19440 11680 19530 11920
rect 19770 11680 19860 11920
rect 20100 11680 20410 11920
rect 8170 11590 20410 11680
rect 8170 11350 8310 11590
rect 8550 11350 8640 11590
rect 8880 11350 8970 11590
rect 9210 11350 9300 11590
rect 9540 11350 9630 11590
rect 9870 11350 9960 11590
rect 10200 11350 10290 11590
rect 10530 11350 10620 11590
rect 10860 11350 10950 11590
rect 11190 11350 11280 11590
rect 11520 11350 11610 11590
rect 11850 11350 11940 11590
rect 12180 11350 12270 11590
rect 12510 11350 12600 11590
rect 12840 11350 12930 11590
rect 13170 11350 13260 11590
rect 13500 11350 13590 11590
rect 13830 11350 13920 11590
rect 14160 11350 14250 11590
rect 14490 11350 14580 11590
rect 14820 11350 14910 11590
rect 15150 11350 15240 11590
rect 15480 11350 15570 11590
rect 15810 11350 15900 11590
rect 16140 11350 16230 11590
rect 16470 11350 16560 11590
rect 16800 11350 16890 11590
rect 17130 11350 17220 11590
rect 17460 11350 17550 11590
rect 17790 11350 17880 11590
rect 18120 11350 18210 11590
rect 18450 11350 18540 11590
rect 18780 11350 18870 11590
rect 19110 11350 19200 11590
rect 19440 11350 19530 11590
rect 19770 11350 19860 11590
rect 20100 11350 20410 11590
rect 8170 11260 20410 11350
rect 8170 11020 8310 11260
rect 8550 11020 8640 11260
rect 8880 11020 8970 11260
rect 9210 11020 9300 11260
rect 9540 11020 9630 11260
rect 9870 11020 9960 11260
rect 10200 11020 10290 11260
rect 10530 11020 10620 11260
rect 10860 11020 10950 11260
rect 11190 11020 11280 11260
rect 11520 11020 11610 11260
rect 11850 11020 11940 11260
rect 12180 11020 12270 11260
rect 12510 11020 12600 11260
rect 12840 11020 12930 11260
rect 13170 11020 13260 11260
rect 13500 11020 13590 11260
rect 13830 11020 13920 11260
rect 14160 11020 14250 11260
rect 14490 11020 14580 11260
rect 14820 11020 14910 11260
rect 15150 11020 15240 11260
rect 15480 11020 15570 11260
rect 15810 11020 15900 11260
rect 16140 11020 16230 11260
rect 16470 11020 16560 11260
rect 16800 11020 16890 11260
rect 17130 11020 17220 11260
rect 17460 11020 17550 11260
rect 17790 11020 17880 11260
rect 18120 11020 18210 11260
rect 18450 11020 18540 11260
rect 18780 11020 18870 11260
rect 19110 11020 19200 11260
rect 19440 11020 19530 11260
rect 19770 11020 19860 11260
rect 20100 11020 20410 11260
rect 8170 10930 20410 11020
rect 8170 10690 8310 10930
rect 8550 10690 8640 10930
rect 8880 10690 8970 10930
rect 9210 10690 9300 10930
rect 9540 10690 9630 10930
rect 9870 10690 9960 10930
rect 10200 10690 10290 10930
rect 10530 10690 10620 10930
rect 10860 10690 10950 10930
rect 11190 10690 11280 10930
rect 11520 10690 11610 10930
rect 11850 10690 11940 10930
rect 12180 10690 12270 10930
rect 12510 10690 12600 10930
rect 12840 10690 12930 10930
rect 13170 10690 13260 10930
rect 13500 10690 13590 10930
rect 13830 10690 13920 10930
rect 14160 10690 14250 10930
rect 14490 10690 14580 10930
rect 14820 10690 14910 10930
rect 15150 10690 15240 10930
rect 15480 10690 15570 10930
rect 15810 10690 15900 10930
rect 16140 10690 16230 10930
rect 16470 10690 16560 10930
rect 16800 10690 16890 10930
rect 17130 10690 17220 10930
rect 17460 10690 17550 10930
rect 17790 10690 17880 10930
rect 18120 10690 18210 10930
rect 18450 10690 18540 10930
rect 18780 10690 18870 10930
rect 19110 10690 19200 10930
rect 19440 10690 19530 10930
rect 19770 10690 19860 10930
rect 20100 10690 20410 10930
rect 8170 10600 20410 10690
rect 8170 10360 8310 10600
rect 8550 10360 8640 10600
rect 8880 10360 8970 10600
rect 9210 10360 9300 10600
rect 9540 10360 9630 10600
rect 9870 10360 9960 10600
rect 10200 10360 10290 10600
rect 10530 10360 10620 10600
rect 10860 10360 10950 10600
rect 11190 10360 11280 10600
rect 11520 10360 11610 10600
rect 11850 10360 11940 10600
rect 12180 10360 12270 10600
rect 12510 10360 12600 10600
rect 12840 10360 12930 10600
rect 13170 10360 13260 10600
rect 13500 10360 13590 10600
rect 13830 10360 13920 10600
rect 14160 10360 14250 10600
rect 14490 10360 14580 10600
rect 14820 10360 14910 10600
rect 15150 10360 15240 10600
rect 15480 10360 15570 10600
rect 15810 10360 15900 10600
rect 16140 10360 16230 10600
rect 16470 10360 16560 10600
rect 16800 10360 16890 10600
rect 17130 10360 17220 10600
rect 17460 10360 17550 10600
rect 17790 10360 17880 10600
rect 18120 10360 18210 10600
rect 18450 10360 18540 10600
rect 18780 10360 18870 10600
rect 19110 10360 19200 10600
rect 19440 10360 19530 10600
rect 19770 10360 19860 10600
rect 20100 10360 20410 10600
rect 8170 10270 20410 10360
rect 8170 10030 8310 10270
rect 8550 10030 8640 10270
rect 8880 10030 8970 10270
rect 9210 10030 9300 10270
rect 9540 10030 9630 10270
rect 9870 10030 9960 10270
rect 10200 10030 10290 10270
rect 10530 10030 10620 10270
rect 10860 10030 10950 10270
rect 11190 10030 11280 10270
rect 11520 10030 11610 10270
rect 11850 10030 11940 10270
rect 12180 10030 12270 10270
rect 12510 10030 12600 10270
rect 12840 10030 12930 10270
rect 13170 10030 13260 10270
rect 13500 10030 13590 10270
rect 13830 10030 13920 10270
rect 14160 10030 14250 10270
rect 14490 10030 14580 10270
rect 14820 10030 14910 10270
rect 15150 10030 15240 10270
rect 15480 10030 15570 10270
rect 15810 10030 15900 10270
rect 16140 10030 16230 10270
rect 16470 10030 16560 10270
rect 16800 10030 16890 10270
rect 17130 10030 17220 10270
rect 17460 10030 17550 10270
rect 17790 10030 17880 10270
rect 18120 10030 18210 10270
rect 18450 10030 18540 10270
rect 18780 10030 18870 10270
rect 19110 10030 19200 10270
rect 19440 10030 19530 10270
rect 19770 10030 19860 10270
rect 20100 10030 20410 10270
rect 8170 9940 20410 10030
rect 8170 9700 8310 9940
rect 8550 9700 8640 9940
rect 8880 9700 8970 9940
rect 9210 9700 9300 9940
rect 9540 9700 9630 9940
rect 9870 9700 9960 9940
rect 10200 9700 10290 9940
rect 10530 9700 10620 9940
rect 10860 9700 10950 9940
rect 11190 9700 11280 9940
rect 11520 9700 11610 9940
rect 11850 9700 11940 9940
rect 12180 9700 12270 9940
rect 12510 9700 12600 9940
rect 12840 9700 12930 9940
rect 13170 9700 13260 9940
rect 13500 9700 13590 9940
rect 13830 9700 13920 9940
rect 14160 9700 14250 9940
rect 14490 9700 14580 9940
rect 14820 9700 14910 9940
rect 15150 9700 15240 9940
rect 15480 9700 15570 9940
rect 15810 9700 15900 9940
rect 16140 9700 16230 9940
rect 16470 9700 16560 9940
rect 16800 9700 16890 9940
rect 17130 9700 17220 9940
rect 17460 9700 17550 9940
rect 17790 9700 17880 9940
rect 18120 9700 18210 9940
rect 18450 9700 18540 9940
rect 18780 9700 18870 9940
rect 19110 9700 19200 9940
rect 19440 9700 19530 9940
rect 19770 9700 19860 9940
rect 20100 9700 20410 9940
rect 8170 9610 20410 9700
rect 8170 9370 8310 9610
rect 8550 9370 8640 9610
rect 8880 9370 8970 9610
rect 9210 9370 9300 9610
rect 9540 9370 9630 9610
rect 9870 9370 9960 9610
rect 10200 9370 10290 9610
rect 10530 9370 10620 9610
rect 10860 9370 10950 9610
rect 11190 9370 11280 9610
rect 11520 9370 11610 9610
rect 11850 9370 11940 9610
rect 12180 9370 12270 9610
rect 12510 9370 12600 9610
rect 12840 9370 12930 9610
rect 13170 9370 13260 9610
rect 13500 9370 13590 9610
rect 13830 9370 13920 9610
rect 14160 9370 14250 9610
rect 14490 9370 14580 9610
rect 14820 9370 14910 9610
rect 15150 9370 15240 9610
rect 15480 9370 15570 9610
rect 15810 9370 15900 9610
rect 16140 9370 16230 9610
rect 16470 9370 16560 9610
rect 16800 9370 16890 9610
rect 17130 9370 17220 9610
rect 17460 9370 17550 9610
rect 17790 9370 17880 9610
rect 18120 9370 18210 9610
rect 18450 9370 18540 9610
rect 18780 9370 18870 9610
rect 19110 9370 19200 9610
rect 19440 9370 19530 9610
rect 19770 9370 19860 9610
rect 20100 9370 20410 9610
rect 8170 9280 20410 9370
rect 8170 9040 8310 9280
rect 8550 9040 8640 9280
rect 8880 9040 8970 9280
rect 9210 9040 9300 9280
rect 9540 9040 9630 9280
rect 9870 9040 9960 9280
rect 10200 9040 10290 9280
rect 10530 9040 10620 9280
rect 10860 9040 10950 9280
rect 11190 9040 11280 9280
rect 11520 9040 11610 9280
rect 11850 9040 11940 9280
rect 12180 9040 12270 9280
rect 12510 9040 12600 9280
rect 12840 9040 12930 9280
rect 13170 9040 13260 9280
rect 13500 9040 13590 9280
rect 13830 9040 13920 9280
rect 14160 9040 14250 9280
rect 14490 9040 14580 9280
rect 14820 9040 14910 9280
rect 15150 9040 15240 9280
rect 15480 9040 15570 9280
rect 15810 9040 15900 9280
rect 16140 9040 16230 9280
rect 16470 9040 16560 9280
rect 16800 9040 16890 9280
rect 17130 9040 17220 9280
rect 17460 9040 17550 9280
rect 17790 9040 17880 9280
rect 18120 9040 18210 9280
rect 18450 9040 18540 9280
rect 18780 9040 18870 9280
rect 19110 9040 19200 9280
rect 19440 9040 19530 9280
rect 19770 9040 19860 9280
rect 20100 9040 20410 9280
rect 8170 8720 20410 9040
rect 31130 7830 37830 7880
rect 31130 7590 31180 7830
rect 31420 7590 31510 7830
rect 31750 7590 31840 7830
rect 32080 7590 32170 7830
rect 32410 7590 32500 7830
rect 32740 7590 32830 7830
rect 33070 7590 33160 7830
rect 33400 7590 33490 7830
rect 33730 7590 33820 7830
rect 34060 7590 34150 7830
rect 34390 7590 34480 7830
rect 34720 7590 34810 7830
rect 35050 7590 35140 7830
rect 35380 7590 35470 7830
rect 35710 7590 35800 7830
rect 36040 7590 36130 7830
rect 36370 7590 36460 7830
rect 36700 7590 36790 7830
rect 37030 7590 37120 7830
rect 37360 7590 37450 7830
rect 37690 7590 37830 7830
rect 31130 7500 37830 7590
rect 31130 7260 31180 7500
rect 31420 7260 31510 7500
rect 31750 7260 31840 7500
rect 32080 7260 32170 7500
rect 32410 7260 32500 7500
rect 32740 7260 32830 7500
rect 33070 7260 33160 7500
rect 33400 7260 33490 7500
rect 33730 7260 33820 7500
rect 34060 7260 34150 7500
rect 34390 7260 34480 7500
rect 34720 7260 34810 7500
rect 35050 7260 35140 7500
rect 35380 7260 35470 7500
rect 35710 7260 35800 7500
rect 36040 7260 36130 7500
rect 36370 7260 36460 7500
rect 36700 7260 36790 7500
rect 37030 7260 37120 7500
rect 37360 7260 37450 7500
rect 37690 7260 37830 7500
rect 31130 7170 37830 7260
rect 31130 6930 31180 7170
rect 31420 6930 31510 7170
rect 31750 6930 31840 7170
rect 32080 6930 32170 7170
rect 32410 6930 32500 7170
rect 32740 6930 32830 7170
rect 33070 6930 33160 7170
rect 33400 6930 33490 7170
rect 33730 6930 33820 7170
rect 34060 6930 34150 7170
rect 34390 6930 34480 7170
rect 34720 6930 34810 7170
rect 35050 6930 35140 7170
rect 35380 6930 35470 7170
rect 35710 6930 35800 7170
rect 36040 6930 36130 7170
rect 36370 6930 36460 7170
rect 36700 6930 36790 7170
rect 37030 6930 37120 7170
rect 37360 6930 37450 7170
rect 37690 6930 37830 7170
rect 31130 6840 37830 6930
rect 31130 6600 31180 6840
rect 31420 6600 31510 6840
rect 31750 6600 31840 6840
rect 32080 6600 32170 6840
rect 32410 6600 32500 6840
rect 32740 6600 32830 6840
rect 33070 6600 33160 6840
rect 33400 6600 33490 6840
rect 33730 6600 33820 6840
rect 34060 6600 34150 6840
rect 34390 6600 34480 6840
rect 34720 6600 34810 6840
rect 35050 6600 35140 6840
rect 35380 6600 35470 6840
rect 35710 6600 35800 6840
rect 36040 6600 36130 6840
rect 36370 6600 36460 6840
rect 36700 6600 36790 6840
rect 37030 6600 37120 6840
rect 37360 6600 37450 6840
rect 37690 6600 37830 6840
rect 31130 6510 37830 6600
rect 31130 6270 31180 6510
rect 31420 6270 31510 6510
rect 31750 6270 31840 6510
rect 32080 6270 32170 6510
rect 32410 6270 32500 6510
rect 32740 6270 32830 6510
rect 33070 6270 33160 6510
rect 33400 6270 33490 6510
rect 33730 6270 33820 6510
rect 34060 6270 34150 6510
rect 34390 6270 34480 6510
rect 34720 6270 34810 6510
rect 35050 6270 35140 6510
rect 35380 6270 35470 6510
rect 35710 6270 35800 6510
rect 36040 6270 36130 6510
rect 36370 6270 36460 6510
rect 36700 6270 36790 6510
rect 37030 6270 37120 6510
rect 37360 6270 37450 6510
rect 37690 6270 37830 6510
rect 31130 6180 37830 6270
rect 31130 5940 31180 6180
rect 31420 5940 31510 6180
rect 31750 5940 31840 6180
rect 32080 5940 32170 6180
rect 32410 5940 32500 6180
rect 32740 5940 32830 6180
rect 33070 5940 33160 6180
rect 33400 5940 33490 6180
rect 33730 5940 33820 6180
rect 34060 5940 34150 6180
rect 34390 5940 34480 6180
rect 34720 5940 34810 6180
rect 35050 5940 35140 6180
rect 35380 5940 35470 6180
rect 35710 5940 35800 6180
rect 36040 5940 36130 6180
rect 36370 5940 36460 6180
rect 36700 5940 36790 6180
rect 37030 5940 37120 6180
rect 37360 5940 37450 6180
rect 37690 5940 37830 6180
rect 31130 5850 37830 5940
rect 31130 5610 31180 5850
rect 31420 5610 31510 5850
rect 31750 5610 31840 5850
rect 32080 5610 32170 5850
rect 32410 5610 32500 5850
rect 32740 5610 32830 5850
rect 33070 5610 33160 5850
rect 33400 5610 33490 5850
rect 33730 5610 33820 5850
rect 34060 5610 34150 5850
rect 34390 5610 34480 5850
rect 34720 5610 34810 5850
rect 35050 5610 35140 5850
rect 35380 5610 35470 5850
rect 35710 5610 35800 5850
rect 36040 5610 36130 5850
rect 36370 5610 36460 5850
rect 36700 5610 36790 5850
rect 37030 5610 37120 5850
rect 37360 5610 37450 5850
rect 37690 5610 37830 5850
rect 31130 5520 37830 5610
rect 31130 5280 31180 5520
rect 31420 5280 31510 5520
rect 31750 5280 31840 5520
rect 32080 5280 32170 5520
rect 32410 5280 32500 5520
rect 32740 5280 32830 5520
rect 33070 5280 33160 5520
rect 33400 5280 33490 5520
rect 33730 5280 33820 5520
rect 34060 5280 34150 5520
rect 34390 5280 34480 5520
rect 34720 5280 34810 5520
rect 35050 5280 35140 5520
rect 35380 5280 35470 5520
rect 35710 5280 35800 5520
rect 36040 5280 36130 5520
rect 36370 5280 36460 5520
rect 36700 5280 36790 5520
rect 37030 5280 37120 5520
rect 37360 5280 37450 5520
rect 37690 5280 37830 5520
rect 31130 5190 37830 5280
rect 31130 4950 31180 5190
rect 31420 4950 31510 5190
rect 31750 4950 31840 5190
rect 32080 4950 32170 5190
rect 32410 4950 32500 5190
rect 32740 4950 32830 5190
rect 33070 4950 33160 5190
rect 33400 4950 33490 5190
rect 33730 4950 33820 5190
rect 34060 4950 34150 5190
rect 34390 4950 34480 5190
rect 34720 4950 34810 5190
rect 35050 4950 35140 5190
rect 35380 4950 35470 5190
rect 35710 4950 35800 5190
rect 36040 4950 36130 5190
rect 36370 4950 36460 5190
rect 36700 4950 36790 5190
rect 37030 4950 37120 5190
rect 37360 4950 37450 5190
rect 37690 4950 37830 5190
rect 31130 4860 37830 4950
rect 31130 4620 31180 4860
rect 31420 4620 31510 4860
rect 31750 4620 31840 4860
rect 32080 4620 32170 4860
rect 32410 4620 32500 4860
rect 32740 4620 32830 4860
rect 33070 4620 33160 4860
rect 33400 4620 33490 4860
rect 33730 4620 33820 4860
rect 34060 4620 34150 4860
rect 34390 4620 34480 4860
rect 34720 4620 34810 4860
rect 35050 4620 35140 4860
rect 35380 4620 35470 4860
rect 35710 4620 35800 4860
rect 36040 4620 36130 4860
rect 36370 4620 36460 4860
rect 36700 4620 36790 4860
rect 37030 4620 37120 4860
rect 37360 4620 37450 4860
rect 37690 4620 37830 4860
rect 31130 4530 37830 4620
rect 31130 4290 31180 4530
rect 31420 4290 31510 4530
rect 31750 4290 31840 4530
rect 32080 4290 32170 4530
rect 32410 4290 32500 4530
rect 32740 4290 32830 4530
rect 33070 4290 33160 4530
rect 33400 4290 33490 4530
rect 33730 4290 33820 4530
rect 34060 4290 34150 4530
rect 34390 4290 34480 4530
rect 34720 4290 34810 4530
rect 35050 4290 35140 4530
rect 35380 4290 35470 4530
rect 35710 4290 35800 4530
rect 36040 4290 36130 4530
rect 36370 4290 36460 4530
rect 36700 4290 36790 4530
rect 37030 4290 37120 4530
rect 37360 4290 37450 4530
rect 37690 4290 37830 4530
rect 31130 4200 37830 4290
rect 31130 3960 31180 4200
rect 31420 3960 31510 4200
rect 31750 3960 31840 4200
rect 32080 3960 32170 4200
rect 32410 3960 32500 4200
rect 32740 3960 32830 4200
rect 33070 3960 33160 4200
rect 33400 3960 33490 4200
rect 33730 3960 33820 4200
rect 34060 3960 34150 4200
rect 34390 3960 34480 4200
rect 34720 3960 34810 4200
rect 35050 3960 35140 4200
rect 35380 3960 35470 4200
rect 35710 3960 35800 4200
rect 36040 3960 36130 4200
rect 36370 3960 36460 4200
rect 36700 3960 36790 4200
rect 37030 3960 37120 4200
rect 37360 3960 37450 4200
rect 37690 3960 37830 4200
rect 31130 3870 37830 3960
rect 31130 3630 31180 3870
rect 31420 3630 31510 3870
rect 31750 3630 31840 3870
rect 32080 3630 32170 3870
rect 32410 3630 32500 3870
rect 32740 3630 32830 3870
rect 33070 3630 33160 3870
rect 33400 3630 33490 3870
rect 33730 3630 33820 3870
rect 34060 3630 34150 3870
rect 34390 3630 34480 3870
rect 34720 3630 34810 3870
rect 35050 3630 35140 3870
rect 35380 3630 35470 3870
rect 35710 3630 35800 3870
rect 36040 3630 36130 3870
rect 36370 3630 36460 3870
rect 36700 3630 36790 3870
rect 37030 3630 37120 3870
rect 37360 3630 37450 3870
rect 37690 3630 37830 3870
rect 31130 3540 37830 3630
rect 31130 3300 31180 3540
rect 31420 3300 31510 3540
rect 31750 3300 31840 3540
rect 32080 3300 32170 3540
rect 32410 3300 32500 3540
rect 32740 3300 32830 3540
rect 33070 3300 33160 3540
rect 33400 3300 33490 3540
rect 33730 3300 33820 3540
rect 34060 3300 34150 3540
rect 34390 3300 34480 3540
rect 34720 3300 34810 3540
rect 35050 3300 35140 3540
rect 35380 3300 35470 3540
rect 35710 3300 35800 3540
rect 36040 3300 36130 3540
rect 36370 3300 36460 3540
rect 36700 3300 36790 3540
rect 37030 3300 37120 3540
rect 37360 3300 37450 3540
rect 37690 3300 37830 3540
rect 31130 3210 37830 3300
rect 31130 2970 31180 3210
rect 31420 2970 31510 3210
rect 31750 2970 31840 3210
rect 32080 2970 32170 3210
rect 32410 2970 32500 3210
rect 32740 2970 32830 3210
rect 33070 2970 33160 3210
rect 33400 2970 33490 3210
rect 33730 2970 33820 3210
rect 34060 2970 34150 3210
rect 34390 2970 34480 3210
rect 34720 2970 34810 3210
rect 35050 2970 35140 3210
rect 35380 2970 35470 3210
rect 35710 2970 35800 3210
rect 36040 2970 36130 3210
rect 36370 2970 36460 3210
rect 36700 2970 36790 3210
rect 37030 2970 37120 3210
rect 37360 2970 37450 3210
rect 37690 2970 37830 3210
rect 31130 2880 37830 2970
rect 31130 2640 31180 2880
rect 31420 2640 31510 2880
rect 31750 2640 31840 2880
rect 32080 2640 32170 2880
rect 32410 2640 32500 2880
rect 32740 2640 32830 2880
rect 33070 2640 33160 2880
rect 33400 2640 33490 2880
rect 33730 2640 33820 2880
rect 34060 2640 34150 2880
rect 34390 2640 34480 2880
rect 34720 2640 34810 2880
rect 35050 2640 35140 2880
rect 35380 2640 35470 2880
rect 35710 2640 35800 2880
rect 36040 2640 36130 2880
rect 36370 2640 36460 2880
rect 36700 2640 36790 2880
rect 37030 2640 37120 2880
rect 37360 2640 37450 2880
rect 37690 2640 37830 2880
rect 31130 2550 37830 2640
rect 31130 2310 31180 2550
rect 31420 2310 31510 2550
rect 31750 2310 31840 2550
rect 32080 2310 32170 2550
rect 32410 2310 32500 2550
rect 32740 2310 32830 2550
rect 33070 2310 33160 2550
rect 33400 2310 33490 2550
rect 33730 2310 33820 2550
rect 34060 2310 34150 2550
rect 34390 2310 34480 2550
rect 34720 2310 34810 2550
rect 35050 2310 35140 2550
rect 35380 2310 35470 2550
rect 35710 2310 35800 2550
rect 36040 2310 36130 2550
rect 36370 2310 36460 2550
rect 36700 2310 36790 2550
rect 37030 2310 37120 2550
rect 37360 2310 37450 2550
rect 37690 2310 37830 2550
rect 31130 2220 37830 2310
rect 31130 1980 31180 2220
rect 31420 1980 31510 2220
rect 31750 1980 31840 2220
rect 32080 1980 32170 2220
rect 32410 1980 32500 2220
rect 32740 1980 32830 2220
rect 33070 1980 33160 2220
rect 33400 1980 33490 2220
rect 33730 1980 33820 2220
rect 34060 1980 34150 2220
rect 34390 1980 34480 2220
rect 34720 1980 34810 2220
rect 35050 1980 35140 2220
rect 35380 1980 35470 2220
rect 35710 1980 35800 2220
rect 36040 1980 36130 2220
rect 36370 1980 36460 2220
rect 36700 1980 36790 2220
rect 37030 1980 37120 2220
rect 37360 1980 37450 2220
rect 37690 1980 37830 2220
rect 31130 1890 37830 1980
rect 31130 1650 31180 1890
rect 31420 1650 31510 1890
rect 31750 1650 31840 1890
rect 32080 1650 32170 1890
rect 32410 1650 32500 1890
rect 32740 1650 32830 1890
rect 33070 1650 33160 1890
rect 33400 1650 33490 1890
rect 33730 1650 33820 1890
rect 34060 1650 34150 1890
rect 34390 1650 34480 1890
rect 34720 1650 34810 1890
rect 35050 1650 35140 1890
rect 35380 1650 35470 1890
rect 35710 1650 35800 1890
rect 36040 1650 36130 1890
rect 36370 1650 36460 1890
rect 36700 1650 36790 1890
rect 37030 1650 37120 1890
rect 37360 1650 37450 1890
rect 37690 1650 37830 1890
rect 31130 1560 37830 1650
rect 31130 1320 31180 1560
rect 31420 1320 31510 1560
rect 31750 1320 31840 1560
rect 32080 1320 32170 1560
rect 32410 1320 32500 1560
rect 32740 1320 32830 1560
rect 33070 1320 33160 1560
rect 33400 1320 33490 1560
rect 33730 1320 33820 1560
rect 34060 1320 34150 1560
rect 34390 1320 34480 1560
rect 34720 1320 34810 1560
rect 35050 1320 35140 1560
rect 35380 1320 35470 1560
rect 35710 1320 35800 1560
rect 36040 1320 36130 1560
rect 36370 1320 36460 1560
rect 36700 1320 36790 1560
rect 37030 1320 37120 1560
rect 37360 1320 37450 1560
rect 37690 1320 37830 1560
rect 31130 1180 37830 1320
rect 31130 230 37830 280
rect 31130 -10 31180 230
rect 31420 -10 31510 230
rect 31750 -10 31840 230
rect 32080 -10 32170 230
rect 32410 -10 32500 230
rect 32740 -10 32830 230
rect 33070 -10 33160 230
rect 33400 -10 33490 230
rect 33730 -10 33820 230
rect 34060 -10 34150 230
rect 34390 -10 34480 230
rect 34720 -10 34810 230
rect 35050 -10 35140 230
rect 35380 -10 35470 230
rect 35710 -10 35800 230
rect 36040 -10 36130 230
rect 36370 -10 36460 230
rect 36700 -10 36790 230
rect 37030 -10 37120 230
rect 37360 -10 37450 230
rect 37690 -10 37830 230
rect 31130 -100 37830 -10
rect 31130 -340 31180 -100
rect 31420 -340 31510 -100
rect 31750 -340 31840 -100
rect 32080 -340 32170 -100
rect 32410 -340 32500 -100
rect 32740 -340 32830 -100
rect 33070 -340 33160 -100
rect 33400 -340 33490 -100
rect 33730 -340 33820 -100
rect 34060 -340 34150 -100
rect 34390 -340 34480 -100
rect 34720 -340 34810 -100
rect 35050 -340 35140 -100
rect 35380 -340 35470 -100
rect 35710 -340 35800 -100
rect 36040 -340 36130 -100
rect 36370 -340 36460 -100
rect 36700 -340 36790 -100
rect 37030 -340 37120 -100
rect 37360 -340 37450 -100
rect 37690 -340 37830 -100
rect 31130 -430 37830 -340
rect 31130 -670 31180 -430
rect 31420 -670 31510 -430
rect 31750 -670 31840 -430
rect 32080 -670 32170 -430
rect 32410 -670 32500 -430
rect 32740 -670 32830 -430
rect 33070 -670 33160 -430
rect 33400 -670 33490 -430
rect 33730 -670 33820 -430
rect 34060 -670 34150 -430
rect 34390 -670 34480 -430
rect 34720 -670 34810 -430
rect 35050 -670 35140 -430
rect 35380 -670 35470 -430
rect 35710 -670 35800 -430
rect 36040 -670 36130 -430
rect 36370 -670 36460 -430
rect 36700 -670 36790 -430
rect 37030 -670 37120 -430
rect 37360 -670 37450 -430
rect 37690 -670 37830 -430
rect 31130 -760 37830 -670
rect 31130 -1000 31180 -760
rect 31420 -1000 31510 -760
rect 31750 -1000 31840 -760
rect 32080 -1000 32170 -760
rect 32410 -1000 32500 -760
rect 32740 -1000 32830 -760
rect 33070 -1000 33160 -760
rect 33400 -1000 33490 -760
rect 33730 -1000 33820 -760
rect 34060 -1000 34150 -760
rect 34390 -1000 34480 -760
rect 34720 -1000 34810 -760
rect 35050 -1000 35140 -760
rect 35380 -1000 35470 -760
rect 35710 -1000 35800 -760
rect 36040 -1000 36130 -760
rect 36370 -1000 36460 -760
rect 36700 -1000 36790 -760
rect 37030 -1000 37120 -760
rect 37360 -1000 37450 -760
rect 37690 -1000 37830 -760
rect 31130 -1090 37830 -1000
rect 31130 -1330 31180 -1090
rect 31420 -1330 31510 -1090
rect 31750 -1330 31840 -1090
rect 32080 -1330 32170 -1090
rect 32410 -1330 32500 -1090
rect 32740 -1330 32830 -1090
rect 33070 -1330 33160 -1090
rect 33400 -1330 33490 -1090
rect 33730 -1330 33820 -1090
rect 34060 -1330 34150 -1090
rect 34390 -1330 34480 -1090
rect 34720 -1330 34810 -1090
rect 35050 -1330 35140 -1090
rect 35380 -1330 35470 -1090
rect 35710 -1330 35800 -1090
rect 36040 -1330 36130 -1090
rect 36370 -1330 36460 -1090
rect 36700 -1330 36790 -1090
rect 37030 -1330 37120 -1090
rect 37360 -1330 37450 -1090
rect 37690 -1330 37830 -1090
rect 31130 -1420 37830 -1330
rect 31130 -1660 31180 -1420
rect 31420 -1660 31510 -1420
rect 31750 -1660 31840 -1420
rect 32080 -1660 32170 -1420
rect 32410 -1660 32500 -1420
rect 32740 -1660 32830 -1420
rect 33070 -1660 33160 -1420
rect 33400 -1660 33490 -1420
rect 33730 -1660 33820 -1420
rect 34060 -1660 34150 -1420
rect 34390 -1660 34480 -1420
rect 34720 -1660 34810 -1420
rect 35050 -1660 35140 -1420
rect 35380 -1660 35470 -1420
rect 35710 -1660 35800 -1420
rect 36040 -1660 36130 -1420
rect 36370 -1660 36460 -1420
rect 36700 -1660 36790 -1420
rect 37030 -1660 37120 -1420
rect 37360 -1660 37450 -1420
rect 37690 -1660 37830 -1420
rect 31130 -1750 37830 -1660
rect 31130 -1990 31180 -1750
rect 31420 -1990 31510 -1750
rect 31750 -1990 31840 -1750
rect 32080 -1990 32170 -1750
rect 32410 -1990 32500 -1750
rect 32740 -1990 32830 -1750
rect 33070 -1990 33160 -1750
rect 33400 -1990 33490 -1750
rect 33730 -1990 33820 -1750
rect 34060 -1990 34150 -1750
rect 34390 -1990 34480 -1750
rect 34720 -1990 34810 -1750
rect 35050 -1990 35140 -1750
rect 35380 -1990 35470 -1750
rect 35710 -1990 35800 -1750
rect 36040 -1990 36130 -1750
rect 36370 -1990 36460 -1750
rect 36700 -1990 36790 -1750
rect 37030 -1990 37120 -1750
rect 37360 -1990 37450 -1750
rect 37690 -1990 37830 -1750
rect 31130 -2080 37830 -1990
rect 31130 -2320 31180 -2080
rect 31420 -2320 31510 -2080
rect 31750 -2320 31840 -2080
rect 32080 -2320 32170 -2080
rect 32410 -2320 32500 -2080
rect 32740 -2320 32830 -2080
rect 33070 -2320 33160 -2080
rect 33400 -2320 33490 -2080
rect 33730 -2320 33820 -2080
rect 34060 -2320 34150 -2080
rect 34390 -2320 34480 -2080
rect 34720 -2320 34810 -2080
rect 35050 -2320 35140 -2080
rect 35380 -2320 35470 -2080
rect 35710 -2320 35800 -2080
rect 36040 -2320 36130 -2080
rect 36370 -2320 36460 -2080
rect 36700 -2320 36790 -2080
rect 37030 -2320 37120 -2080
rect 37360 -2320 37450 -2080
rect 37690 -2320 37830 -2080
rect 31130 -2410 37830 -2320
rect 31130 -2650 31180 -2410
rect 31420 -2650 31510 -2410
rect 31750 -2650 31840 -2410
rect 32080 -2650 32170 -2410
rect 32410 -2650 32500 -2410
rect 32740 -2650 32830 -2410
rect 33070 -2650 33160 -2410
rect 33400 -2650 33490 -2410
rect 33730 -2650 33820 -2410
rect 34060 -2650 34150 -2410
rect 34390 -2650 34480 -2410
rect 34720 -2650 34810 -2410
rect 35050 -2650 35140 -2410
rect 35380 -2650 35470 -2410
rect 35710 -2650 35800 -2410
rect 36040 -2650 36130 -2410
rect 36370 -2650 36460 -2410
rect 36700 -2650 36790 -2410
rect 37030 -2650 37120 -2410
rect 37360 -2650 37450 -2410
rect 37690 -2650 37830 -2410
rect 31130 -2740 37830 -2650
rect 31130 -2980 31180 -2740
rect 31420 -2980 31510 -2740
rect 31750 -2980 31840 -2740
rect 32080 -2980 32170 -2740
rect 32410 -2980 32500 -2740
rect 32740 -2980 32830 -2740
rect 33070 -2980 33160 -2740
rect 33400 -2980 33490 -2740
rect 33730 -2980 33820 -2740
rect 34060 -2980 34150 -2740
rect 34390 -2980 34480 -2740
rect 34720 -2980 34810 -2740
rect 35050 -2980 35140 -2740
rect 35380 -2980 35470 -2740
rect 35710 -2980 35800 -2740
rect 36040 -2980 36130 -2740
rect 36370 -2980 36460 -2740
rect 36700 -2980 36790 -2740
rect 37030 -2980 37120 -2740
rect 37360 -2980 37450 -2740
rect 37690 -2980 37830 -2740
rect 31130 -3070 37830 -2980
rect 31130 -3310 31180 -3070
rect 31420 -3310 31510 -3070
rect 31750 -3310 31840 -3070
rect 32080 -3310 32170 -3070
rect 32410 -3310 32500 -3070
rect 32740 -3310 32830 -3070
rect 33070 -3310 33160 -3070
rect 33400 -3310 33490 -3070
rect 33730 -3310 33820 -3070
rect 34060 -3310 34150 -3070
rect 34390 -3310 34480 -3070
rect 34720 -3310 34810 -3070
rect 35050 -3310 35140 -3070
rect 35380 -3310 35470 -3070
rect 35710 -3310 35800 -3070
rect 36040 -3310 36130 -3070
rect 36370 -3310 36460 -3070
rect 36700 -3310 36790 -3070
rect 37030 -3310 37120 -3070
rect 37360 -3310 37450 -3070
rect 37690 -3310 37830 -3070
rect 31130 -3400 37830 -3310
rect 31130 -3640 31180 -3400
rect 31420 -3640 31510 -3400
rect 31750 -3640 31840 -3400
rect 32080 -3640 32170 -3400
rect 32410 -3640 32500 -3400
rect 32740 -3640 32830 -3400
rect 33070 -3640 33160 -3400
rect 33400 -3640 33490 -3400
rect 33730 -3640 33820 -3400
rect 34060 -3640 34150 -3400
rect 34390 -3640 34480 -3400
rect 34720 -3640 34810 -3400
rect 35050 -3640 35140 -3400
rect 35380 -3640 35470 -3400
rect 35710 -3640 35800 -3400
rect 36040 -3640 36130 -3400
rect 36370 -3640 36460 -3400
rect 36700 -3640 36790 -3400
rect 37030 -3640 37120 -3400
rect 37360 -3640 37450 -3400
rect 37690 -3640 37830 -3400
rect 31130 -3730 37830 -3640
rect 31130 -3970 31180 -3730
rect 31420 -3970 31510 -3730
rect 31750 -3970 31840 -3730
rect 32080 -3970 32170 -3730
rect 32410 -3970 32500 -3730
rect 32740 -3970 32830 -3730
rect 33070 -3970 33160 -3730
rect 33400 -3970 33490 -3730
rect 33730 -3970 33820 -3730
rect 34060 -3970 34150 -3730
rect 34390 -3970 34480 -3730
rect 34720 -3970 34810 -3730
rect 35050 -3970 35140 -3730
rect 35380 -3970 35470 -3730
rect 35710 -3970 35800 -3730
rect 36040 -3970 36130 -3730
rect 36370 -3970 36460 -3730
rect 36700 -3970 36790 -3730
rect 37030 -3970 37120 -3730
rect 37360 -3970 37450 -3730
rect 37690 -3970 37830 -3730
rect 31130 -4060 37830 -3970
rect 31130 -4300 31180 -4060
rect 31420 -4300 31510 -4060
rect 31750 -4300 31840 -4060
rect 32080 -4300 32170 -4060
rect 32410 -4300 32500 -4060
rect 32740 -4300 32830 -4060
rect 33070 -4300 33160 -4060
rect 33400 -4300 33490 -4060
rect 33730 -4300 33820 -4060
rect 34060 -4300 34150 -4060
rect 34390 -4300 34480 -4060
rect 34720 -4300 34810 -4060
rect 35050 -4300 35140 -4060
rect 35380 -4300 35470 -4060
rect 35710 -4300 35800 -4060
rect 36040 -4300 36130 -4060
rect 36370 -4300 36460 -4060
rect 36700 -4300 36790 -4060
rect 37030 -4300 37120 -4060
rect 37360 -4300 37450 -4060
rect 37690 -4300 37830 -4060
rect 31130 -4390 37830 -4300
rect 31130 -4630 31180 -4390
rect 31420 -4630 31510 -4390
rect 31750 -4630 31840 -4390
rect 32080 -4630 32170 -4390
rect 32410 -4630 32500 -4390
rect 32740 -4630 32830 -4390
rect 33070 -4630 33160 -4390
rect 33400 -4630 33490 -4390
rect 33730 -4630 33820 -4390
rect 34060 -4630 34150 -4390
rect 34390 -4630 34480 -4390
rect 34720 -4630 34810 -4390
rect 35050 -4630 35140 -4390
rect 35380 -4630 35470 -4390
rect 35710 -4630 35800 -4390
rect 36040 -4630 36130 -4390
rect 36370 -4630 36460 -4390
rect 36700 -4630 36790 -4390
rect 37030 -4630 37120 -4390
rect 37360 -4630 37450 -4390
rect 37690 -4630 37830 -4390
rect -1320 -4840 230 -4660
rect -1320 -5080 -1180 -4840
rect -940 -5080 -850 -4840
rect -610 -5080 -520 -4840
rect -280 -5080 -190 -4840
rect 50 -5080 230 -4840
rect -1320 -5170 230 -5080
rect -1320 -5410 -1180 -5170
rect -940 -5410 -850 -5170
rect -610 -5410 -520 -5170
rect -280 -5410 -190 -5170
rect 50 -5410 230 -5170
rect -1320 -5500 230 -5410
rect -1320 -5740 -1180 -5500
rect -940 -5740 -850 -5500
rect -610 -5740 -520 -5500
rect -280 -5740 -190 -5500
rect 50 -5740 230 -5500
rect -1320 -5830 230 -5740
rect -1320 -6070 -1180 -5830
rect -940 -6070 -850 -5830
rect -610 -6070 -520 -5830
rect -280 -6070 -190 -5830
rect 50 -6070 230 -5830
rect -1320 -6210 230 -6070
rect 14550 -4840 16100 -4660
rect 14550 -5080 14730 -4840
rect 14970 -5080 15060 -4840
rect 15300 -5080 15390 -4840
rect 15630 -5080 15720 -4840
rect 15960 -5080 16100 -4840
rect 14550 -5170 16100 -5080
rect 14550 -5410 14730 -5170
rect 14970 -5410 15060 -5170
rect 15300 -5410 15390 -5170
rect 15630 -5410 15720 -5170
rect 15960 -5410 16100 -5170
rect 14550 -5500 16100 -5410
rect 14550 -5740 14730 -5500
rect 14970 -5740 15060 -5500
rect 15300 -5740 15390 -5500
rect 15630 -5740 15720 -5500
rect 15960 -5740 16100 -5500
rect 14550 -5830 16100 -5740
rect 14550 -6070 14730 -5830
rect 14970 -6070 15060 -5830
rect 15300 -6070 15390 -5830
rect 15630 -6070 15720 -5830
rect 15960 -6070 16100 -5830
rect 14550 -6210 16100 -6070
rect 31130 -4720 37830 -4630
rect 31130 -4960 31180 -4720
rect 31420 -4960 31510 -4720
rect 31750 -4960 31840 -4720
rect 32080 -4960 32170 -4720
rect 32410 -4960 32500 -4720
rect 32740 -4960 32830 -4720
rect 33070 -4960 33160 -4720
rect 33400 -4960 33490 -4720
rect 33730 -4960 33820 -4720
rect 34060 -4960 34150 -4720
rect 34390 -4960 34480 -4720
rect 34720 -4960 34810 -4720
rect 35050 -4960 35140 -4720
rect 35380 -4960 35470 -4720
rect 35710 -4960 35800 -4720
rect 36040 -4960 36130 -4720
rect 36370 -4960 36460 -4720
rect 36700 -4960 36790 -4720
rect 37030 -4960 37120 -4720
rect 37360 -4960 37450 -4720
rect 37690 -4960 37830 -4720
rect 31130 -5050 37830 -4960
rect 31130 -5290 31180 -5050
rect 31420 -5290 31510 -5050
rect 31750 -5290 31840 -5050
rect 32080 -5290 32170 -5050
rect 32410 -5290 32500 -5050
rect 32740 -5290 32830 -5050
rect 33070 -5290 33160 -5050
rect 33400 -5290 33490 -5050
rect 33730 -5290 33820 -5050
rect 34060 -5290 34150 -5050
rect 34390 -5290 34480 -5050
rect 34720 -5290 34810 -5050
rect 35050 -5290 35140 -5050
rect 35380 -5290 35470 -5050
rect 35710 -5290 35800 -5050
rect 36040 -5290 36130 -5050
rect 36370 -5290 36460 -5050
rect 36700 -5290 36790 -5050
rect 37030 -5290 37120 -5050
rect 37360 -5290 37450 -5050
rect 37690 -5290 37830 -5050
rect 31130 -5380 37830 -5290
rect 31130 -5620 31180 -5380
rect 31420 -5620 31510 -5380
rect 31750 -5620 31840 -5380
rect 32080 -5620 32170 -5380
rect 32410 -5620 32500 -5380
rect 32740 -5620 32830 -5380
rect 33070 -5620 33160 -5380
rect 33400 -5620 33490 -5380
rect 33730 -5620 33820 -5380
rect 34060 -5620 34150 -5380
rect 34390 -5620 34480 -5380
rect 34720 -5620 34810 -5380
rect 35050 -5620 35140 -5380
rect 35380 -5620 35470 -5380
rect 35710 -5620 35800 -5380
rect 36040 -5620 36130 -5380
rect 36370 -5620 36460 -5380
rect 36700 -5620 36790 -5380
rect 37030 -5620 37120 -5380
rect 37360 -5620 37450 -5380
rect 37690 -5620 37830 -5380
rect 31130 -5710 37830 -5620
rect 31130 -5950 31180 -5710
rect 31420 -5950 31510 -5710
rect 31750 -5950 31840 -5710
rect 32080 -5950 32170 -5710
rect 32410 -5950 32500 -5710
rect 32740 -5950 32830 -5710
rect 33070 -5950 33160 -5710
rect 33400 -5950 33490 -5710
rect 33730 -5950 33820 -5710
rect 34060 -5950 34150 -5710
rect 34390 -5950 34480 -5710
rect 34720 -5950 34810 -5710
rect 35050 -5950 35140 -5710
rect 35380 -5950 35470 -5710
rect 35710 -5950 35800 -5710
rect 36040 -5950 36130 -5710
rect 36370 -5950 36460 -5710
rect 36700 -5950 36790 -5710
rect 37030 -5950 37120 -5710
rect 37360 -5950 37450 -5710
rect 37690 -5950 37830 -5710
rect 31130 -6040 37830 -5950
rect 31130 -6280 31180 -6040
rect 31420 -6280 31510 -6040
rect 31750 -6280 31840 -6040
rect 32080 -6280 32170 -6040
rect 32410 -6280 32500 -6040
rect 32740 -6280 32830 -6040
rect 33070 -6280 33160 -6040
rect 33400 -6280 33490 -6040
rect 33730 -6280 33820 -6040
rect 34060 -6280 34150 -6040
rect 34390 -6280 34480 -6040
rect 34720 -6280 34810 -6040
rect 35050 -6280 35140 -6040
rect 35380 -6280 35470 -6040
rect 35710 -6280 35800 -6040
rect 36040 -6280 36130 -6040
rect 36370 -6280 36460 -6040
rect 36700 -6280 36790 -6040
rect 37030 -6280 37120 -6040
rect 37360 -6280 37450 -6040
rect 37690 -6280 37830 -6040
rect 31130 -6420 37830 -6280
<< mimcapcontact >>
rect -5200 20590 -4960 20830
rect -4870 20590 -4630 20830
rect -4540 20590 -4300 20830
rect -4210 20590 -3970 20830
rect -3880 20590 -3640 20830
rect -3550 20590 -3310 20830
rect -3220 20590 -2980 20830
rect -2890 20590 -2650 20830
rect -2560 20590 -2320 20830
rect -2230 20590 -1990 20830
rect -1900 20590 -1660 20830
rect -1570 20590 -1330 20830
rect -1240 20590 -1000 20830
rect -910 20590 -670 20830
rect -580 20590 -340 20830
rect -250 20590 -10 20830
rect 80 20590 320 20830
rect 410 20590 650 20830
rect 740 20590 980 20830
rect 1070 20590 1310 20830
rect 1400 20590 1640 20830
rect 1730 20590 1970 20830
rect 2060 20590 2300 20830
rect 2390 20590 2630 20830
rect 2720 20590 2960 20830
rect 3050 20590 3290 20830
rect 3380 20590 3620 20830
rect 3710 20590 3950 20830
rect 4040 20590 4280 20830
rect 4370 20590 4610 20830
rect 4700 20590 4940 20830
rect 5030 20590 5270 20830
rect 5360 20590 5600 20830
rect 5690 20590 5930 20830
rect 6020 20590 6260 20830
rect 6350 20590 6590 20830
rect -5200 20260 -4960 20500
rect -4870 20260 -4630 20500
rect -4540 20260 -4300 20500
rect -4210 20260 -3970 20500
rect -3880 20260 -3640 20500
rect -3550 20260 -3310 20500
rect -3220 20260 -2980 20500
rect -2890 20260 -2650 20500
rect -2560 20260 -2320 20500
rect -2230 20260 -1990 20500
rect -1900 20260 -1660 20500
rect -1570 20260 -1330 20500
rect -1240 20260 -1000 20500
rect -910 20260 -670 20500
rect -580 20260 -340 20500
rect -250 20260 -10 20500
rect 80 20260 320 20500
rect 410 20260 650 20500
rect 740 20260 980 20500
rect 1070 20260 1310 20500
rect 1400 20260 1640 20500
rect 1730 20260 1970 20500
rect 2060 20260 2300 20500
rect 2390 20260 2630 20500
rect 2720 20260 2960 20500
rect 3050 20260 3290 20500
rect 3380 20260 3620 20500
rect 3710 20260 3950 20500
rect 4040 20260 4280 20500
rect 4370 20260 4610 20500
rect 4700 20260 4940 20500
rect 5030 20260 5270 20500
rect 5360 20260 5600 20500
rect 5690 20260 5930 20500
rect 6020 20260 6260 20500
rect 6350 20260 6590 20500
rect -5200 19930 -4960 20170
rect -4870 19930 -4630 20170
rect -4540 19930 -4300 20170
rect -4210 19930 -3970 20170
rect -3880 19930 -3640 20170
rect -3550 19930 -3310 20170
rect -3220 19930 -2980 20170
rect -2890 19930 -2650 20170
rect -2560 19930 -2320 20170
rect -2230 19930 -1990 20170
rect -1900 19930 -1660 20170
rect -1570 19930 -1330 20170
rect -1240 19930 -1000 20170
rect -910 19930 -670 20170
rect -580 19930 -340 20170
rect -250 19930 -10 20170
rect 80 19930 320 20170
rect 410 19930 650 20170
rect 740 19930 980 20170
rect 1070 19930 1310 20170
rect 1400 19930 1640 20170
rect 1730 19930 1970 20170
rect 2060 19930 2300 20170
rect 2390 19930 2630 20170
rect 2720 19930 2960 20170
rect 3050 19930 3290 20170
rect 3380 19930 3620 20170
rect 3710 19930 3950 20170
rect 4040 19930 4280 20170
rect 4370 19930 4610 20170
rect 4700 19930 4940 20170
rect 5030 19930 5270 20170
rect 5360 19930 5600 20170
rect 5690 19930 5930 20170
rect 6020 19930 6260 20170
rect 6350 19930 6590 20170
rect -5200 19600 -4960 19840
rect -4870 19600 -4630 19840
rect -4540 19600 -4300 19840
rect -4210 19600 -3970 19840
rect -3880 19600 -3640 19840
rect -3550 19600 -3310 19840
rect -3220 19600 -2980 19840
rect -2890 19600 -2650 19840
rect -2560 19600 -2320 19840
rect -2230 19600 -1990 19840
rect -1900 19600 -1660 19840
rect -1570 19600 -1330 19840
rect -1240 19600 -1000 19840
rect -910 19600 -670 19840
rect -580 19600 -340 19840
rect -250 19600 -10 19840
rect 80 19600 320 19840
rect 410 19600 650 19840
rect 740 19600 980 19840
rect 1070 19600 1310 19840
rect 1400 19600 1640 19840
rect 1730 19600 1970 19840
rect 2060 19600 2300 19840
rect 2390 19600 2630 19840
rect 2720 19600 2960 19840
rect 3050 19600 3290 19840
rect 3380 19600 3620 19840
rect 3710 19600 3950 19840
rect 4040 19600 4280 19840
rect 4370 19600 4610 19840
rect 4700 19600 4940 19840
rect 5030 19600 5270 19840
rect 5360 19600 5600 19840
rect 5690 19600 5930 19840
rect 6020 19600 6260 19840
rect 6350 19600 6590 19840
rect -5200 19270 -4960 19510
rect -4870 19270 -4630 19510
rect -4540 19270 -4300 19510
rect -4210 19270 -3970 19510
rect -3880 19270 -3640 19510
rect -3550 19270 -3310 19510
rect -3220 19270 -2980 19510
rect -2890 19270 -2650 19510
rect -2560 19270 -2320 19510
rect -2230 19270 -1990 19510
rect -1900 19270 -1660 19510
rect -1570 19270 -1330 19510
rect -1240 19270 -1000 19510
rect -910 19270 -670 19510
rect -580 19270 -340 19510
rect -250 19270 -10 19510
rect 80 19270 320 19510
rect 410 19270 650 19510
rect 740 19270 980 19510
rect 1070 19270 1310 19510
rect 1400 19270 1640 19510
rect 1730 19270 1970 19510
rect 2060 19270 2300 19510
rect 2390 19270 2630 19510
rect 2720 19270 2960 19510
rect 3050 19270 3290 19510
rect 3380 19270 3620 19510
rect 3710 19270 3950 19510
rect 4040 19270 4280 19510
rect 4370 19270 4610 19510
rect 4700 19270 4940 19510
rect 5030 19270 5270 19510
rect 5360 19270 5600 19510
rect 5690 19270 5930 19510
rect 6020 19270 6260 19510
rect 6350 19270 6590 19510
rect -5200 18940 -4960 19180
rect -4870 18940 -4630 19180
rect -4540 18940 -4300 19180
rect -4210 18940 -3970 19180
rect -3880 18940 -3640 19180
rect -3550 18940 -3310 19180
rect -3220 18940 -2980 19180
rect -2890 18940 -2650 19180
rect -2560 18940 -2320 19180
rect -2230 18940 -1990 19180
rect -1900 18940 -1660 19180
rect -1570 18940 -1330 19180
rect -1240 18940 -1000 19180
rect -910 18940 -670 19180
rect -580 18940 -340 19180
rect -250 18940 -10 19180
rect 80 18940 320 19180
rect 410 18940 650 19180
rect 740 18940 980 19180
rect 1070 18940 1310 19180
rect 1400 18940 1640 19180
rect 1730 18940 1970 19180
rect 2060 18940 2300 19180
rect 2390 18940 2630 19180
rect 2720 18940 2960 19180
rect 3050 18940 3290 19180
rect 3380 18940 3620 19180
rect 3710 18940 3950 19180
rect 4040 18940 4280 19180
rect 4370 18940 4610 19180
rect 4700 18940 4940 19180
rect 5030 18940 5270 19180
rect 5360 18940 5600 19180
rect 5690 18940 5930 19180
rect 6020 18940 6260 19180
rect 6350 18940 6590 19180
rect -5200 18610 -4960 18850
rect -4870 18610 -4630 18850
rect -4540 18610 -4300 18850
rect -4210 18610 -3970 18850
rect -3880 18610 -3640 18850
rect -3550 18610 -3310 18850
rect -3220 18610 -2980 18850
rect -2890 18610 -2650 18850
rect -2560 18610 -2320 18850
rect -2230 18610 -1990 18850
rect -1900 18610 -1660 18850
rect -1570 18610 -1330 18850
rect -1240 18610 -1000 18850
rect -910 18610 -670 18850
rect -580 18610 -340 18850
rect -250 18610 -10 18850
rect 80 18610 320 18850
rect 410 18610 650 18850
rect 740 18610 980 18850
rect 1070 18610 1310 18850
rect 1400 18610 1640 18850
rect 1730 18610 1970 18850
rect 2060 18610 2300 18850
rect 2390 18610 2630 18850
rect 2720 18610 2960 18850
rect 3050 18610 3290 18850
rect 3380 18610 3620 18850
rect 3710 18610 3950 18850
rect 4040 18610 4280 18850
rect 4370 18610 4610 18850
rect 4700 18610 4940 18850
rect 5030 18610 5270 18850
rect 5360 18610 5600 18850
rect 5690 18610 5930 18850
rect 6020 18610 6260 18850
rect 6350 18610 6590 18850
rect -5200 18280 -4960 18520
rect -4870 18280 -4630 18520
rect -4540 18280 -4300 18520
rect -4210 18280 -3970 18520
rect -3880 18280 -3640 18520
rect -3550 18280 -3310 18520
rect -3220 18280 -2980 18520
rect -2890 18280 -2650 18520
rect -2560 18280 -2320 18520
rect -2230 18280 -1990 18520
rect -1900 18280 -1660 18520
rect -1570 18280 -1330 18520
rect -1240 18280 -1000 18520
rect -910 18280 -670 18520
rect -580 18280 -340 18520
rect -250 18280 -10 18520
rect 80 18280 320 18520
rect 410 18280 650 18520
rect 740 18280 980 18520
rect 1070 18280 1310 18520
rect 1400 18280 1640 18520
rect 1730 18280 1970 18520
rect 2060 18280 2300 18520
rect 2390 18280 2630 18520
rect 2720 18280 2960 18520
rect 3050 18280 3290 18520
rect 3380 18280 3620 18520
rect 3710 18280 3950 18520
rect 4040 18280 4280 18520
rect 4370 18280 4610 18520
rect 4700 18280 4940 18520
rect 5030 18280 5270 18520
rect 5360 18280 5600 18520
rect 5690 18280 5930 18520
rect 6020 18280 6260 18520
rect 6350 18280 6590 18520
rect -5200 17950 -4960 18190
rect -4870 17950 -4630 18190
rect -4540 17950 -4300 18190
rect -4210 17950 -3970 18190
rect -3880 17950 -3640 18190
rect -3550 17950 -3310 18190
rect -3220 17950 -2980 18190
rect -2890 17950 -2650 18190
rect -2560 17950 -2320 18190
rect -2230 17950 -1990 18190
rect -1900 17950 -1660 18190
rect -1570 17950 -1330 18190
rect -1240 17950 -1000 18190
rect -910 17950 -670 18190
rect -580 17950 -340 18190
rect -250 17950 -10 18190
rect 80 17950 320 18190
rect 410 17950 650 18190
rect 740 17950 980 18190
rect 1070 17950 1310 18190
rect 1400 17950 1640 18190
rect 1730 17950 1970 18190
rect 2060 17950 2300 18190
rect 2390 17950 2630 18190
rect 2720 17950 2960 18190
rect 3050 17950 3290 18190
rect 3380 17950 3620 18190
rect 3710 17950 3950 18190
rect 4040 17950 4280 18190
rect 4370 17950 4610 18190
rect 4700 17950 4940 18190
rect 5030 17950 5270 18190
rect 5360 17950 5600 18190
rect 5690 17950 5930 18190
rect 6020 17950 6260 18190
rect 6350 17950 6590 18190
rect -5200 17620 -4960 17860
rect -4870 17620 -4630 17860
rect -4540 17620 -4300 17860
rect -4210 17620 -3970 17860
rect -3880 17620 -3640 17860
rect -3550 17620 -3310 17860
rect -3220 17620 -2980 17860
rect -2890 17620 -2650 17860
rect -2560 17620 -2320 17860
rect -2230 17620 -1990 17860
rect -1900 17620 -1660 17860
rect -1570 17620 -1330 17860
rect -1240 17620 -1000 17860
rect -910 17620 -670 17860
rect -580 17620 -340 17860
rect -250 17620 -10 17860
rect 80 17620 320 17860
rect 410 17620 650 17860
rect 740 17620 980 17860
rect 1070 17620 1310 17860
rect 1400 17620 1640 17860
rect 1730 17620 1970 17860
rect 2060 17620 2300 17860
rect 2390 17620 2630 17860
rect 2720 17620 2960 17860
rect 3050 17620 3290 17860
rect 3380 17620 3620 17860
rect 3710 17620 3950 17860
rect 4040 17620 4280 17860
rect 4370 17620 4610 17860
rect 4700 17620 4940 17860
rect 5030 17620 5270 17860
rect 5360 17620 5600 17860
rect 5690 17620 5930 17860
rect 6020 17620 6260 17860
rect 6350 17620 6590 17860
rect -5200 17290 -4960 17530
rect -4870 17290 -4630 17530
rect -4540 17290 -4300 17530
rect -4210 17290 -3970 17530
rect -3880 17290 -3640 17530
rect -3550 17290 -3310 17530
rect -3220 17290 -2980 17530
rect -2890 17290 -2650 17530
rect -2560 17290 -2320 17530
rect -2230 17290 -1990 17530
rect -1900 17290 -1660 17530
rect -1570 17290 -1330 17530
rect -1240 17290 -1000 17530
rect -910 17290 -670 17530
rect -580 17290 -340 17530
rect -250 17290 -10 17530
rect 80 17290 320 17530
rect 410 17290 650 17530
rect 740 17290 980 17530
rect 1070 17290 1310 17530
rect 1400 17290 1640 17530
rect 1730 17290 1970 17530
rect 2060 17290 2300 17530
rect 2390 17290 2630 17530
rect 2720 17290 2960 17530
rect 3050 17290 3290 17530
rect 3380 17290 3620 17530
rect 3710 17290 3950 17530
rect 4040 17290 4280 17530
rect 4370 17290 4610 17530
rect 4700 17290 4940 17530
rect 5030 17290 5270 17530
rect 5360 17290 5600 17530
rect 5690 17290 5930 17530
rect 6020 17290 6260 17530
rect 6350 17290 6590 17530
rect -5200 16960 -4960 17200
rect -4870 16960 -4630 17200
rect -4540 16960 -4300 17200
rect -4210 16960 -3970 17200
rect -3880 16960 -3640 17200
rect -3550 16960 -3310 17200
rect -3220 16960 -2980 17200
rect -2890 16960 -2650 17200
rect -2560 16960 -2320 17200
rect -2230 16960 -1990 17200
rect -1900 16960 -1660 17200
rect -1570 16960 -1330 17200
rect -1240 16960 -1000 17200
rect -910 16960 -670 17200
rect -580 16960 -340 17200
rect -250 16960 -10 17200
rect 80 16960 320 17200
rect 410 16960 650 17200
rect 740 16960 980 17200
rect 1070 16960 1310 17200
rect 1400 16960 1640 17200
rect 1730 16960 1970 17200
rect 2060 16960 2300 17200
rect 2390 16960 2630 17200
rect 2720 16960 2960 17200
rect 3050 16960 3290 17200
rect 3380 16960 3620 17200
rect 3710 16960 3950 17200
rect 4040 16960 4280 17200
rect 4370 16960 4610 17200
rect 4700 16960 4940 17200
rect 5030 16960 5270 17200
rect 5360 16960 5600 17200
rect 5690 16960 5930 17200
rect 6020 16960 6260 17200
rect 6350 16960 6590 17200
rect -5200 16630 -4960 16870
rect -4870 16630 -4630 16870
rect -4540 16630 -4300 16870
rect -4210 16630 -3970 16870
rect -3880 16630 -3640 16870
rect -3550 16630 -3310 16870
rect -3220 16630 -2980 16870
rect -2890 16630 -2650 16870
rect -2560 16630 -2320 16870
rect -2230 16630 -1990 16870
rect -1900 16630 -1660 16870
rect -1570 16630 -1330 16870
rect -1240 16630 -1000 16870
rect -910 16630 -670 16870
rect -580 16630 -340 16870
rect -250 16630 -10 16870
rect 80 16630 320 16870
rect 410 16630 650 16870
rect 740 16630 980 16870
rect 1070 16630 1310 16870
rect 1400 16630 1640 16870
rect 1730 16630 1970 16870
rect 2060 16630 2300 16870
rect 2390 16630 2630 16870
rect 2720 16630 2960 16870
rect 3050 16630 3290 16870
rect 3380 16630 3620 16870
rect 3710 16630 3950 16870
rect 4040 16630 4280 16870
rect 4370 16630 4610 16870
rect 4700 16630 4940 16870
rect 5030 16630 5270 16870
rect 5360 16630 5600 16870
rect 5690 16630 5930 16870
rect 6020 16630 6260 16870
rect 6350 16630 6590 16870
rect -5200 16300 -4960 16540
rect -4870 16300 -4630 16540
rect -4540 16300 -4300 16540
rect -4210 16300 -3970 16540
rect -3880 16300 -3640 16540
rect -3550 16300 -3310 16540
rect -3220 16300 -2980 16540
rect -2890 16300 -2650 16540
rect -2560 16300 -2320 16540
rect -2230 16300 -1990 16540
rect -1900 16300 -1660 16540
rect -1570 16300 -1330 16540
rect -1240 16300 -1000 16540
rect -910 16300 -670 16540
rect -580 16300 -340 16540
rect -250 16300 -10 16540
rect 80 16300 320 16540
rect 410 16300 650 16540
rect 740 16300 980 16540
rect 1070 16300 1310 16540
rect 1400 16300 1640 16540
rect 1730 16300 1970 16540
rect 2060 16300 2300 16540
rect 2390 16300 2630 16540
rect 2720 16300 2960 16540
rect 3050 16300 3290 16540
rect 3380 16300 3620 16540
rect 3710 16300 3950 16540
rect 4040 16300 4280 16540
rect 4370 16300 4610 16540
rect 4700 16300 4940 16540
rect 5030 16300 5270 16540
rect 5360 16300 5600 16540
rect 5690 16300 5930 16540
rect 6020 16300 6260 16540
rect 6350 16300 6590 16540
rect -5200 15970 -4960 16210
rect -4870 15970 -4630 16210
rect -4540 15970 -4300 16210
rect -4210 15970 -3970 16210
rect -3880 15970 -3640 16210
rect -3550 15970 -3310 16210
rect -3220 15970 -2980 16210
rect -2890 15970 -2650 16210
rect -2560 15970 -2320 16210
rect -2230 15970 -1990 16210
rect -1900 15970 -1660 16210
rect -1570 15970 -1330 16210
rect -1240 15970 -1000 16210
rect -910 15970 -670 16210
rect -580 15970 -340 16210
rect -250 15970 -10 16210
rect 80 15970 320 16210
rect 410 15970 650 16210
rect 740 15970 980 16210
rect 1070 15970 1310 16210
rect 1400 15970 1640 16210
rect 1730 15970 1970 16210
rect 2060 15970 2300 16210
rect 2390 15970 2630 16210
rect 2720 15970 2960 16210
rect 3050 15970 3290 16210
rect 3380 15970 3620 16210
rect 3710 15970 3950 16210
rect 4040 15970 4280 16210
rect 4370 15970 4610 16210
rect 4700 15970 4940 16210
rect 5030 15970 5270 16210
rect 5360 15970 5600 16210
rect 5690 15970 5930 16210
rect 6020 15970 6260 16210
rect 6350 15970 6590 16210
rect -5200 15640 -4960 15880
rect -4870 15640 -4630 15880
rect -4540 15640 -4300 15880
rect -4210 15640 -3970 15880
rect -3880 15640 -3640 15880
rect -3550 15640 -3310 15880
rect -3220 15640 -2980 15880
rect -2890 15640 -2650 15880
rect -2560 15640 -2320 15880
rect -2230 15640 -1990 15880
rect -1900 15640 -1660 15880
rect -1570 15640 -1330 15880
rect -1240 15640 -1000 15880
rect -910 15640 -670 15880
rect -580 15640 -340 15880
rect -250 15640 -10 15880
rect 80 15640 320 15880
rect 410 15640 650 15880
rect 740 15640 980 15880
rect 1070 15640 1310 15880
rect 1400 15640 1640 15880
rect 1730 15640 1970 15880
rect 2060 15640 2300 15880
rect 2390 15640 2630 15880
rect 2720 15640 2960 15880
rect 3050 15640 3290 15880
rect 3380 15640 3620 15880
rect 3710 15640 3950 15880
rect 4040 15640 4280 15880
rect 4370 15640 4610 15880
rect 4700 15640 4940 15880
rect 5030 15640 5270 15880
rect 5360 15640 5600 15880
rect 5690 15640 5930 15880
rect 6020 15640 6260 15880
rect 6350 15640 6590 15880
rect -5200 15310 -4960 15550
rect -4870 15310 -4630 15550
rect -4540 15310 -4300 15550
rect -4210 15310 -3970 15550
rect -3880 15310 -3640 15550
rect -3550 15310 -3310 15550
rect -3220 15310 -2980 15550
rect -2890 15310 -2650 15550
rect -2560 15310 -2320 15550
rect -2230 15310 -1990 15550
rect -1900 15310 -1660 15550
rect -1570 15310 -1330 15550
rect -1240 15310 -1000 15550
rect -910 15310 -670 15550
rect -580 15310 -340 15550
rect -250 15310 -10 15550
rect 80 15310 320 15550
rect 410 15310 650 15550
rect 740 15310 980 15550
rect 1070 15310 1310 15550
rect 1400 15310 1640 15550
rect 1730 15310 1970 15550
rect 2060 15310 2300 15550
rect 2390 15310 2630 15550
rect 2720 15310 2960 15550
rect 3050 15310 3290 15550
rect 3380 15310 3620 15550
rect 3710 15310 3950 15550
rect 4040 15310 4280 15550
rect 4370 15310 4610 15550
rect 4700 15310 4940 15550
rect 5030 15310 5270 15550
rect 5360 15310 5600 15550
rect 5690 15310 5930 15550
rect 6020 15310 6260 15550
rect 6350 15310 6590 15550
rect -5200 14980 -4960 15220
rect -4870 14980 -4630 15220
rect -4540 14980 -4300 15220
rect -4210 14980 -3970 15220
rect -3880 14980 -3640 15220
rect -3550 14980 -3310 15220
rect -3220 14980 -2980 15220
rect -2890 14980 -2650 15220
rect -2560 14980 -2320 15220
rect -2230 14980 -1990 15220
rect -1900 14980 -1660 15220
rect -1570 14980 -1330 15220
rect -1240 14980 -1000 15220
rect -910 14980 -670 15220
rect -580 14980 -340 15220
rect -250 14980 -10 15220
rect 80 14980 320 15220
rect 410 14980 650 15220
rect 740 14980 980 15220
rect 1070 14980 1310 15220
rect 1400 14980 1640 15220
rect 1730 14980 1970 15220
rect 2060 14980 2300 15220
rect 2390 14980 2630 15220
rect 2720 14980 2960 15220
rect 3050 14980 3290 15220
rect 3380 14980 3620 15220
rect 3710 14980 3950 15220
rect 4040 14980 4280 15220
rect 4370 14980 4610 15220
rect 4700 14980 4940 15220
rect 5030 14980 5270 15220
rect 5360 14980 5600 15220
rect 5690 14980 5930 15220
rect 6020 14980 6260 15220
rect 6350 14980 6590 15220
rect -5200 14650 -4960 14890
rect -4870 14650 -4630 14890
rect -4540 14650 -4300 14890
rect -4210 14650 -3970 14890
rect -3880 14650 -3640 14890
rect -3550 14650 -3310 14890
rect -3220 14650 -2980 14890
rect -2890 14650 -2650 14890
rect -2560 14650 -2320 14890
rect -2230 14650 -1990 14890
rect -1900 14650 -1660 14890
rect -1570 14650 -1330 14890
rect -1240 14650 -1000 14890
rect -910 14650 -670 14890
rect -580 14650 -340 14890
rect -250 14650 -10 14890
rect 80 14650 320 14890
rect 410 14650 650 14890
rect 740 14650 980 14890
rect 1070 14650 1310 14890
rect 1400 14650 1640 14890
rect 1730 14650 1970 14890
rect 2060 14650 2300 14890
rect 2390 14650 2630 14890
rect 2720 14650 2960 14890
rect 3050 14650 3290 14890
rect 3380 14650 3620 14890
rect 3710 14650 3950 14890
rect 4040 14650 4280 14890
rect 4370 14650 4610 14890
rect 4700 14650 4940 14890
rect 5030 14650 5270 14890
rect 5360 14650 5600 14890
rect 5690 14650 5930 14890
rect 6020 14650 6260 14890
rect 6350 14650 6590 14890
rect -5200 14320 -4960 14560
rect -4870 14320 -4630 14560
rect -4540 14320 -4300 14560
rect -4210 14320 -3970 14560
rect -3880 14320 -3640 14560
rect -3550 14320 -3310 14560
rect -3220 14320 -2980 14560
rect -2890 14320 -2650 14560
rect -2560 14320 -2320 14560
rect -2230 14320 -1990 14560
rect -1900 14320 -1660 14560
rect -1570 14320 -1330 14560
rect -1240 14320 -1000 14560
rect -910 14320 -670 14560
rect -580 14320 -340 14560
rect -250 14320 -10 14560
rect 80 14320 320 14560
rect 410 14320 650 14560
rect 740 14320 980 14560
rect 1070 14320 1310 14560
rect 1400 14320 1640 14560
rect 1730 14320 1970 14560
rect 2060 14320 2300 14560
rect 2390 14320 2630 14560
rect 2720 14320 2960 14560
rect 3050 14320 3290 14560
rect 3380 14320 3620 14560
rect 3710 14320 3950 14560
rect 4040 14320 4280 14560
rect 4370 14320 4610 14560
rect 4700 14320 4940 14560
rect 5030 14320 5270 14560
rect 5360 14320 5600 14560
rect 5690 14320 5930 14560
rect 6020 14320 6260 14560
rect 6350 14320 6590 14560
rect -5200 13990 -4960 14230
rect -4870 13990 -4630 14230
rect -4540 13990 -4300 14230
rect -4210 13990 -3970 14230
rect -3880 13990 -3640 14230
rect -3550 13990 -3310 14230
rect -3220 13990 -2980 14230
rect -2890 13990 -2650 14230
rect -2560 13990 -2320 14230
rect -2230 13990 -1990 14230
rect -1900 13990 -1660 14230
rect -1570 13990 -1330 14230
rect -1240 13990 -1000 14230
rect -910 13990 -670 14230
rect -580 13990 -340 14230
rect -250 13990 -10 14230
rect 80 13990 320 14230
rect 410 13990 650 14230
rect 740 13990 980 14230
rect 1070 13990 1310 14230
rect 1400 13990 1640 14230
rect 1730 13990 1970 14230
rect 2060 13990 2300 14230
rect 2390 13990 2630 14230
rect 2720 13990 2960 14230
rect 3050 13990 3290 14230
rect 3380 13990 3620 14230
rect 3710 13990 3950 14230
rect 4040 13990 4280 14230
rect 4370 13990 4610 14230
rect 4700 13990 4940 14230
rect 5030 13990 5270 14230
rect 5360 13990 5600 14230
rect 5690 13990 5930 14230
rect 6020 13990 6260 14230
rect 6350 13990 6590 14230
rect -5200 13660 -4960 13900
rect -4870 13660 -4630 13900
rect -4540 13660 -4300 13900
rect -4210 13660 -3970 13900
rect -3880 13660 -3640 13900
rect -3550 13660 -3310 13900
rect -3220 13660 -2980 13900
rect -2890 13660 -2650 13900
rect -2560 13660 -2320 13900
rect -2230 13660 -1990 13900
rect -1900 13660 -1660 13900
rect -1570 13660 -1330 13900
rect -1240 13660 -1000 13900
rect -910 13660 -670 13900
rect -580 13660 -340 13900
rect -250 13660 -10 13900
rect 80 13660 320 13900
rect 410 13660 650 13900
rect 740 13660 980 13900
rect 1070 13660 1310 13900
rect 1400 13660 1640 13900
rect 1730 13660 1970 13900
rect 2060 13660 2300 13900
rect 2390 13660 2630 13900
rect 2720 13660 2960 13900
rect 3050 13660 3290 13900
rect 3380 13660 3620 13900
rect 3710 13660 3950 13900
rect 4040 13660 4280 13900
rect 4370 13660 4610 13900
rect 4700 13660 4940 13900
rect 5030 13660 5270 13900
rect 5360 13660 5600 13900
rect 5690 13660 5930 13900
rect 6020 13660 6260 13900
rect 6350 13660 6590 13900
rect -5200 13330 -4960 13570
rect -4870 13330 -4630 13570
rect -4540 13330 -4300 13570
rect -4210 13330 -3970 13570
rect -3880 13330 -3640 13570
rect -3550 13330 -3310 13570
rect -3220 13330 -2980 13570
rect -2890 13330 -2650 13570
rect -2560 13330 -2320 13570
rect -2230 13330 -1990 13570
rect -1900 13330 -1660 13570
rect -1570 13330 -1330 13570
rect -1240 13330 -1000 13570
rect -910 13330 -670 13570
rect -580 13330 -340 13570
rect -250 13330 -10 13570
rect 80 13330 320 13570
rect 410 13330 650 13570
rect 740 13330 980 13570
rect 1070 13330 1310 13570
rect 1400 13330 1640 13570
rect 1730 13330 1970 13570
rect 2060 13330 2300 13570
rect 2390 13330 2630 13570
rect 2720 13330 2960 13570
rect 3050 13330 3290 13570
rect 3380 13330 3620 13570
rect 3710 13330 3950 13570
rect 4040 13330 4280 13570
rect 4370 13330 4610 13570
rect 4700 13330 4940 13570
rect 5030 13330 5270 13570
rect 5360 13330 5600 13570
rect 5690 13330 5930 13570
rect 6020 13330 6260 13570
rect 6350 13330 6590 13570
rect -5200 13000 -4960 13240
rect -4870 13000 -4630 13240
rect -4540 13000 -4300 13240
rect -4210 13000 -3970 13240
rect -3880 13000 -3640 13240
rect -3550 13000 -3310 13240
rect -3220 13000 -2980 13240
rect -2890 13000 -2650 13240
rect -2560 13000 -2320 13240
rect -2230 13000 -1990 13240
rect -1900 13000 -1660 13240
rect -1570 13000 -1330 13240
rect -1240 13000 -1000 13240
rect -910 13000 -670 13240
rect -580 13000 -340 13240
rect -250 13000 -10 13240
rect 80 13000 320 13240
rect 410 13000 650 13240
rect 740 13000 980 13240
rect 1070 13000 1310 13240
rect 1400 13000 1640 13240
rect 1730 13000 1970 13240
rect 2060 13000 2300 13240
rect 2390 13000 2630 13240
rect 2720 13000 2960 13240
rect 3050 13000 3290 13240
rect 3380 13000 3620 13240
rect 3710 13000 3950 13240
rect 4040 13000 4280 13240
rect 4370 13000 4610 13240
rect 4700 13000 4940 13240
rect 5030 13000 5270 13240
rect 5360 13000 5600 13240
rect 5690 13000 5930 13240
rect 6020 13000 6260 13240
rect 6350 13000 6590 13240
rect -5200 12670 -4960 12910
rect -4870 12670 -4630 12910
rect -4540 12670 -4300 12910
rect -4210 12670 -3970 12910
rect -3880 12670 -3640 12910
rect -3550 12670 -3310 12910
rect -3220 12670 -2980 12910
rect -2890 12670 -2650 12910
rect -2560 12670 -2320 12910
rect -2230 12670 -1990 12910
rect -1900 12670 -1660 12910
rect -1570 12670 -1330 12910
rect -1240 12670 -1000 12910
rect -910 12670 -670 12910
rect -580 12670 -340 12910
rect -250 12670 -10 12910
rect 80 12670 320 12910
rect 410 12670 650 12910
rect 740 12670 980 12910
rect 1070 12670 1310 12910
rect 1400 12670 1640 12910
rect 1730 12670 1970 12910
rect 2060 12670 2300 12910
rect 2390 12670 2630 12910
rect 2720 12670 2960 12910
rect 3050 12670 3290 12910
rect 3380 12670 3620 12910
rect 3710 12670 3950 12910
rect 4040 12670 4280 12910
rect 4370 12670 4610 12910
rect 4700 12670 4940 12910
rect 5030 12670 5270 12910
rect 5360 12670 5600 12910
rect 5690 12670 5930 12910
rect 6020 12670 6260 12910
rect 6350 12670 6590 12910
rect -5200 12340 -4960 12580
rect -4870 12340 -4630 12580
rect -4540 12340 -4300 12580
rect -4210 12340 -3970 12580
rect -3880 12340 -3640 12580
rect -3550 12340 -3310 12580
rect -3220 12340 -2980 12580
rect -2890 12340 -2650 12580
rect -2560 12340 -2320 12580
rect -2230 12340 -1990 12580
rect -1900 12340 -1660 12580
rect -1570 12340 -1330 12580
rect -1240 12340 -1000 12580
rect -910 12340 -670 12580
rect -580 12340 -340 12580
rect -250 12340 -10 12580
rect 80 12340 320 12580
rect 410 12340 650 12580
rect 740 12340 980 12580
rect 1070 12340 1310 12580
rect 1400 12340 1640 12580
rect 1730 12340 1970 12580
rect 2060 12340 2300 12580
rect 2390 12340 2630 12580
rect 2720 12340 2960 12580
rect 3050 12340 3290 12580
rect 3380 12340 3620 12580
rect 3710 12340 3950 12580
rect 4040 12340 4280 12580
rect 4370 12340 4610 12580
rect 4700 12340 4940 12580
rect 5030 12340 5270 12580
rect 5360 12340 5600 12580
rect 5690 12340 5930 12580
rect 6020 12340 6260 12580
rect 6350 12340 6590 12580
rect -5200 12010 -4960 12250
rect -4870 12010 -4630 12250
rect -4540 12010 -4300 12250
rect -4210 12010 -3970 12250
rect -3880 12010 -3640 12250
rect -3550 12010 -3310 12250
rect -3220 12010 -2980 12250
rect -2890 12010 -2650 12250
rect -2560 12010 -2320 12250
rect -2230 12010 -1990 12250
rect -1900 12010 -1660 12250
rect -1570 12010 -1330 12250
rect -1240 12010 -1000 12250
rect -910 12010 -670 12250
rect -580 12010 -340 12250
rect -250 12010 -10 12250
rect 80 12010 320 12250
rect 410 12010 650 12250
rect 740 12010 980 12250
rect 1070 12010 1310 12250
rect 1400 12010 1640 12250
rect 1730 12010 1970 12250
rect 2060 12010 2300 12250
rect 2390 12010 2630 12250
rect 2720 12010 2960 12250
rect 3050 12010 3290 12250
rect 3380 12010 3620 12250
rect 3710 12010 3950 12250
rect 4040 12010 4280 12250
rect 4370 12010 4610 12250
rect 4700 12010 4940 12250
rect 5030 12010 5270 12250
rect 5360 12010 5600 12250
rect 5690 12010 5930 12250
rect 6020 12010 6260 12250
rect 6350 12010 6590 12250
rect -5200 11680 -4960 11920
rect -4870 11680 -4630 11920
rect -4540 11680 -4300 11920
rect -4210 11680 -3970 11920
rect -3880 11680 -3640 11920
rect -3550 11680 -3310 11920
rect -3220 11680 -2980 11920
rect -2890 11680 -2650 11920
rect -2560 11680 -2320 11920
rect -2230 11680 -1990 11920
rect -1900 11680 -1660 11920
rect -1570 11680 -1330 11920
rect -1240 11680 -1000 11920
rect -910 11680 -670 11920
rect -580 11680 -340 11920
rect -250 11680 -10 11920
rect 80 11680 320 11920
rect 410 11680 650 11920
rect 740 11680 980 11920
rect 1070 11680 1310 11920
rect 1400 11680 1640 11920
rect 1730 11680 1970 11920
rect 2060 11680 2300 11920
rect 2390 11680 2630 11920
rect 2720 11680 2960 11920
rect 3050 11680 3290 11920
rect 3380 11680 3620 11920
rect 3710 11680 3950 11920
rect 4040 11680 4280 11920
rect 4370 11680 4610 11920
rect 4700 11680 4940 11920
rect 5030 11680 5270 11920
rect 5360 11680 5600 11920
rect 5690 11680 5930 11920
rect 6020 11680 6260 11920
rect 6350 11680 6590 11920
rect -5200 11350 -4960 11590
rect -4870 11350 -4630 11590
rect -4540 11350 -4300 11590
rect -4210 11350 -3970 11590
rect -3880 11350 -3640 11590
rect -3550 11350 -3310 11590
rect -3220 11350 -2980 11590
rect -2890 11350 -2650 11590
rect -2560 11350 -2320 11590
rect -2230 11350 -1990 11590
rect -1900 11350 -1660 11590
rect -1570 11350 -1330 11590
rect -1240 11350 -1000 11590
rect -910 11350 -670 11590
rect -580 11350 -340 11590
rect -250 11350 -10 11590
rect 80 11350 320 11590
rect 410 11350 650 11590
rect 740 11350 980 11590
rect 1070 11350 1310 11590
rect 1400 11350 1640 11590
rect 1730 11350 1970 11590
rect 2060 11350 2300 11590
rect 2390 11350 2630 11590
rect 2720 11350 2960 11590
rect 3050 11350 3290 11590
rect 3380 11350 3620 11590
rect 3710 11350 3950 11590
rect 4040 11350 4280 11590
rect 4370 11350 4610 11590
rect 4700 11350 4940 11590
rect 5030 11350 5270 11590
rect 5360 11350 5600 11590
rect 5690 11350 5930 11590
rect 6020 11350 6260 11590
rect 6350 11350 6590 11590
rect -5200 11020 -4960 11260
rect -4870 11020 -4630 11260
rect -4540 11020 -4300 11260
rect -4210 11020 -3970 11260
rect -3880 11020 -3640 11260
rect -3550 11020 -3310 11260
rect -3220 11020 -2980 11260
rect -2890 11020 -2650 11260
rect -2560 11020 -2320 11260
rect -2230 11020 -1990 11260
rect -1900 11020 -1660 11260
rect -1570 11020 -1330 11260
rect -1240 11020 -1000 11260
rect -910 11020 -670 11260
rect -580 11020 -340 11260
rect -250 11020 -10 11260
rect 80 11020 320 11260
rect 410 11020 650 11260
rect 740 11020 980 11260
rect 1070 11020 1310 11260
rect 1400 11020 1640 11260
rect 1730 11020 1970 11260
rect 2060 11020 2300 11260
rect 2390 11020 2630 11260
rect 2720 11020 2960 11260
rect 3050 11020 3290 11260
rect 3380 11020 3620 11260
rect 3710 11020 3950 11260
rect 4040 11020 4280 11260
rect 4370 11020 4610 11260
rect 4700 11020 4940 11260
rect 5030 11020 5270 11260
rect 5360 11020 5600 11260
rect 5690 11020 5930 11260
rect 6020 11020 6260 11260
rect 6350 11020 6590 11260
rect -5200 10690 -4960 10930
rect -4870 10690 -4630 10930
rect -4540 10690 -4300 10930
rect -4210 10690 -3970 10930
rect -3880 10690 -3640 10930
rect -3550 10690 -3310 10930
rect -3220 10690 -2980 10930
rect -2890 10690 -2650 10930
rect -2560 10690 -2320 10930
rect -2230 10690 -1990 10930
rect -1900 10690 -1660 10930
rect -1570 10690 -1330 10930
rect -1240 10690 -1000 10930
rect -910 10690 -670 10930
rect -580 10690 -340 10930
rect -250 10690 -10 10930
rect 80 10690 320 10930
rect 410 10690 650 10930
rect 740 10690 980 10930
rect 1070 10690 1310 10930
rect 1400 10690 1640 10930
rect 1730 10690 1970 10930
rect 2060 10690 2300 10930
rect 2390 10690 2630 10930
rect 2720 10690 2960 10930
rect 3050 10690 3290 10930
rect 3380 10690 3620 10930
rect 3710 10690 3950 10930
rect 4040 10690 4280 10930
rect 4370 10690 4610 10930
rect 4700 10690 4940 10930
rect 5030 10690 5270 10930
rect 5360 10690 5600 10930
rect 5690 10690 5930 10930
rect 6020 10690 6260 10930
rect 6350 10690 6590 10930
rect -5200 10360 -4960 10600
rect -4870 10360 -4630 10600
rect -4540 10360 -4300 10600
rect -4210 10360 -3970 10600
rect -3880 10360 -3640 10600
rect -3550 10360 -3310 10600
rect -3220 10360 -2980 10600
rect -2890 10360 -2650 10600
rect -2560 10360 -2320 10600
rect -2230 10360 -1990 10600
rect -1900 10360 -1660 10600
rect -1570 10360 -1330 10600
rect -1240 10360 -1000 10600
rect -910 10360 -670 10600
rect -580 10360 -340 10600
rect -250 10360 -10 10600
rect 80 10360 320 10600
rect 410 10360 650 10600
rect 740 10360 980 10600
rect 1070 10360 1310 10600
rect 1400 10360 1640 10600
rect 1730 10360 1970 10600
rect 2060 10360 2300 10600
rect 2390 10360 2630 10600
rect 2720 10360 2960 10600
rect 3050 10360 3290 10600
rect 3380 10360 3620 10600
rect 3710 10360 3950 10600
rect 4040 10360 4280 10600
rect 4370 10360 4610 10600
rect 4700 10360 4940 10600
rect 5030 10360 5270 10600
rect 5360 10360 5600 10600
rect 5690 10360 5930 10600
rect 6020 10360 6260 10600
rect 6350 10360 6590 10600
rect -5200 10030 -4960 10270
rect -4870 10030 -4630 10270
rect -4540 10030 -4300 10270
rect -4210 10030 -3970 10270
rect -3880 10030 -3640 10270
rect -3550 10030 -3310 10270
rect -3220 10030 -2980 10270
rect -2890 10030 -2650 10270
rect -2560 10030 -2320 10270
rect -2230 10030 -1990 10270
rect -1900 10030 -1660 10270
rect -1570 10030 -1330 10270
rect -1240 10030 -1000 10270
rect -910 10030 -670 10270
rect -580 10030 -340 10270
rect -250 10030 -10 10270
rect 80 10030 320 10270
rect 410 10030 650 10270
rect 740 10030 980 10270
rect 1070 10030 1310 10270
rect 1400 10030 1640 10270
rect 1730 10030 1970 10270
rect 2060 10030 2300 10270
rect 2390 10030 2630 10270
rect 2720 10030 2960 10270
rect 3050 10030 3290 10270
rect 3380 10030 3620 10270
rect 3710 10030 3950 10270
rect 4040 10030 4280 10270
rect 4370 10030 4610 10270
rect 4700 10030 4940 10270
rect 5030 10030 5270 10270
rect 5360 10030 5600 10270
rect 5690 10030 5930 10270
rect 6020 10030 6260 10270
rect 6350 10030 6590 10270
rect -5200 9700 -4960 9940
rect -4870 9700 -4630 9940
rect -4540 9700 -4300 9940
rect -4210 9700 -3970 9940
rect -3880 9700 -3640 9940
rect -3550 9700 -3310 9940
rect -3220 9700 -2980 9940
rect -2890 9700 -2650 9940
rect -2560 9700 -2320 9940
rect -2230 9700 -1990 9940
rect -1900 9700 -1660 9940
rect -1570 9700 -1330 9940
rect -1240 9700 -1000 9940
rect -910 9700 -670 9940
rect -580 9700 -340 9940
rect -250 9700 -10 9940
rect 80 9700 320 9940
rect 410 9700 650 9940
rect 740 9700 980 9940
rect 1070 9700 1310 9940
rect 1400 9700 1640 9940
rect 1730 9700 1970 9940
rect 2060 9700 2300 9940
rect 2390 9700 2630 9940
rect 2720 9700 2960 9940
rect 3050 9700 3290 9940
rect 3380 9700 3620 9940
rect 3710 9700 3950 9940
rect 4040 9700 4280 9940
rect 4370 9700 4610 9940
rect 4700 9700 4940 9940
rect 5030 9700 5270 9940
rect 5360 9700 5600 9940
rect 5690 9700 5930 9940
rect 6020 9700 6260 9940
rect 6350 9700 6590 9940
rect -5200 9370 -4960 9610
rect -4870 9370 -4630 9610
rect -4540 9370 -4300 9610
rect -4210 9370 -3970 9610
rect -3880 9370 -3640 9610
rect -3550 9370 -3310 9610
rect -3220 9370 -2980 9610
rect -2890 9370 -2650 9610
rect -2560 9370 -2320 9610
rect -2230 9370 -1990 9610
rect -1900 9370 -1660 9610
rect -1570 9370 -1330 9610
rect -1240 9370 -1000 9610
rect -910 9370 -670 9610
rect -580 9370 -340 9610
rect -250 9370 -10 9610
rect 80 9370 320 9610
rect 410 9370 650 9610
rect 740 9370 980 9610
rect 1070 9370 1310 9610
rect 1400 9370 1640 9610
rect 1730 9370 1970 9610
rect 2060 9370 2300 9610
rect 2390 9370 2630 9610
rect 2720 9370 2960 9610
rect 3050 9370 3290 9610
rect 3380 9370 3620 9610
rect 3710 9370 3950 9610
rect 4040 9370 4280 9610
rect 4370 9370 4610 9610
rect 4700 9370 4940 9610
rect 5030 9370 5270 9610
rect 5360 9370 5600 9610
rect 5690 9370 5930 9610
rect 6020 9370 6260 9610
rect 6350 9370 6590 9610
rect -5200 9040 -4960 9280
rect -4870 9040 -4630 9280
rect -4540 9040 -4300 9280
rect -4210 9040 -3970 9280
rect -3880 9040 -3640 9280
rect -3550 9040 -3310 9280
rect -3220 9040 -2980 9280
rect -2890 9040 -2650 9280
rect -2560 9040 -2320 9280
rect -2230 9040 -1990 9280
rect -1900 9040 -1660 9280
rect -1570 9040 -1330 9280
rect -1240 9040 -1000 9280
rect -910 9040 -670 9280
rect -580 9040 -340 9280
rect -250 9040 -10 9280
rect 80 9040 320 9280
rect 410 9040 650 9280
rect 740 9040 980 9280
rect 1070 9040 1310 9280
rect 1400 9040 1640 9280
rect 1730 9040 1970 9280
rect 2060 9040 2300 9280
rect 2390 9040 2630 9280
rect 2720 9040 2960 9280
rect 3050 9040 3290 9280
rect 3380 9040 3620 9280
rect 3710 9040 3950 9280
rect 4040 9040 4280 9280
rect 4370 9040 4610 9280
rect 4700 9040 4940 9280
rect 5030 9040 5270 9280
rect 5360 9040 5600 9280
rect 5690 9040 5930 9280
rect 6020 9040 6260 9280
rect 6350 9040 6590 9280
rect 8310 20590 8550 20830
rect 8640 20590 8880 20830
rect 8970 20590 9210 20830
rect 9300 20590 9540 20830
rect 9630 20590 9870 20830
rect 9960 20590 10200 20830
rect 10290 20590 10530 20830
rect 10620 20590 10860 20830
rect 10950 20590 11190 20830
rect 11280 20590 11520 20830
rect 11610 20590 11850 20830
rect 11940 20590 12180 20830
rect 12270 20590 12510 20830
rect 12600 20590 12840 20830
rect 12930 20590 13170 20830
rect 13260 20590 13500 20830
rect 13590 20590 13830 20830
rect 13920 20590 14160 20830
rect 14250 20590 14490 20830
rect 14580 20590 14820 20830
rect 14910 20590 15150 20830
rect 15240 20590 15480 20830
rect 15570 20590 15810 20830
rect 15900 20590 16140 20830
rect 16230 20590 16470 20830
rect 16560 20590 16800 20830
rect 16890 20590 17130 20830
rect 17220 20590 17460 20830
rect 17550 20590 17790 20830
rect 17880 20590 18120 20830
rect 18210 20590 18450 20830
rect 18540 20590 18780 20830
rect 18870 20590 19110 20830
rect 19200 20590 19440 20830
rect 19530 20590 19770 20830
rect 19860 20590 20100 20830
rect 8310 20260 8550 20500
rect 8640 20260 8880 20500
rect 8970 20260 9210 20500
rect 9300 20260 9540 20500
rect 9630 20260 9870 20500
rect 9960 20260 10200 20500
rect 10290 20260 10530 20500
rect 10620 20260 10860 20500
rect 10950 20260 11190 20500
rect 11280 20260 11520 20500
rect 11610 20260 11850 20500
rect 11940 20260 12180 20500
rect 12270 20260 12510 20500
rect 12600 20260 12840 20500
rect 12930 20260 13170 20500
rect 13260 20260 13500 20500
rect 13590 20260 13830 20500
rect 13920 20260 14160 20500
rect 14250 20260 14490 20500
rect 14580 20260 14820 20500
rect 14910 20260 15150 20500
rect 15240 20260 15480 20500
rect 15570 20260 15810 20500
rect 15900 20260 16140 20500
rect 16230 20260 16470 20500
rect 16560 20260 16800 20500
rect 16890 20260 17130 20500
rect 17220 20260 17460 20500
rect 17550 20260 17790 20500
rect 17880 20260 18120 20500
rect 18210 20260 18450 20500
rect 18540 20260 18780 20500
rect 18870 20260 19110 20500
rect 19200 20260 19440 20500
rect 19530 20260 19770 20500
rect 19860 20260 20100 20500
rect 8310 19930 8550 20170
rect 8640 19930 8880 20170
rect 8970 19930 9210 20170
rect 9300 19930 9540 20170
rect 9630 19930 9870 20170
rect 9960 19930 10200 20170
rect 10290 19930 10530 20170
rect 10620 19930 10860 20170
rect 10950 19930 11190 20170
rect 11280 19930 11520 20170
rect 11610 19930 11850 20170
rect 11940 19930 12180 20170
rect 12270 19930 12510 20170
rect 12600 19930 12840 20170
rect 12930 19930 13170 20170
rect 13260 19930 13500 20170
rect 13590 19930 13830 20170
rect 13920 19930 14160 20170
rect 14250 19930 14490 20170
rect 14580 19930 14820 20170
rect 14910 19930 15150 20170
rect 15240 19930 15480 20170
rect 15570 19930 15810 20170
rect 15900 19930 16140 20170
rect 16230 19930 16470 20170
rect 16560 19930 16800 20170
rect 16890 19930 17130 20170
rect 17220 19930 17460 20170
rect 17550 19930 17790 20170
rect 17880 19930 18120 20170
rect 18210 19930 18450 20170
rect 18540 19930 18780 20170
rect 18870 19930 19110 20170
rect 19200 19930 19440 20170
rect 19530 19930 19770 20170
rect 19860 19930 20100 20170
rect 8310 19600 8550 19840
rect 8640 19600 8880 19840
rect 8970 19600 9210 19840
rect 9300 19600 9540 19840
rect 9630 19600 9870 19840
rect 9960 19600 10200 19840
rect 10290 19600 10530 19840
rect 10620 19600 10860 19840
rect 10950 19600 11190 19840
rect 11280 19600 11520 19840
rect 11610 19600 11850 19840
rect 11940 19600 12180 19840
rect 12270 19600 12510 19840
rect 12600 19600 12840 19840
rect 12930 19600 13170 19840
rect 13260 19600 13500 19840
rect 13590 19600 13830 19840
rect 13920 19600 14160 19840
rect 14250 19600 14490 19840
rect 14580 19600 14820 19840
rect 14910 19600 15150 19840
rect 15240 19600 15480 19840
rect 15570 19600 15810 19840
rect 15900 19600 16140 19840
rect 16230 19600 16470 19840
rect 16560 19600 16800 19840
rect 16890 19600 17130 19840
rect 17220 19600 17460 19840
rect 17550 19600 17790 19840
rect 17880 19600 18120 19840
rect 18210 19600 18450 19840
rect 18540 19600 18780 19840
rect 18870 19600 19110 19840
rect 19200 19600 19440 19840
rect 19530 19600 19770 19840
rect 19860 19600 20100 19840
rect 8310 19270 8550 19510
rect 8640 19270 8880 19510
rect 8970 19270 9210 19510
rect 9300 19270 9540 19510
rect 9630 19270 9870 19510
rect 9960 19270 10200 19510
rect 10290 19270 10530 19510
rect 10620 19270 10860 19510
rect 10950 19270 11190 19510
rect 11280 19270 11520 19510
rect 11610 19270 11850 19510
rect 11940 19270 12180 19510
rect 12270 19270 12510 19510
rect 12600 19270 12840 19510
rect 12930 19270 13170 19510
rect 13260 19270 13500 19510
rect 13590 19270 13830 19510
rect 13920 19270 14160 19510
rect 14250 19270 14490 19510
rect 14580 19270 14820 19510
rect 14910 19270 15150 19510
rect 15240 19270 15480 19510
rect 15570 19270 15810 19510
rect 15900 19270 16140 19510
rect 16230 19270 16470 19510
rect 16560 19270 16800 19510
rect 16890 19270 17130 19510
rect 17220 19270 17460 19510
rect 17550 19270 17790 19510
rect 17880 19270 18120 19510
rect 18210 19270 18450 19510
rect 18540 19270 18780 19510
rect 18870 19270 19110 19510
rect 19200 19270 19440 19510
rect 19530 19270 19770 19510
rect 19860 19270 20100 19510
rect 8310 18940 8550 19180
rect 8640 18940 8880 19180
rect 8970 18940 9210 19180
rect 9300 18940 9540 19180
rect 9630 18940 9870 19180
rect 9960 18940 10200 19180
rect 10290 18940 10530 19180
rect 10620 18940 10860 19180
rect 10950 18940 11190 19180
rect 11280 18940 11520 19180
rect 11610 18940 11850 19180
rect 11940 18940 12180 19180
rect 12270 18940 12510 19180
rect 12600 18940 12840 19180
rect 12930 18940 13170 19180
rect 13260 18940 13500 19180
rect 13590 18940 13830 19180
rect 13920 18940 14160 19180
rect 14250 18940 14490 19180
rect 14580 18940 14820 19180
rect 14910 18940 15150 19180
rect 15240 18940 15480 19180
rect 15570 18940 15810 19180
rect 15900 18940 16140 19180
rect 16230 18940 16470 19180
rect 16560 18940 16800 19180
rect 16890 18940 17130 19180
rect 17220 18940 17460 19180
rect 17550 18940 17790 19180
rect 17880 18940 18120 19180
rect 18210 18940 18450 19180
rect 18540 18940 18780 19180
rect 18870 18940 19110 19180
rect 19200 18940 19440 19180
rect 19530 18940 19770 19180
rect 19860 18940 20100 19180
rect 8310 18610 8550 18850
rect 8640 18610 8880 18850
rect 8970 18610 9210 18850
rect 9300 18610 9540 18850
rect 9630 18610 9870 18850
rect 9960 18610 10200 18850
rect 10290 18610 10530 18850
rect 10620 18610 10860 18850
rect 10950 18610 11190 18850
rect 11280 18610 11520 18850
rect 11610 18610 11850 18850
rect 11940 18610 12180 18850
rect 12270 18610 12510 18850
rect 12600 18610 12840 18850
rect 12930 18610 13170 18850
rect 13260 18610 13500 18850
rect 13590 18610 13830 18850
rect 13920 18610 14160 18850
rect 14250 18610 14490 18850
rect 14580 18610 14820 18850
rect 14910 18610 15150 18850
rect 15240 18610 15480 18850
rect 15570 18610 15810 18850
rect 15900 18610 16140 18850
rect 16230 18610 16470 18850
rect 16560 18610 16800 18850
rect 16890 18610 17130 18850
rect 17220 18610 17460 18850
rect 17550 18610 17790 18850
rect 17880 18610 18120 18850
rect 18210 18610 18450 18850
rect 18540 18610 18780 18850
rect 18870 18610 19110 18850
rect 19200 18610 19440 18850
rect 19530 18610 19770 18850
rect 19860 18610 20100 18850
rect 8310 18280 8550 18520
rect 8640 18280 8880 18520
rect 8970 18280 9210 18520
rect 9300 18280 9540 18520
rect 9630 18280 9870 18520
rect 9960 18280 10200 18520
rect 10290 18280 10530 18520
rect 10620 18280 10860 18520
rect 10950 18280 11190 18520
rect 11280 18280 11520 18520
rect 11610 18280 11850 18520
rect 11940 18280 12180 18520
rect 12270 18280 12510 18520
rect 12600 18280 12840 18520
rect 12930 18280 13170 18520
rect 13260 18280 13500 18520
rect 13590 18280 13830 18520
rect 13920 18280 14160 18520
rect 14250 18280 14490 18520
rect 14580 18280 14820 18520
rect 14910 18280 15150 18520
rect 15240 18280 15480 18520
rect 15570 18280 15810 18520
rect 15900 18280 16140 18520
rect 16230 18280 16470 18520
rect 16560 18280 16800 18520
rect 16890 18280 17130 18520
rect 17220 18280 17460 18520
rect 17550 18280 17790 18520
rect 17880 18280 18120 18520
rect 18210 18280 18450 18520
rect 18540 18280 18780 18520
rect 18870 18280 19110 18520
rect 19200 18280 19440 18520
rect 19530 18280 19770 18520
rect 19860 18280 20100 18520
rect 8310 17950 8550 18190
rect 8640 17950 8880 18190
rect 8970 17950 9210 18190
rect 9300 17950 9540 18190
rect 9630 17950 9870 18190
rect 9960 17950 10200 18190
rect 10290 17950 10530 18190
rect 10620 17950 10860 18190
rect 10950 17950 11190 18190
rect 11280 17950 11520 18190
rect 11610 17950 11850 18190
rect 11940 17950 12180 18190
rect 12270 17950 12510 18190
rect 12600 17950 12840 18190
rect 12930 17950 13170 18190
rect 13260 17950 13500 18190
rect 13590 17950 13830 18190
rect 13920 17950 14160 18190
rect 14250 17950 14490 18190
rect 14580 17950 14820 18190
rect 14910 17950 15150 18190
rect 15240 17950 15480 18190
rect 15570 17950 15810 18190
rect 15900 17950 16140 18190
rect 16230 17950 16470 18190
rect 16560 17950 16800 18190
rect 16890 17950 17130 18190
rect 17220 17950 17460 18190
rect 17550 17950 17790 18190
rect 17880 17950 18120 18190
rect 18210 17950 18450 18190
rect 18540 17950 18780 18190
rect 18870 17950 19110 18190
rect 19200 17950 19440 18190
rect 19530 17950 19770 18190
rect 19860 17950 20100 18190
rect 8310 17620 8550 17860
rect 8640 17620 8880 17860
rect 8970 17620 9210 17860
rect 9300 17620 9540 17860
rect 9630 17620 9870 17860
rect 9960 17620 10200 17860
rect 10290 17620 10530 17860
rect 10620 17620 10860 17860
rect 10950 17620 11190 17860
rect 11280 17620 11520 17860
rect 11610 17620 11850 17860
rect 11940 17620 12180 17860
rect 12270 17620 12510 17860
rect 12600 17620 12840 17860
rect 12930 17620 13170 17860
rect 13260 17620 13500 17860
rect 13590 17620 13830 17860
rect 13920 17620 14160 17860
rect 14250 17620 14490 17860
rect 14580 17620 14820 17860
rect 14910 17620 15150 17860
rect 15240 17620 15480 17860
rect 15570 17620 15810 17860
rect 15900 17620 16140 17860
rect 16230 17620 16470 17860
rect 16560 17620 16800 17860
rect 16890 17620 17130 17860
rect 17220 17620 17460 17860
rect 17550 17620 17790 17860
rect 17880 17620 18120 17860
rect 18210 17620 18450 17860
rect 18540 17620 18780 17860
rect 18870 17620 19110 17860
rect 19200 17620 19440 17860
rect 19530 17620 19770 17860
rect 19860 17620 20100 17860
rect 8310 17290 8550 17530
rect 8640 17290 8880 17530
rect 8970 17290 9210 17530
rect 9300 17290 9540 17530
rect 9630 17290 9870 17530
rect 9960 17290 10200 17530
rect 10290 17290 10530 17530
rect 10620 17290 10860 17530
rect 10950 17290 11190 17530
rect 11280 17290 11520 17530
rect 11610 17290 11850 17530
rect 11940 17290 12180 17530
rect 12270 17290 12510 17530
rect 12600 17290 12840 17530
rect 12930 17290 13170 17530
rect 13260 17290 13500 17530
rect 13590 17290 13830 17530
rect 13920 17290 14160 17530
rect 14250 17290 14490 17530
rect 14580 17290 14820 17530
rect 14910 17290 15150 17530
rect 15240 17290 15480 17530
rect 15570 17290 15810 17530
rect 15900 17290 16140 17530
rect 16230 17290 16470 17530
rect 16560 17290 16800 17530
rect 16890 17290 17130 17530
rect 17220 17290 17460 17530
rect 17550 17290 17790 17530
rect 17880 17290 18120 17530
rect 18210 17290 18450 17530
rect 18540 17290 18780 17530
rect 18870 17290 19110 17530
rect 19200 17290 19440 17530
rect 19530 17290 19770 17530
rect 19860 17290 20100 17530
rect 8310 16960 8550 17200
rect 8640 16960 8880 17200
rect 8970 16960 9210 17200
rect 9300 16960 9540 17200
rect 9630 16960 9870 17200
rect 9960 16960 10200 17200
rect 10290 16960 10530 17200
rect 10620 16960 10860 17200
rect 10950 16960 11190 17200
rect 11280 16960 11520 17200
rect 11610 16960 11850 17200
rect 11940 16960 12180 17200
rect 12270 16960 12510 17200
rect 12600 16960 12840 17200
rect 12930 16960 13170 17200
rect 13260 16960 13500 17200
rect 13590 16960 13830 17200
rect 13920 16960 14160 17200
rect 14250 16960 14490 17200
rect 14580 16960 14820 17200
rect 14910 16960 15150 17200
rect 15240 16960 15480 17200
rect 15570 16960 15810 17200
rect 15900 16960 16140 17200
rect 16230 16960 16470 17200
rect 16560 16960 16800 17200
rect 16890 16960 17130 17200
rect 17220 16960 17460 17200
rect 17550 16960 17790 17200
rect 17880 16960 18120 17200
rect 18210 16960 18450 17200
rect 18540 16960 18780 17200
rect 18870 16960 19110 17200
rect 19200 16960 19440 17200
rect 19530 16960 19770 17200
rect 19860 16960 20100 17200
rect 8310 16630 8550 16870
rect 8640 16630 8880 16870
rect 8970 16630 9210 16870
rect 9300 16630 9540 16870
rect 9630 16630 9870 16870
rect 9960 16630 10200 16870
rect 10290 16630 10530 16870
rect 10620 16630 10860 16870
rect 10950 16630 11190 16870
rect 11280 16630 11520 16870
rect 11610 16630 11850 16870
rect 11940 16630 12180 16870
rect 12270 16630 12510 16870
rect 12600 16630 12840 16870
rect 12930 16630 13170 16870
rect 13260 16630 13500 16870
rect 13590 16630 13830 16870
rect 13920 16630 14160 16870
rect 14250 16630 14490 16870
rect 14580 16630 14820 16870
rect 14910 16630 15150 16870
rect 15240 16630 15480 16870
rect 15570 16630 15810 16870
rect 15900 16630 16140 16870
rect 16230 16630 16470 16870
rect 16560 16630 16800 16870
rect 16890 16630 17130 16870
rect 17220 16630 17460 16870
rect 17550 16630 17790 16870
rect 17880 16630 18120 16870
rect 18210 16630 18450 16870
rect 18540 16630 18780 16870
rect 18870 16630 19110 16870
rect 19200 16630 19440 16870
rect 19530 16630 19770 16870
rect 19860 16630 20100 16870
rect 8310 16300 8550 16540
rect 8640 16300 8880 16540
rect 8970 16300 9210 16540
rect 9300 16300 9540 16540
rect 9630 16300 9870 16540
rect 9960 16300 10200 16540
rect 10290 16300 10530 16540
rect 10620 16300 10860 16540
rect 10950 16300 11190 16540
rect 11280 16300 11520 16540
rect 11610 16300 11850 16540
rect 11940 16300 12180 16540
rect 12270 16300 12510 16540
rect 12600 16300 12840 16540
rect 12930 16300 13170 16540
rect 13260 16300 13500 16540
rect 13590 16300 13830 16540
rect 13920 16300 14160 16540
rect 14250 16300 14490 16540
rect 14580 16300 14820 16540
rect 14910 16300 15150 16540
rect 15240 16300 15480 16540
rect 15570 16300 15810 16540
rect 15900 16300 16140 16540
rect 16230 16300 16470 16540
rect 16560 16300 16800 16540
rect 16890 16300 17130 16540
rect 17220 16300 17460 16540
rect 17550 16300 17790 16540
rect 17880 16300 18120 16540
rect 18210 16300 18450 16540
rect 18540 16300 18780 16540
rect 18870 16300 19110 16540
rect 19200 16300 19440 16540
rect 19530 16300 19770 16540
rect 19860 16300 20100 16540
rect 8310 15970 8550 16210
rect 8640 15970 8880 16210
rect 8970 15970 9210 16210
rect 9300 15970 9540 16210
rect 9630 15970 9870 16210
rect 9960 15970 10200 16210
rect 10290 15970 10530 16210
rect 10620 15970 10860 16210
rect 10950 15970 11190 16210
rect 11280 15970 11520 16210
rect 11610 15970 11850 16210
rect 11940 15970 12180 16210
rect 12270 15970 12510 16210
rect 12600 15970 12840 16210
rect 12930 15970 13170 16210
rect 13260 15970 13500 16210
rect 13590 15970 13830 16210
rect 13920 15970 14160 16210
rect 14250 15970 14490 16210
rect 14580 15970 14820 16210
rect 14910 15970 15150 16210
rect 15240 15970 15480 16210
rect 15570 15970 15810 16210
rect 15900 15970 16140 16210
rect 16230 15970 16470 16210
rect 16560 15970 16800 16210
rect 16890 15970 17130 16210
rect 17220 15970 17460 16210
rect 17550 15970 17790 16210
rect 17880 15970 18120 16210
rect 18210 15970 18450 16210
rect 18540 15970 18780 16210
rect 18870 15970 19110 16210
rect 19200 15970 19440 16210
rect 19530 15970 19770 16210
rect 19860 15970 20100 16210
rect 8310 15640 8550 15880
rect 8640 15640 8880 15880
rect 8970 15640 9210 15880
rect 9300 15640 9540 15880
rect 9630 15640 9870 15880
rect 9960 15640 10200 15880
rect 10290 15640 10530 15880
rect 10620 15640 10860 15880
rect 10950 15640 11190 15880
rect 11280 15640 11520 15880
rect 11610 15640 11850 15880
rect 11940 15640 12180 15880
rect 12270 15640 12510 15880
rect 12600 15640 12840 15880
rect 12930 15640 13170 15880
rect 13260 15640 13500 15880
rect 13590 15640 13830 15880
rect 13920 15640 14160 15880
rect 14250 15640 14490 15880
rect 14580 15640 14820 15880
rect 14910 15640 15150 15880
rect 15240 15640 15480 15880
rect 15570 15640 15810 15880
rect 15900 15640 16140 15880
rect 16230 15640 16470 15880
rect 16560 15640 16800 15880
rect 16890 15640 17130 15880
rect 17220 15640 17460 15880
rect 17550 15640 17790 15880
rect 17880 15640 18120 15880
rect 18210 15640 18450 15880
rect 18540 15640 18780 15880
rect 18870 15640 19110 15880
rect 19200 15640 19440 15880
rect 19530 15640 19770 15880
rect 19860 15640 20100 15880
rect 8310 15310 8550 15550
rect 8640 15310 8880 15550
rect 8970 15310 9210 15550
rect 9300 15310 9540 15550
rect 9630 15310 9870 15550
rect 9960 15310 10200 15550
rect 10290 15310 10530 15550
rect 10620 15310 10860 15550
rect 10950 15310 11190 15550
rect 11280 15310 11520 15550
rect 11610 15310 11850 15550
rect 11940 15310 12180 15550
rect 12270 15310 12510 15550
rect 12600 15310 12840 15550
rect 12930 15310 13170 15550
rect 13260 15310 13500 15550
rect 13590 15310 13830 15550
rect 13920 15310 14160 15550
rect 14250 15310 14490 15550
rect 14580 15310 14820 15550
rect 14910 15310 15150 15550
rect 15240 15310 15480 15550
rect 15570 15310 15810 15550
rect 15900 15310 16140 15550
rect 16230 15310 16470 15550
rect 16560 15310 16800 15550
rect 16890 15310 17130 15550
rect 17220 15310 17460 15550
rect 17550 15310 17790 15550
rect 17880 15310 18120 15550
rect 18210 15310 18450 15550
rect 18540 15310 18780 15550
rect 18870 15310 19110 15550
rect 19200 15310 19440 15550
rect 19530 15310 19770 15550
rect 19860 15310 20100 15550
rect 8310 14980 8550 15220
rect 8640 14980 8880 15220
rect 8970 14980 9210 15220
rect 9300 14980 9540 15220
rect 9630 14980 9870 15220
rect 9960 14980 10200 15220
rect 10290 14980 10530 15220
rect 10620 14980 10860 15220
rect 10950 14980 11190 15220
rect 11280 14980 11520 15220
rect 11610 14980 11850 15220
rect 11940 14980 12180 15220
rect 12270 14980 12510 15220
rect 12600 14980 12840 15220
rect 12930 14980 13170 15220
rect 13260 14980 13500 15220
rect 13590 14980 13830 15220
rect 13920 14980 14160 15220
rect 14250 14980 14490 15220
rect 14580 14980 14820 15220
rect 14910 14980 15150 15220
rect 15240 14980 15480 15220
rect 15570 14980 15810 15220
rect 15900 14980 16140 15220
rect 16230 14980 16470 15220
rect 16560 14980 16800 15220
rect 16890 14980 17130 15220
rect 17220 14980 17460 15220
rect 17550 14980 17790 15220
rect 17880 14980 18120 15220
rect 18210 14980 18450 15220
rect 18540 14980 18780 15220
rect 18870 14980 19110 15220
rect 19200 14980 19440 15220
rect 19530 14980 19770 15220
rect 19860 14980 20100 15220
rect 8310 14650 8550 14890
rect 8640 14650 8880 14890
rect 8970 14650 9210 14890
rect 9300 14650 9540 14890
rect 9630 14650 9870 14890
rect 9960 14650 10200 14890
rect 10290 14650 10530 14890
rect 10620 14650 10860 14890
rect 10950 14650 11190 14890
rect 11280 14650 11520 14890
rect 11610 14650 11850 14890
rect 11940 14650 12180 14890
rect 12270 14650 12510 14890
rect 12600 14650 12840 14890
rect 12930 14650 13170 14890
rect 13260 14650 13500 14890
rect 13590 14650 13830 14890
rect 13920 14650 14160 14890
rect 14250 14650 14490 14890
rect 14580 14650 14820 14890
rect 14910 14650 15150 14890
rect 15240 14650 15480 14890
rect 15570 14650 15810 14890
rect 15900 14650 16140 14890
rect 16230 14650 16470 14890
rect 16560 14650 16800 14890
rect 16890 14650 17130 14890
rect 17220 14650 17460 14890
rect 17550 14650 17790 14890
rect 17880 14650 18120 14890
rect 18210 14650 18450 14890
rect 18540 14650 18780 14890
rect 18870 14650 19110 14890
rect 19200 14650 19440 14890
rect 19530 14650 19770 14890
rect 19860 14650 20100 14890
rect 8310 14320 8550 14560
rect 8640 14320 8880 14560
rect 8970 14320 9210 14560
rect 9300 14320 9540 14560
rect 9630 14320 9870 14560
rect 9960 14320 10200 14560
rect 10290 14320 10530 14560
rect 10620 14320 10860 14560
rect 10950 14320 11190 14560
rect 11280 14320 11520 14560
rect 11610 14320 11850 14560
rect 11940 14320 12180 14560
rect 12270 14320 12510 14560
rect 12600 14320 12840 14560
rect 12930 14320 13170 14560
rect 13260 14320 13500 14560
rect 13590 14320 13830 14560
rect 13920 14320 14160 14560
rect 14250 14320 14490 14560
rect 14580 14320 14820 14560
rect 14910 14320 15150 14560
rect 15240 14320 15480 14560
rect 15570 14320 15810 14560
rect 15900 14320 16140 14560
rect 16230 14320 16470 14560
rect 16560 14320 16800 14560
rect 16890 14320 17130 14560
rect 17220 14320 17460 14560
rect 17550 14320 17790 14560
rect 17880 14320 18120 14560
rect 18210 14320 18450 14560
rect 18540 14320 18780 14560
rect 18870 14320 19110 14560
rect 19200 14320 19440 14560
rect 19530 14320 19770 14560
rect 19860 14320 20100 14560
rect 8310 13990 8550 14230
rect 8640 13990 8880 14230
rect 8970 13990 9210 14230
rect 9300 13990 9540 14230
rect 9630 13990 9870 14230
rect 9960 13990 10200 14230
rect 10290 13990 10530 14230
rect 10620 13990 10860 14230
rect 10950 13990 11190 14230
rect 11280 13990 11520 14230
rect 11610 13990 11850 14230
rect 11940 13990 12180 14230
rect 12270 13990 12510 14230
rect 12600 13990 12840 14230
rect 12930 13990 13170 14230
rect 13260 13990 13500 14230
rect 13590 13990 13830 14230
rect 13920 13990 14160 14230
rect 14250 13990 14490 14230
rect 14580 13990 14820 14230
rect 14910 13990 15150 14230
rect 15240 13990 15480 14230
rect 15570 13990 15810 14230
rect 15900 13990 16140 14230
rect 16230 13990 16470 14230
rect 16560 13990 16800 14230
rect 16890 13990 17130 14230
rect 17220 13990 17460 14230
rect 17550 13990 17790 14230
rect 17880 13990 18120 14230
rect 18210 13990 18450 14230
rect 18540 13990 18780 14230
rect 18870 13990 19110 14230
rect 19200 13990 19440 14230
rect 19530 13990 19770 14230
rect 19860 13990 20100 14230
rect 8310 13660 8550 13900
rect 8640 13660 8880 13900
rect 8970 13660 9210 13900
rect 9300 13660 9540 13900
rect 9630 13660 9870 13900
rect 9960 13660 10200 13900
rect 10290 13660 10530 13900
rect 10620 13660 10860 13900
rect 10950 13660 11190 13900
rect 11280 13660 11520 13900
rect 11610 13660 11850 13900
rect 11940 13660 12180 13900
rect 12270 13660 12510 13900
rect 12600 13660 12840 13900
rect 12930 13660 13170 13900
rect 13260 13660 13500 13900
rect 13590 13660 13830 13900
rect 13920 13660 14160 13900
rect 14250 13660 14490 13900
rect 14580 13660 14820 13900
rect 14910 13660 15150 13900
rect 15240 13660 15480 13900
rect 15570 13660 15810 13900
rect 15900 13660 16140 13900
rect 16230 13660 16470 13900
rect 16560 13660 16800 13900
rect 16890 13660 17130 13900
rect 17220 13660 17460 13900
rect 17550 13660 17790 13900
rect 17880 13660 18120 13900
rect 18210 13660 18450 13900
rect 18540 13660 18780 13900
rect 18870 13660 19110 13900
rect 19200 13660 19440 13900
rect 19530 13660 19770 13900
rect 19860 13660 20100 13900
rect 8310 13330 8550 13570
rect 8640 13330 8880 13570
rect 8970 13330 9210 13570
rect 9300 13330 9540 13570
rect 9630 13330 9870 13570
rect 9960 13330 10200 13570
rect 10290 13330 10530 13570
rect 10620 13330 10860 13570
rect 10950 13330 11190 13570
rect 11280 13330 11520 13570
rect 11610 13330 11850 13570
rect 11940 13330 12180 13570
rect 12270 13330 12510 13570
rect 12600 13330 12840 13570
rect 12930 13330 13170 13570
rect 13260 13330 13500 13570
rect 13590 13330 13830 13570
rect 13920 13330 14160 13570
rect 14250 13330 14490 13570
rect 14580 13330 14820 13570
rect 14910 13330 15150 13570
rect 15240 13330 15480 13570
rect 15570 13330 15810 13570
rect 15900 13330 16140 13570
rect 16230 13330 16470 13570
rect 16560 13330 16800 13570
rect 16890 13330 17130 13570
rect 17220 13330 17460 13570
rect 17550 13330 17790 13570
rect 17880 13330 18120 13570
rect 18210 13330 18450 13570
rect 18540 13330 18780 13570
rect 18870 13330 19110 13570
rect 19200 13330 19440 13570
rect 19530 13330 19770 13570
rect 19860 13330 20100 13570
rect 8310 13000 8550 13240
rect 8640 13000 8880 13240
rect 8970 13000 9210 13240
rect 9300 13000 9540 13240
rect 9630 13000 9870 13240
rect 9960 13000 10200 13240
rect 10290 13000 10530 13240
rect 10620 13000 10860 13240
rect 10950 13000 11190 13240
rect 11280 13000 11520 13240
rect 11610 13000 11850 13240
rect 11940 13000 12180 13240
rect 12270 13000 12510 13240
rect 12600 13000 12840 13240
rect 12930 13000 13170 13240
rect 13260 13000 13500 13240
rect 13590 13000 13830 13240
rect 13920 13000 14160 13240
rect 14250 13000 14490 13240
rect 14580 13000 14820 13240
rect 14910 13000 15150 13240
rect 15240 13000 15480 13240
rect 15570 13000 15810 13240
rect 15900 13000 16140 13240
rect 16230 13000 16470 13240
rect 16560 13000 16800 13240
rect 16890 13000 17130 13240
rect 17220 13000 17460 13240
rect 17550 13000 17790 13240
rect 17880 13000 18120 13240
rect 18210 13000 18450 13240
rect 18540 13000 18780 13240
rect 18870 13000 19110 13240
rect 19200 13000 19440 13240
rect 19530 13000 19770 13240
rect 19860 13000 20100 13240
rect 8310 12670 8550 12910
rect 8640 12670 8880 12910
rect 8970 12670 9210 12910
rect 9300 12670 9540 12910
rect 9630 12670 9870 12910
rect 9960 12670 10200 12910
rect 10290 12670 10530 12910
rect 10620 12670 10860 12910
rect 10950 12670 11190 12910
rect 11280 12670 11520 12910
rect 11610 12670 11850 12910
rect 11940 12670 12180 12910
rect 12270 12670 12510 12910
rect 12600 12670 12840 12910
rect 12930 12670 13170 12910
rect 13260 12670 13500 12910
rect 13590 12670 13830 12910
rect 13920 12670 14160 12910
rect 14250 12670 14490 12910
rect 14580 12670 14820 12910
rect 14910 12670 15150 12910
rect 15240 12670 15480 12910
rect 15570 12670 15810 12910
rect 15900 12670 16140 12910
rect 16230 12670 16470 12910
rect 16560 12670 16800 12910
rect 16890 12670 17130 12910
rect 17220 12670 17460 12910
rect 17550 12670 17790 12910
rect 17880 12670 18120 12910
rect 18210 12670 18450 12910
rect 18540 12670 18780 12910
rect 18870 12670 19110 12910
rect 19200 12670 19440 12910
rect 19530 12670 19770 12910
rect 19860 12670 20100 12910
rect 8310 12340 8550 12580
rect 8640 12340 8880 12580
rect 8970 12340 9210 12580
rect 9300 12340 9540 12580
rect 9630 12340 9870 12580
rect 9960 12340 10200 12580
rect 10290 12340 10530 12580
rect 10620 12340 10860 12580
rect 10950 12340 11190 12580
rect 11280 12340 11520 12580
rect 11610 12340 11850 12580
rect 11940 12340 12180 12580
rect 12270 12340 12510 12580
rect 12600 12340 12840 12580
rect 12930 12340 13170 12580
rect 13260 12340 13500 12580
rect 13590 12340 13830 12580
rect 13920 12340 14160 12580
rect 14250 12340 14490 12580
rect 14580 12340 14820 12580
rect 14910 12340 15150 12580
rect 15240 12340 15480 12580
rect 15570 12340 15810 12580
rect 15900 12340 16140 12580
rect 16230 12340 16470 12580
rect 16560 12340 16800 12580
rect 16890 12340 17130 12580
rect 17220 12340 17460 12580
rect 17550 12340 17790 12580
rect 17880 12340 18120 12580
rect 18210 12340 18450 12580
rect 18540 12340 18780 12580
rect 18870 12340 19110 12580
rect 19200 12340 19440 12580
rect 19530 12340 19770 12580
rect 19860 12340 20100 12580
rect 8310 12010 8550 12250
rect 8640 12010 8880 12250
rect 8970 12010 9210 12250
rect 9300 12010 9540 12250
rect 9630 12010 9870 12250
rect 9960 12010 10200 12250
rect 10290 12010 10530 12250
rect 10620 12010 10860 12250
rect 10950 12010 11190 12250
rect 11280 12010 11520 12250
rect 11610 12010 11850 12250
rect 11940 12010 12180 12250
rect 12270 12010 12510 12250
rect 12600 12010 12840 12250
rect 12930 12010 13170 12250
rect 13260 12010 13500 12250
rect 13590 12010 13830 12250
rect 13920 12010 14160 12250
rect 14250 12010 14490 12250
rect 14580 12010 14820 12250
rect 14910 12010 15150 12250
rect 15240 12010 15480 12250
rect 15570 12010 15810 12250
rect 15900 12010 16140 12250
rect 16230 12010 16470 12250
rect 16560 12010 16800 12250
rect 16890 12010 17130 12250
rect 17220 12010 17460 12250
rect 17550 12010 17790 12250
rect 17880 12010 18120 12250
rect 18210 12010 18450 12250
rect 18540 12010 18780 12250
rect 18870 12010 19110 12250
rect 19200 12010 19440 12250
rect 19530 12010 19770 12250
rect 19860 12010 20100 12250
rect 8310 11680 8550 11920
rect 8640 11680 8880 11920
rect 8970 11680 9210 11920
rect 9300 11680 9540 11920
rect 9630 11680 9870 11920
rect 9960 11680 10200 11920
rect 10290 11680 10530 11920
rect 10620 11680 10860 11920
rect 10950 11680 11190 11920
rect 11280 11680 11520 11920
rect 11610 11680 11850 11920
rect 11940 11680 12180 11920
rect 12270 11680 12510 11920
rect 12600 11680 12840 11920
rect 12930 11680 13170 11920
rect 13260 11680 13500 11920
rect 13590 11680 13830 11920
rect 13920 11680 14160 11920
rect 14250 11680 14490 11920
rect 14580 11680 14820 11920
rect 14910 11680 15150 11920
rect 15240 11680 15480 11920
rect 15570 11680 15810 11920
rect 15900 11680 16140 11920
rect 16230 11680 16470 11920
rect 16560 11680 16800 11920
rect 16890 11680 17130 11920
rect 17220 11680 17460 11920
rect 17550 11680 17790 11920
rect 17880 11680 18120 11920
rect 18210 11680 18450 11920
rect 18540 11680 18780 11920
rect 18870 11680 19110 11920
rect 19200 11680 19440 11920
rect 19530 11680 19770 11920
rect 19860 11680 20100 11920
rect 8310 11350 8550 11590
rect 8640 11350 8880 11590
rect 8970 11350 9210 11590
rect 9300 11350 9540 11590
rect 9630 11350 9870 11590
rect 9960 11350 10200 11590
rect 10290 11350 10530 11590
rect 10620 11350 10860 11590
rect 10950 11350 11190 11590
rect 11280 11350 11520 11590
rect 11610 11350 11850 11590
rect 11940 11350 12180 11590
rect 12270 11350 12510 11590
rect 12600 11350 12840 11590
rect 12930 11350 13170 11590
rect 13260 11350 13500 11590
rect 13590 11350 13830 11590
rect 13920 11350 14160 11590
rect 14250 11350 14490 11590
rect 14580 11350 14820 11590
rect 14910 11350 15150 11590
rect 15240 11350 15480 11590
rect 15570 11350 15810 11590
rect 15900 11350 16140 11590
rect 16230 11350 16470 11590
rect 16560 11350 16800 11590
rect 16890 11350 17130 11590
rect 17220 11350 17460 11590
rect 17550 11350 17790 11590
rect 17880 11350 18120 11590
rect 18210 11350 18450 11590
rect 18540 11350 18780 11590
rect 18870 11350 19110 11590
rect 19200 11350 19440 11590
rect 19530 11350 19770 11590
rect 19860 11350 20100 11590
rect 8310 11020 8550 11260
rect 8640 11020 8880 11260
rect 8970 11020 9210 11260
rect 9300 11020 9540 11260
rect 9630 11020 9870 11260
rect 9960 11020 10200 11260
rect 10290 11020 10530 11260
rect 10620 11020 10860 11260
rect 10950 11020 11190 11260
rect 11280 11020 11520 11260
rect 11610 11020 11850 11260
rect 11940 11020 12180 11260
rect 12270 11020 12510 11260
rect 12600 11020 12840 11260
rect 12930 11020 13170 11260
rect 13260 11020 13500 11260
rect 13590 11020 13830 11260
rect 13920 11020 14160 11260
rect 14250 11020 14490 11260
rect 14580 11020 14820 11260
rect 14910 11020 15150 11260
rect 15240 11020 15480 11260
rect 15570 11020 15810 11260
rect 15900 11020 16140 11260
rect 16230 11020 16470 11260
rect 16560 11020 16800 11260
rect 16890 11020 17130 11260
rect 17220 11020 17460 11260
rect 17550 11020 17790 11260
rect 17880 11020 18120 11260
rect 18210 11020 18450 11260
rect 18540 11020 18780 11260
rect 18870 11020 19110 11260
rect 19200 11020 19440 11260
rect 19530 11020 19770 11260
rect 19860 11020 20100 11260
rect 8310 10690 8550 10930
rect 8640 10690 8880 10930
rect 8970 10690 9210 10930
rect 9300 10690 9540 10930
rect 9630 10690 9870 10930
rect 9960 10690 10200 10930
rect 10290 10690 10530 10930
rect 10620 10690 10860 10930
rect 10950 10690 11190 10930
rect 11280 10690 11520 10930
rect 11610 10690 11850 10930
rect 11940 10690 12180 10930
rect 12270 10690 12510 10930
rect 12600 10690 12840 10930
rect 12930 10690 13170 10930
rect 13260 10690 13500 10930
rect 13590 10690 13830 10930
rect 13920 10690 14160 10930
rect 14250 10690 14490 10930
rect 14580 10690 14820 10930
rect 14910 10690 15150 10930
rect 15240 10690 15480 10930
rect 15570 10690 15810 10930
rect 15900 10690 16140 10930
rect 16230 10690 16470 10930
rect 16560 10690 16800 10930
rect 16890 10690 17130 10930
rect 17220 10690 17460 10930
rect 17550 10690 17790 10930
rect 17880 10690 18120 10930
rect 18210 10690 18450 10930
rect 18540 10690 18780 10930
rect 18870 10690 19110 10930
rect 19200 10690 19440 10930
rect 19530 10690 19770 10930
rect 19860 10690 20100 10930
rect 8310 10360 8550 10600
rect 8640 10360 8880 10600
rect 8970 10360 9210 10600
rect 9300 10360 9540 10600
rect 9630 10360 9870 10600
rect 9960 10360 10200 10600
rect 10290 10360 10530 10600
rect 10620 10360 10860 10600
rect 10950 10360 11190 10600
rect 11280 10360 11520 10600
rect 11610 10360 11850 10600
rect 11940 10360 12180 10600
rect 12270 10360 12510 10600
rect 12600 10360 12840 10600
rect 12930 10360 13170 10600
rect 13260 10360 13500 10600
rect 13590 10360 13830 10600
rect 13920 10360 14160 10600
rect 14250 10360 14490 10600
rect 14580 10360 14820 10600
rect 14910 10360 15150 10600
rect 15240 10360 15480 10600
rect 15570 10360 15810 10600
rect 15900 10360 16140 10600
rect 16230 10360 16470 10600
rect 16560 10360 16800 10600
rect 16890 10360 17130 10600
rect 17220 10360 17460 10600
rect 17550 10360 17790 10600
rect 17880 10360 18120 10600
rect 18210 10360 18450 10600
rect 18540 10360 18780 10600
rect 18870 10360 19110 10600
rect 19200 10360 19440 10600
rect 19530 10360 19770 10600
rect 19860 10360 20100 10600
rect 8310 10030 8550 10270
rect 8640 10030 8880 10270
rect 8970 10030 9210 10270
rect 9300 10030 9540 10270
rect 9630 10030 9870 10270
rect 9960 10030 10200 10270
rect 10290 10030 10530 10270
rect 10620 10030 10860 10270
rect 10950 10030 11190 10270
rect 11280 10030 11520 10270
rect 11610 10030 11850 10270
rect 11940 10030 12180 10270
rect 12270 10030 12510 10270
rect 12600 10030 12840 10270
rect 12930 10030 13170 10270
rect 13260 10030 13500 10270
rect 13590 10030 13830 10270
rect 13920 10030 14160 10270
rect 14250 10030 14490 10270
rect 14580 10030 14820 10270
rect 14910 10030 15150 10270
rect 15240 10030 15480 10270
rect 15570 10030 15810 10270
rect 15900 10030 16140 10270
rect 16230 10030 16470 10270
rect 16560 10030 16800 10270
rect 16890 10030 17130 10270
rect 17220 10030 17460 10270
rect 17550 10030 17790 10270
rect 17880 10030 18120 10270
rect 18210 10030 18450 10270
rect 18540 10030 18780 10270
rect 18870 10030 19110 10270
rect 19200 10030 19440 10270
rect 19530 10030 19770 10270
rect 19860 10030 20100 10270
rect 8310 9700 8550 9940
rect 8640 9700 8880 9940
rect 8970 9700 9210 9940
rect 9300 9700 9540 9940
rect 9630 9700 9870 9940
rect 9960 9700 10200 9940
rect 10290 9700 10530 9940
rect 10620 9700 10860 9940
rect 10950 9700 11190 9940
rect 11280 9700 11520 9940
rect 11610 9700 11850 9940
rect 11940 9700 12180 9940
rect 12270 9700 12510 9940
rect 12600 9700 12840 9940
rect 12930 9700 13170 9940
rect 13260 9700 13500 9940
rect 13590 9700 13830 9940
rect 13920 9700 14160 9940
rect 14250 9700 14490 9940
rect 14580 9700 14820 9940
rect 14910 9700 15150 9940
rect 15240 9700 15480 9940
rect 15570 9700 15810 9940
rect 15900 9700 16140 9940
rect 16230 9700 16470 9940
rect 16560 9700 16800 9940
rect 16890 9700 17130 9940
rect 17220 9700 17460 9940
rect 17550 9700 17790 9940
rect 17880 9700 18120 9940
rect 18210 9700 18450 9940
rect 18540 9700 18780 9940
rect 18870 9700 19110 9940
rect 19200 9700 19440 9940
rect 19530 9700 19770 9940
rect 19860 9700 20100 9940
rect 8310 9370 8550 9610
rect 8640 9370 8880 9610
rect 8970 9370 9210 9610
rect 9300 9370 9540 9610
rect 9630 9370 9870 9610
rect 9960 9370 10200 9610
rect 10290 9370 10530 9610
rect 10620 9370 10860 9610
rect 10950 9370 11190 9610
rect 11280 9370 11520 9610
rect 11610 9370 11850 9610
rect 11940 9370 12180 9610
rect 12270 9370 12510 9610
rect 12600 9370 12840 9610
rect 12930 9370 13170 9610
rect 13260 9370 13500 9610
rect 13590 9370 13830 9610
rect 13920 9370 14160 9610
rect 14250 9370 14490 9610
rect 14580 9370 14820 9610
rect 14910 9370 15150 9610
rect 15240 9370 15480 9610
rect 15570 9370 15810 9610
rect 15900 9370 16140 9610
rect 16230 9370 16470 9610
rect 16560 9370 16800 9610
rect 16890 9370 17130 9610
rect 17220 9370 17460 9610
rect 17550 9370 17790 9610
rect 17880 9370 18120 9610
rect 18210 9370 18450 9610
rect 18540 9370 18780 9610
rect 18870 9370 19110 9610
rect 19200 9370 19440 9610
rect 19530 9370 19770 9610
rect 19860 9370 20100 9610
rect 8310 9040 8550 9280
rect 8640 9040 8880 9280
rect 8970 9040 9210 9280
rect 9300 9040 9540 9280
rect 9630 9040 9870 9280
rect 9960 9040 10200 9280
rect 10290 9040 10530 9280
rect 10620 9040 10860 9280
rect 10950 9040 11190 9280
rect 11280 9040 11520 9280
rect 11610 9040 11850 9280
rect 11940 9040 12180 9280
rect 12270 9040 12510 9280
rect 12600 9040 12840 9280
rect 12930 9040 13170 9280
rect 13260 9040 13500 9280
rect 13590 9040 13830 9280
rect 13920 9040 14160 9280
rect 14250 9040 14490 9280
rect 14580 9040 14820 9280
rect 14910 9040 15150 9280
rect 15240 9040 15480 9280
rect 15570 9040 15810 9280
rect 15900 9040 16140 9280
rect 16230 9040 16470 9280
rect 16560 9040 16800 9280
rect 16890 9040 17130 9280
rect 17220 9040 17460 9280
rect 17550 9040 17790 9280
rect 17880 9040 18120 9280
rect 18210 9040 18450 9280
rect 18540 9040 18780 9280
rect 18870 9040 19110 9280
rect 19200 9040 19440 9280
rect 19530 9040 19770 9280
rect 19860 9040 20100 9280
rect 31180 7590 31420 7830
rect 31510 7590 31750 7830
rect 31840 7590 32080 7830
rect 32170 7590 32410 7830
rect 32500 7590 32740 7830
rect 32830 7590 33070 7830
rect 33160 7590 33400 7830
rect 33490 7590 33730 7830
rect 33820 7590 34060 7830
rect 34150 7590 34390 7830
rect 34480 7590 34720 7830
rect 34810 7590 35050 7830
rect 35140 7590 35380 7830
rect 35470 7590 35710 7830
rect 35800 7590 36040 7830
rect 36130 7590 36370 7830
rect 36460 7590 36700 7830
rect 36790 7590 37030 7830
rect 37120 7590 37360 7830
rect 37450 7590 37690 7830
rect 31180 7260 31420 7500
rect 31510 7260 31750 7500
rect 31840 7260 32080 7500
rect 32170 7260 32410 7500
rect 32500 7260 32740 7500
rect 32830 7260 33070 7500
rect 33160 7260 33400 7500
rect 33490 7260 33730 7500
rect 33820 7260 34060 7500
rect 34150 7260 34390 7500
rect 34480 7260 34720 7500
rect 34810 7260 35050 7500
rect 35140 7260 35380 7500
rect 35470 7260 35710 7500
rect 35800 7260 36040 7500
rect 36130 7260 36370 7500
rect 36460 7260 36700 7500
rect 36790 7260 37030 7500
rect 37120 7260 37360 7500
rect 37450 7260 37690 7500
rect 31180 6930 31420 7170
rect 31510 6930 31750 7170
rect 31840 6930 32080 7170
rect 32170 6930 32410 7170
rect 32500 6930 32740 7170
rect 32830 6930 33070 7170
rect 33160 6930 33400 7170
rect 33490 6930 33730 7170
rect 33820 6930 34060 7170
rect 34150 6930 34390 7170
rect 34480 6930 34720 7170
rect 34810 6930 35050 7170
rect 35140 6930 35380 7170
rect 35470 6930 35710 7170
rect 35800 6930 36040 7170
rect 36130 6930 36370 7170
rect 36460 6930 36700 7170
rect 36790 6930 37030 7170
rect 37120 6930 37360 7170
rect 37450 6930 37690 7170
rect 31180 6600 31420 6840
rect 31510 6600 31750 6840
rect 31840 6600 32080 6840
rect 32170 6600 32410 6840
rect 32500 6600 32740 6840
rect 32830 6600 33070 6840
rect 33160 6600 33400 6840
rect 33490 6600 33730 6840
rect 33820 6600 34060 6840
rect 34150 6600 34390 6840
rect 34480 6600 34720 6840
rect 34810 6600 35050 6840
rect 35140 6600 35380 6840
rect 35470 6600 35710 6840
rect 35800 6600 36040 6840
rect 36130 6600 36370 6840
rect 36460 6600 36700 6840
rect 36790 6600 37030 6840
rect 37120 6600 37360 6840
rect 37450 6600 37690 6840
rect 31180 6270 31420 6510
rect 31510 6270 31750 6510
rect 31840 6270 32080 6510
rect 32170 6270 32410 6510
rect 32500 6270 32740 6510
rect 32830 6270 33070 6510
rect 33160 6270 33400 6510
rect 33490 6270 33730 6510
rect 33820 6270 34060 6510
rect 34150 6270 34390 6510
rect 34480 6270 34720 6510
rect 34810 6270 35050 6510
rect 35140 6270 35380 6510
rect 35470 6270 35710 6510
rect 35800 6270 36040 6510
rect 36130 6270 36370 6510
rect 36460 6270 36700 6510
rect 36790 6270 37030 6510
rect 37120 6270 37360 6510
rect 37450 6270 37690 6510
rect 31180 5940 31420 6180
rect 31510 5940 31750 6180
rect 31840 5940 32080 6180
rect 32170 5940 32410 6180
rect 32500 5940 32740 6180
rect 32830 5940 33070 6180
rect 33160 5940 33400 6180
rect 33490 5940 33730 6180
rect 33820 5940 34060 6180
rect 34150 5940 34390 6180
rect 34480 5940 34720 6180
rect 34810 5940 35050 6180
rect 35140 5940 35380 6180
rect 35470 5940 35710 6180
rect 35800 5940 36040 6180
rect 36130 5940 36370 6180
rect 36460 5940 36700 6180
rect 36790 5940 37030 6180
rect 37120 5940 37360 6180
rect 37450 5940 37690 6180
rect 31180 5610 31420 5850
rect 31510 5610 31750 5850
rect 31840 5610 32080 5850
rect 32170 5610 32410 5850
rect 32500 5610 32740 5850
rect 32830 5610 33070 5850
rect 33160 5610 33400 5850
rect 33490 5610 33730 5850
rect 33820 5610 34060 5850
rect 34150 5610 34390 5850
rect 34480 5610 34720 5850
rect 34810 5610 35050 5850
rect 35140 5610 35380 5850
rect 35470 5610 35710 5850
rect 35800 5610 36040 5850
rect 36130 5610 36370 5850
rect 36460 5610 36700 5850
rect 36790 5610 37030 5850
rect 37120 5610 37360 5850
rect 37450 5610 37690 5850
rect 31180 5280 31420 5520
rect 31510 5280 31750 5520
rect 31840 5280 32080 5520
rect 32170 5280 32410 5520
rect 32500 5280 32740 5520
rect 32830 5280 33070 5520
rect 33160 5280 33400 5520
rect 33490 5280 33730 5520
rect 33820 5280 34060 5520
rect 34150 5280 34390 5520
rect 34480 5280 34720 5520
rect 34810 5280 35050 5520
rect 35140 5280 35380 5520
rect 35470 5280 35710 5520
rect 35800 5280 36040 5520
rect 36130 5280 36370 5520
rect 36460 5280 36700 5520
rect 36790 5280 37030 5520
rect 37120 5280 37360 5520
rect 37450 5280 37690 5520
rect 31180 4950 31420 5190
rect 31510 4950 31750 5190
rect 31840 4950 32080 5190
rect 32170 4950 32410 5190
rect 32500 4950 32740 5190
rect 32830 4950 33070 5190
rect 33160 4950 33400 5190
rect 33490 4950 33730 5190
rect 33820 4950 34060 5190
rect 34150 4950 34390 5190
rect 34480 4950 34720 5190
rect 34810 4950 35050 5190
rect 35140 4950 35380 5190
rect 35470 4950 35710 5190
rect 35800 4950 36040 5190
rect 36130 4950 36370 5190
rect 36460 4950 36700 5190
rect 36790 4950 37030 5190
rect 37120 4950 37360 5190
rect 37450 4950 37690 5190
rect 31180 4620 31420 4860
rect 31510 4620 31750 4860
rect 31840 4620 32080 4860
rect 32170 4620 32410 4860
rect 32500 4620 32740 4860
rect 32830 4620 33070 4860
rect 33160 4620 33400 4860
rect 33490 4620 33730 4860
rect 33820 4620 34060 4860
rect 34150 4620 34390 4860
rect 34480 4620 34720 4860
rect 34810 4620 35050 4860
rect 35140 4620 35380 4860
rect 35470 4620 35710 4860
rect 35800 4620 36040 4860
rect 36130 4620 36370 4860
rect 36460 4620 36700 4860
rect 36790 4620 37030 4860
rect 37120 4620 37360 4860
rect 37450 4620 37690 4860
rect 31180 4290 31420 4530
rect 31510 4290 31750 4530
rect 31840 4290 32080 4530
rect 32170 4290 32410 4530
rect 32500 4290 32740 4530
rect 32830 4290 33070 4530
rect 33160 4290 33400 4530
rect 33490 4290 33730 4530
rect 33820 4290 34060 4530
rect 34150 4290 34390 4530
rect 34480 4290 34720 4530
rect 34810 4290 35050 4530
rect 35140 4290 35380 4530
rect 35470 4290 35710 4530
rect 35800 4290 36040 4530
rect 36130 4290 36370 4530
rect 36460 4290 36700 4530
rect 36790 4290 37030 4530
rect 37120 4290 37360 4530
rect 37450 4290 37690 4530
rect 31180 3960 31420 4200
rect 31510 3960 31750 4200
rect 31840 3960 32080 4200
rect 32170 3960 32410 4200
rect 32500 3960 32740 4200
rect 32830 3960 33070 4200
rect 33160 3960 33400 4200
rect 33490 3960 33730 4200
rect 33820 3960 34060 4200
rect 34150 3960 34390 4200
rect 34480 3960 34720 4200
rect 34810 3960 35050 4200
rect 35140 3960 35380 4200
rect 35470 3960 35710 4200
rect 35800 3960 36040 4200
rect 36130 3960 36370 4200
rect 36460 3960 36700 4200
rect 36790 3960 37030 4200
rect 37120 3960 37360 4200
rect 37450 3960 37690 4200
rect 31180 3630 31420 3870
rect 31510 3630 31750 3870
rect 31840 3630 32080 3870
rect 32170 3630 32410 3870
rect 32500 3630 32740 3870
rect 32830 3630 33070 3870
rect 33160 3630 33400 3870
rect 33490 3630 33730 3870
rect 33820 3630 34060 3870
rect 34150 3630 34390 3870
rect 34480 3630 34720 3870
rect 34810 3630 35050 3870
rect 35140 3630 35380 3870
rect 35470 3630 35710 3870
rect 35800 3630 36040 3870
rect 36130 3630 36370 3870
rect 36460 3630 36700 3870
rect 36790 3630 37030 3870
rect 37120 3630 37360 3870
rect 37450 3630 37690 3870
rect 31180 3300 31420 3540
rect 31510 3300 31750 3540
rect 31840 3300 32080 3540
rect 32170 3300 32410 3540
rect 32500 3300 32740 3540
rect 32830 3300 33070 3540
rect 33160 3300 33400 3540
rect 33490 3300 33730 3540
rect 33820 3300 34060 3540
rect 34150 3300 34390 3540
rect 34480 3300 34720 3540
rect 34810 3300 35050 3540
rect 35140 3300 35380 3540
rect 35470 3300 35710 3540
rect 35800 3300 36040 3540
rect 36130 3300 36370 3540
rect 36460 3300 36700 3540
rect 36790 3300 37030 3540
rect 37120 3300 37360 3540
rect 37450 3300 37690 3540
rect 31180 2970 31420 3210
rect 31510 2970 31750 3210
rect 31840 2970 32080 3210
rect 32170 2970 32410 3210
rect 32500 2970 32740 3210
rect 32830 2970 33070 3210
rect 33160 2970 33400 3210
rect 33490 2970 33730 3210
rect 33820 2970 34060 3210
rect 34150 2970 34390 3210
rect 34480 2970 34720 3210
rect 34810 2970 35050 3210
rect 35140 2970 35380 3210
rect 35470 2970 35710 3210
rect 35800 2970 36040 3210
rect 36130 2970 36370 3210
rect 36460 2970 36700 3210
rect 36790 2970 37030 3210
rect 37120 2970 37360 3210
rect 37450 2970 37690 3210
rect 31180 2640 31420 2880
rect 31510 2640 31750 2880
rect 31840 2640 32080 2880
rect 32170 2640 32410 2880
rect 32500 2640 32740 2880
rect 32830 2640 33070 2880
rect 33160 2640 33400 2880
rect 33490 2640 33730 2880
rect 33820 2640 34060 2880
rect 34150 2640 34390 2880
rect 34480 2640 34720 2880
rect 34810 2640 35050 2880
rect 35140 2640 35380 2880
rect 35470 2640 35710 2880
rect 35800 2640 36040 2880
rect 36130 2640 36370 2880
rect 36460 2640 36700 2880
rect 36790 2640 37030 2880
rect 37120 2640 37360 2880
rect 37450 2640 37690 2880
rect 31180 2310 31420 2550
rect 31510 2310 31750 2550
rect 31840 2310 32080 2550
rect 32170 2310 32410 2550
rect 32500 2310 32740 2550
rect 32830 2310 33070 2550
rect 33160 2310 33400 2550
rect 33490 2310 33730 2550
rect 33820 2310 34060 2550
rect 34150 2310 34390 2550
rect 34480 2310 34720 2550
rect 34810 2310 35050 2550
rect 35140 2310 35380 2550
rect 35470 2310 35710 2550
rect 35800 2310 36040 2550
rect 36130 2310 36370 2550
rect 36460 2310 36700 2550
rect 36790 2310 37030 2550
rect 37120 2310 37360 2550
rect 37450 2310 37690 2550
rect 31180 1980 31420 2220
rect 31510 1980 31750 2220
rect 31840 1980 32080 2220
rect 32170 1980 32410 2220
rect 32500 1980 32740 2220
rect 32830 1980 33070 2220
rect 33160 1980 33400 2220
rect 33490 1980 33730 2220
rect 33820 1980 34060 2220
rect 34150 1980 34390 2220
rect 34480 1980 34720 2220
rect 34810 1980 35050 2220
rect 35140 1980 35380 2220
rect 35470 1980 35710 2220
rect 35800 1980 36040 2220
rect 36130 1980 36370 2220
rect 36460 1980 36700 2220
rect 36790 1980 37030 2220
rect 37120 1980 37360 2220
rect 37450 1980 37690 2220
rect 31180 1650 31420 1890
rect 31510 1650 31750 1890
rect 31840 1650 32080 1890
rect 32170 1650 32410 1890
rect 32500 1650 32740 1890
rect 32830 1650 33070 1890
rect 33160 1650 33400 1890
rect 33490 1650 33730 1890
rect 33820 1650 34060 1890
rect 34150 1650 34390 1890
rect 34480 1650 34720 1890
rect 34810 1650 35050 1890
rect 35140 1650 35380 1890
rect 35470 1650 35710 1890
rect 35800 1650 36040 1890
rect 36130 1650 36370 1890
rect 36460 1650 36700 1890
rect 36790 1650 37030 1890
rect 37120 1650 37360 1890
rect 37450 1650 37690 1890
rect 31180 1320 31420 1560
rect 31510 1320 31750 1560
rect 31840 1320 32080 1560
rect 32170 1320 32410 1560
rect 32500 1320 32740 1560
rect 32830 1320 33070 1560
rect 33160 1320 33400 1560
rect 33490 1320 33730 1560
rect 33820 1320 34060 1560
rect 34150 1320 34390 1560
rect 34480 1320 34720 1560
rect 34810 1320 35050 1560
rect 35140 1320 35380 1560
rect 35470 1320 35710 1560
rect 35800 1320 36040 1560
rect 36130 1320 36370 1560
rect 36460 1320 36700 1560
rect 36790 1320 37030 1560
rect 37120 1320 37360 1560
rect 37450 1320 37690 1560
rect 31180 -10 31420 230
rect 31510 -10 31750 230
rect 31840 -10 32080 230
rect 32170 -10 32410 230
rect 32500 -10 32740 230
rect 32830 -10 33070 230
rect 33160 -10 33400 230
rect 33490 -10 33730 230
rect 33820 -10 34060 230
rect 34150 -10 34390 230
rect 34480 -10 34720 230
rect 34810 -10 35050 230
rect 35140 -10 35380 230
rect 35470 -10 35710 230
rect 35800 -10 36040 230
rect 36130 -10 36370 230
rect 36460 -10 36700 230
rect 36790 -10 37030 230
rect 37120 -10 37360 230
rect 37450 -10 37690 230
rect 31180 -340 31420 -100
rect 31510 -340 31750 -100
rect 31840 -340 32080 -100
rect 32170 -340 32410 -100
rect 32500 -340 32740 -100
rect 32830 -340 33070 -100
rect 33160 -340 33400 -100
rect 33490 -340 33730 -100
rect 33820 -340 34060 -100
rect 34150 -340 34390 -100
rect 34480 -340 34720 -100
rect 34810 -340 35050 -100
rect 35140 -340 35380 -100
rect 35470 -340 35710 -100
rect 35800 -340 36040 -100
rect 36130 -340 36370 -100
rect 36460 -340 36700 -100
rect 36790 -340 37030 -100
rect 37120 -340 37360 -100
rect 37450 -340 37690 -100
rect 31180 -670 31420 -430
rect 31510 -670 31750 -430
rect 31840 -670 32080 -430
rect 32170 -670 32410 -430
rect 32500 -670 32740 -430
rect 32830 -670 33070 -430
rect 33160 -670 33400 -430
rect 33490 -670 33730 -430
rect 33820 -670 34060 -430
rect 34150 -670 34390 -430
rect 34480 -670 34720 -430
rect 34810 -670 35050 -430
rect 35140 -670 35380 -430
rect 35470 -670 35710 -430
rect 35800 -670 36040 -430
rect 36130 -670 36370 -430
rect 36460 -670 36700 -430
rect 36790 -670 37030 -430
rect 37120 -670 37360 -430
rect 37450 -670 37690 -430
rect 31180 -1000 31420 -760
rect 31510 -1000 31750 -760
rect 31840 -1000 32080 -760
rect 32170 -1000 32410 -760
rect 32500 -1000 32740 -760
rect 32830 -1000 33070 -760
rect 33160 -1000 33400 -760
rect 33490 -1000 33730 -760
rect 33820 -1000 34060 -760
rect 34150 -1000 34390 -760
rect 34480 -1000 34720 -760
rect 34810 -1000 35050 -760
rect 35140 -1000 35380 -760
rect 35470 -1000 35710 -760
rect 35800 -1000 36040 -760
rect 36130 -1000 36370 -760
rect 36460 -1000 36700 -760
rect 36790 -1000 37030 -760
rect 37120 -1000 37360 -760
rect 37450 -1000 37690 -760
rect 31180 -1330 31420 -1090
rect 31510 -1330 31750 -1090
rect 31840 -1330 32080 -1090
rect 32170 -1330 32410 -1090
rect 32500 -1330 32740 -1090
rect 32830 -1330 33070 -1090
rect 33160 -1330 33400 -1090
rect 33490 -1330 33730 -1090
rect 33820 -1330 34060 -1090
rect 34150 -1330 34390 -1090
rect 34480 -1330 34720 -1090
rect 34810 -1330 35050 -1090
rect 35140 -1330 35380 -1090
rect 35470 -1330 35710 -1090
rect 35800 -1330 36040 -1090
rect 36130 -1330 36370 -1090
rect 36460 -1330 36700 -1090
rect 36790 -1330 37030 -1090
rect 37120 -1330 37360 -1090
rect 37450 -1330 37690 -1090
rect 31180 -1660 31420 -1420
rect 31510 -1660 31750 -1420
rect 31840 -1660 32080 -1420
rect 32170 -1660 32410 -1420
rect 32500 -1660 32740 -1420
rect 32830 -1660 33070 -1420
rect 33160 -1660 33400 -1420
rect 33490 -1660 33730 -1420
rect 33820 -1660 34060 -1420
rect 34150 -1660 34390 -1420
rect 34480 -1660 34720 -1420
rect 34810 -1660 35050 -1420
rect 35140 -1660 35380 -1420
rect 35470 -1660 35710 -1420
rect 35800 -1660 36040 -1420
rect 36130 -1660 36370 -1420
rect 36460 -1660 36700 -1420
rect 36790 -1660 37030 -1420
rect 37120 -1660 37360 -1420
rect 37450 -1660 37690 -1420
rect 31180 -1990 31420 -1750
rect 31510 -1990 31750 -1750
rect 31840 -1990 32080 -1750
rect 32170 -1990 32410 -1750
rect 32500 -1990 32740 -1750
rect 32830 -1990 33070 -1750
rect 33160 -1990 33400 -1750
rect 33490 -1990 33730 -1750
rect 33820 -1990 34060 -1750
rect 34150 -1990 34390 -1750
rect 34480 -1990 34720 -1750
rect 34810 -1990 35050 -1750
rect 35140 -1990 35380 -1750
rect 35470 -1990 35710 -1750
rect 35800 -1990 36040 -1750
rect 36130 -1990 36370 -1750
rect 36460 -1990 36700 -1750
rect 36790 -1990 37030 -1750
rect 37120 -1990 37360 -1750
rect 37450 -1990 37690 -1750
rect 31180 -2320 31420 -2080
rect 31510 -2320 31750 -2080
rect 31840 -2320 32080 -2080
rect 32170 -2320 32410 -2080
rect 32500 -2320 32740 -2080
rect 32830 -2320 33070 -2080
rect 33160 -2320 33400 -2080
rect 33490 -2320 33730 -2080
rect 33820 -2320 34060 -2080
rect 34150 -2320 34390 -2080
rect 34480 -2320 34720 -2080
rect 34810 -2320 35050 -2080
rect 35140 -2320 35380 -2080
rect 35470 -2320 35710 -2080
rect 35800 -2320 36040 -2080
rect 36130 -2320 36370 -2080
rect 36460 -2320 36700 -2080
rect 36790 -2320 37030 -2080
rect 37120 -2320 37360 -2080
rect 37450 -2320 37690 -2080
rect 31180 -2650 31420 -2410
rect 31510 -2650 31750 -2410
rect 31840 -2650 32080 -2410
rect 32170 -2650 32410 -2410
rect 32500 -2650 32740 -2410
rect 32830 -2650 33070 -2410
rect 33160 -2650 33400 -2410
rect 33490 -2650 33730 -2410
rect 33820 -2650 34060 -2410
rect 34150 -2650 34390 -2410
rect 34480 -2650 34720 -2410
rect 34810 -2650 35050 -2410
rect 35140 -2650 35380 -2410
rect 35470 -2650 35710 -2410
rect 35800 -2650 36040 -2410
rect 36130 -2650 36370 -2410
rect 36460 -2650 36700 -2410
rect 36790 -2650 37030 -2410
rect 37120 -2650 37360 -2410
rect 37450 -2650 37690 -2410
rect 31180 -2980 31420 -2740
rect 31510 -2980 31750 -2740
rect 31840 -2980 32080 -2740
rect 32170 -2980 32410 -2740
rect 32500 -2980 32740 -2740
rect 32830 -2980 33070 -2740
rect 33160 -2980 33400 -2740
rect 33490 -2980 33730 -2740
rect 33820 -2980 34060 -2740
rect 34150 -2980 34390 -2740
rect 34480 -2980 34720 -2740
rect 34810 -2980 35050 -2740
rect 35140 -2980 35380 -2740
rect 35470 -2980 35710 -2740
rect 35800 -2980 36040 -2740
rect 36130 -2980 36370 -2740
rect 36460 -2980 36700 -2740
rect 36790 -2980 37030 -2740
rect 37120 -2980 37360 -2740
rect 37450 -2980 37690 -2740
rect 31180 -3310 31420 -3070
rect 31510 -3310 31750 -3070
rect 31840 -3310 32080 -3070
rect 32170 -3310 32410 -3070
rect 32500 -3310 32740 -3070
rect 32830 -3310 33070 -3070
rect 33160 -3310 33400 -3070
rect 33490 -3310 33730 -3070
rect 33820 -3310 34060 -3070
rect 34150 -3310 34390 -3070
rect 34480 -3310 34720 -3070
rect 34810 -3310 35050 -3070
rect 35140 -3310 35380 -3070
rect 35470 -3310 35710 -3070
rect 35800 -3310 36040 -3070
rect 36130 -3310 36370 -3070
rect 36460 -3310 36700 -3070
rect 36790 -3310 37030 -3070
rect 37120 -3310 37360 -3070
rect 37450 -3310 37690 -3070
rect 31180 -3640 31420 -3400
rect 31510 -3640 31750 -3400
rect 31840 -3640 32080 -3400
rect 32170 -3640 32410 -3400
rect 32500 -3640 32740 -3400
rect 32830 -3640 33070 -3400
rect 33160 -3640 33400 -3400
rect 33490 -3640 33730 -3400
rect 33820 -3640 34060 -3400
rect 34150 -3640 34390 -3400
rect 34480 -3640 34720 -3400
rect 34810 -3640 35050 -3400
rect 35140 -3640 35380 -3400
rect 35470 -3640 35710 -3400
rect 35800 -3640 36040 -3400
rect 36130 -3640 36370 -3400
rect 36460 -3640 36700 -3400
rect 36790 -3640 37030 -3400
rect 37120 -3640 37360 -3400
rect 37450 -3640 37690 -3400
rect 31180 -3970 31420 -3730
rect 31510 -3970 31750 -3730
rect 31840 -3970 32080 -3730
rect 32170 -3970 32410 -3730
rect 32500 -3970 32740 -3730
rect 32830 -3970 33070 -3730
rect 33160 -3970 33400 -3730
rect 33490 -3970 33730 -3730
rect 33820 -3970 34060 -3730
rect 34150 -3970 34390 -3730
rect 34480 -3970 34720 -3730
rect 34810 -3970 35050 -3730
rect 35140 -3970 35380 -3730
rect 35470 -3970 35710 -3730
rect 35800 -3970 36040 -3730
rect 36130 -3970 36370 -3730
rect 36460 -3970 36700 -3730
rect 36790 -3970 37030 -3730
rect 37120 -3970 37360 -3730
rect 37450 -3970 37690 -3730
rect 31180 -4300 31420 -4060
rect 31510 -4300 31750 -4060
rect 31840 -4300 32080 -4060
rect 32170 -4300 32410 -4060
rect 32500 -4300 32740 -4060
rect 32830 -4300 33070 -4060
rect 33160 -4300 33400 -4060
rect 33490 -4300 33730 -4060
rect 33820 -4300 34060 -4060
rect 34150 -4300 34390 -4060
rect 34480 -4300 34720 -4060
rect 34810 -4300 35050 -4060
rect 35140 -4300 35380 -4060
rect 35470 -4300 35710 -4060
rect 35800 -4300 36040 -4060
rect 36130 -4300 36370 -4060
rect 36460 -4300 36700 -4060
rect 36790 -4300 37030 -4060
rect 37120 -4300 37360 -4060
rect 37450 -4300 37690 -4060
rect 31180 -4630 31420 -4390
rect 31510 -4630 31750 -4390
rect 31840 -4630 32080 -4390
rect 32170 -4630 32410 -4390
rect 32500 -4630 32740 -4390
rect 32830 -4630 33070 -4390
rect 33160 -4630 33400 -4390
rect 33490 -4630 33730 -4390
rect 33820 -4630 34060 -4390
rect 34150 -4630 34390 -4390
rect 34480 -4630 34720 -4390
rect 34810 -4630 35050 -4390
rect 35140 -4630 35380 -4390
rect 35470 -4630 35710 -4390
rect 35800 -4630 36040 -4390
rect 36130 -4630 36370 -4390
rect 36460 -4630 36700 -4390
rect 36790 -4630 37030 -4390
rect 37120 -4630 37360 -4390
rect 37450 -4630 37690 -4390
rect -1180 -5080 -940 -4840
rect -850 -5080 -610 -4840
rect -520 -5080 -280 -4840
rect -190 -5080 50 -4840
rect -1180 -5410 -940 -5170
rect -850 -5410 -610 -5170
rect -520 -5410 -280 -5170
rect -190 -5410 50 -5170
rect -1180 -5740 -940 -5500
rect -850 -5740 -610 -5500
rect -520 -5740 -280 -5500
rect -190 -5740 50 -5500
rect -1180 -6070 -940 -5830
rect -850 -6070 -610 -5830
rect -520 -6070 -280 -5830
rect -190 -6070 50 -5830
rect 14730 -5080 14970 -4840
rect 15060 -5080 15300 -4840
rect 15390 -5080 15630 -4840
rect 15720 -5080 15960 -4840
rect 14730 -5410 14970 -5170
rect 15060 -5410 15300 -5170
rect 15390 -5410 15630 -5170
rect 15720 -5410 15960 -5170
rect 14730 -5740 14970 -5500
rect 15060 -5740 15300 -5500
rect 15390 -5740 15630 -5500
rect 15720 -5740 15960 -5500
rect 14730 -6070 14970 -5830
rect 15060 -6070 15300 -5830
rect 15390 -6070 15630 -5830
rect 15720 -6070 15960 -5830
rect 31180 -4960 31420 -4720
rect 31510 -4960 31750 -4720
rect 31840 -4960 32080 -4720
rect 32170 -4960 32410 -4720
rect 32500 -4960 32740 -4720
rect 32830 -4960 33070 -4720
rect 33160 -4960 33400 -4720
rect 33490 -4960 33730 -4720
rect 33820 -4960 34060 -4720
rect 34150 -4960 34390 -4720
rect 34480 -4960 34720 -4720
rect 34810 -4960 35050 -4720
rect 35140 -4960 35380 -4720
rect 35470 -4960 35710 -4720
rect 35800 -4960 36040 -4720
rect 36130 -4960 36370 -4720
rect 36460 -4960 36700 -4720
rect 36790 -4960 37030 -4720
rect 37120 -4960 37360 -4720
rect 37450 -4960 37690 -4720
rect 31180 -5290 31420 -5050
rect 31510 -5290 31750 -5050
rect 31840 -5290 32080 -5050
rect 32170 -5290 32410 -5050
rect 32500 -5290 32740 -5050
rect 32830 -5290 33070 -5050
rect 33160 -5290 33400 -5050
rect 33490 -5290 33730 -5050
rect 33820 -5290 34060 -5050
rect 34150 -5290 34390 -5050
rect 34480 -5290 34720 -5050
rect 34810 -5290 35050 -5050
rect 35140 -5290 35380 -5050
rect 35470 -5290 35710 -5050
rect 35800 -5290 36040 -5050
rect 36130 -5290 36370 -5050
rect 36460 -5290 36700 -5050
rect 36790 -5290 37030 -5050
rect 37120 -5290 37360 -5050
rect 37450 -5290 37690 -5050
rect 31180 -5620 31420 -5380
rect 31510 -5620 31750 -5380
rect 31840 -5620 32080 -5380
rect 32170 -5620 32410 -5380
rect 32500 -5620 32740 -5380
rect 32830 -5620 33070 -5380
rect 33160 -5620 33400 -5380
rect 33490 -5620 33730 -5380
rect 33820 -5620 34060 -5380
rect 34150 -5620 34390 -5380
rect 34480 -5620 34720 -5380
rect 34810 -5620 35050 -5380
rect 35140 -5620 35380 -5380
rect 35470 -5620 35710 -5380
rect 35800 -5620 36040 -5380
rect 36130 -5620 36370 -5380
rect 36460 -5620 36700 -5380
rect 36790 -5620 37030 -5380
rect 37120 -5620 37360 -5380
rect 37450 -5620 37690 -5380
rect 31180 -5950 31420 -5710
rect 31510 -5950 31750 -5710
rect 31840 -5950 32080 -5710
rect 32170 -5950 32410 -5710
rect 32500 -5950 32740 -5710
rect 32830 -5950 33070 -5710
rect 33160 -5950 33400 -5710
rect 33490 -5950 33730 -5710
rect 33820 -5950 34060 -5710
rect 34150 -5950 34390 -5710
rect 34480 -5950 34720 -5710
rect 34810 -5950 35050 -5710
rect 35140 -5950 35380 -5710
rect 35470 -5950 35710 -5710
rect 35800 -5950 36040 -5710
rect 36130 -5950 36370 -5710
rect 36460 -5950 36700 -5710
rect 36790 -5950 37030 -5710
rect 37120 -5950 37360 -5710
rect 37450 -5950 37690 -5710
rect 31180 -6280 31420 -6040
rect 31510 -6280 31750 -6040
rect 31840 -6280 32080 -6040
rect 32170 -6280 32410 -6040
rect 32500 -6280 32740 -6040
rect 32830 -6280 33070 -6040
rect 33160 -6280 33400 -6040
rect 33490 -6280 33730 -6040
rect 33820 -6280 34060 -6040
rect 34150 -6280 34390 -6040
rect 34480 -6280 34720 -6040
rect 34810 -6280 35050 -6040
rect 35140 -6280 35380 -6040
rect 35470 -6280 35710 -6040
rect 35800 -6280 36040 -6040
rect 36130 -6280 36370 -6040
rect 36460 -6280 36700 -6040
rect 36790 -6280 37030 -6040
rect 37120 -6280 37360 -6040
rect 37450 -6280 37690 -6040
<< metal4 >>
rect -5550 21610 6760 21640
rect -5550 21580 -5180 21610
rect -4940 21580 -4850 21610
rect -4610 21580 -4520 21610
rect -4280 21580 -4190 21610
rect -3950 21580 -3860 21610
rect -3620 21580 -3530 21610
rect -3290 21580 -3200 21610
rect -2960 21580 -2870 21610
rect -2630 21580 -2540 21610
rect -2300 21580 -2170 21610
rect -1930 21580 -1840 21610
rect -1600 21580 -1510 21610
rect -1270 21580 -1180 21610
rect -940 21580 -850 21610
rect -610 21580 -520 21610
rect -280 21580 -190 21610
rect 50 21580 140 21610
rect 380 21580 470 21610
rect 710 21580 840 21610
rect 1080 21580 1170 21610
rect 1410 21580 1500 21610
rect 1740 21580 1830 21610
rect 2070 21580 2160 21610
rect 2400 21580 2490 21610
rect 2730 21580 2820 21610
rect 3060 21580 3150 21610
rect 3390 21580 3480 21610
rect 3720 21580 3850 21610
rect 4090 21580 4180 21610
rect 4420 21580 4510 21610
rect 4750 21580 4840 21610
rect 5080 21580 5170 21610
rect 5410 21580 5500 21610
rect 5740 21580 5830 21610
rect 6070 21580 6160 21610
rect 6400 21580 6490 21610
rect -5550 21510 -5260 21580
rect -5190 21510 -5180 21580
rect -4920 21510 -4900 21580
rect -4560 21510 -4540 21580
rect -4280 21510 -4270 21580
rect -4200 21510 -4190 21580
rect -3930 21510 -3910 21580
rect -3570 21510 -3550 21580
rect -3290 21510 -3280 21580
rect -3210 21510 -3200 21580
rect -2940 21510 -2920 21580
rect -2580 21510 -2560 21580
rect -2300 21510 -2250 21580
rect -2180 21510 -2170 21580
rect -1910 21510 -1890 21580
rect -1550 21510 -1530 21580
rect -1270 21510 -1260 21580
rect -1190 21510 -1180 21580
rect -920 21510 -900 21580
rect -560 21510 -540 21580
rect -280 21510 -270 21580
rect -200 21510 -190 21580
rect 70 21510 90 21580
rect 430 21510 450 21580
rect 710 21510 760 21580
rect 830 21510 840 21580
rect 1100 21510 1120 21580
rect 1460 21510 1480 21580
rect 1740 21510 1750 21580
rect 1820 21510 1830 21580
rect 2090 21510 2110 21580
rect 2450 21510 2470 21580
rect 2730 21510 2740 21580
rect 2810 21510 2820 21580
rect 3080 21510 3100 21580
rect 3440 21510 3460 21580
rect 3720 21510 3770 21580
rect 3840 21510 3850 21580
rect 4110 21510 4130 21580
rect 4470 21510 4490 21580
rect 4750 21510 4760 21580
rect 4830 21510 4840 21580
rect 5100 21510 5120 21580
rect 5460 21510 5480 21580
rect 5740 21510 5750 21580
rect 5820 21510 5830 21580
rect 6090 21510 6110 21580
rect 6450 21510 6470 21580
rect -5550 21490 -5180 21510
rect -4940 21490 -4850 21510
rect -4610 21490 -4520 21510
rect -4280 21490 -4190 21510
rect -3950 21490 -3860 21510
rect -3620 21490 -3530 21510
rect -3290 21490 -3200 21510
rect -2960 21490 -2870 21510
rect -2630 21490 -2540 21510
rect -2300 21490 -2170 21510
rect -1930 21490 -1840 21510
rect -1600 21490 -1510 21510
rect -1270 21490 -1180 21510
rect -940 21490 -850 21510
rect -610 21490 -520 21510
rect -280 21490 -190 21510
rect 50 21490 140 21510
rect 380 21490 470 21510
rect 710 21490 840 21510
rect 1080 21490 1170 21510
rect 1410 21490 1500 21510
rect 1740 21490 1830 21510
rect 2070 21490 2160 21510
rect 2400 21490 2490 21510
rect 2730 21490 2820 21510
rect 3060 21490 3150 21510
rect 3390 21490 3480 21510
rect 3720 21490 3850 21510
rect 4090 21490 4180 21510
rect 4420 21490 4510 21510
rect 4750 21490 4840 21510
rect 5080 21490 5170 21510
rect 5410 21490 5500 21510
rect 5740 21490 5830 21510
rect 6070 21490 6160 21510
rect 6400 21490 6490 21510
rect -5550 21420 -5260 21490
rect -5190 21420 -5180 21490
rect -4920 21420 -4900 21490
rect -4560 21420 -4540 21490
rect -4280 21420 -4270 21490
rect -4200 21420 -4190 21490
rect -3930 21420 -3910 21490
rect -3570 21420 -3550 21490
rect -3290 21420 -3280 21490
rect -3210 21420 -3200 21490
rect -2940 21420 -2920 21490
rect -2580 21420 -2560 21490
rect -2300 21420 -2250 21490
rect -2180 21420 -2170 21490
rect -1910 21420 -1890 21490
rect -1550 21420 -1530 21490
rect -1270 21420 -1260 21490
rect -1190 21420 -1180 21490
rect -920 21420 -900 21490
rect -560 21420 -540 21490
rect -280 21420 -270 21490
rect -200 21420 -190 21490
rect 70 21420 90 21490
rect 430 21420 450 21490
rect 710 21420 760 21490
rect 830 21420 840 21490
rect 1100 21420 1120 21490
rect 1460 21420 1480 21490
rect 1740 21420 1750 21490
rect 1820 21420 1830 21490
rect 2090 21420 2110 21490
rect 2450 21420 2470 21490
rect 2730 21420 2740 21490
rect 2810 21420 2820 21490
rect 3080 21420 3100 21490
rect 3440 21420 3460 21490
rect 3720 21420 3770 21490
rect 3840 21420 3850 21490
rect 4110 21420 4130 21490
rect 4470 21420 4490 21490
rect 4750 21420 4760 21490
rect 4830 21420 4840 21490
rect 5100 21420 5120 21490
rect 5460 21420 5480 21490
rect 5740 21420 5750 21490
rect 5820 21420 5830 21490
rect 6090 21420 6110 21490
rect 6450 21420 6470 21490
rect -5550 21400 -5180 21420
rect -4940 21400 -4850 21420
rect -4610 21400 -4520 21420
rect -4280 21400 -4190 21420
rect -3950 21400 -3860 21420
rect -3620 21400 -3530 21420
rect -3290 21400 -3200 21420
rect -2960 21400 -2870 21420
rect -2630 21400 -2540 21420
rect -2300 21400 -2170 21420
rect -1930 21400 -1840 21420
rect -1600 21400 -1510 21420
rect -1270 21400 -1180 21420
rect -940 21400 -850 21420
rect -610 21400 -520 21420
rect -280 21400 -190 21420
rect 50 21400 140 21420
rect 380 21400 470 21420
rect 710 21400 840 21420
rect 1080 21400 1170 21420
rect 1410 21400 1500 21420
rect 1740 21400 1830 21420
rect 2070 21400 2160 21420
rect 2400 21400 2490 21420
rect 2730 21400 2820 21420
rect 3060 21400 3150 21420
rect 3390 21400 3480 21420
rect 3720 21400 3850 21420
rect 4090 21400 4180 21420
rect 4420 21400 4510 21420
rect 4750 21400 4840 21420
rect 5080 21400 5170 21420
rect 5410 21400 5500 21420
rect 5740 21400 5830 21420
rect 6070 21400 6160 21420
rect 6400 21400 6490 21420
rect -5550 21330 -5260 21400
rect -5190 21370 -5180 21400
rect -5190 21330 -5170 21370
rect -5100 21330 -5080 21370
rect -5010 21330 -4990 21370
rect -4920 21330 -4900 21400
rect -4830 21330 -4810 21370
rect -4740 21330 -4720 21370
rect -4650 21330 -4630 21370
rect -4560 21330 -4540 21400
rect -4280 21370 -4270 21400
rect -4470 21330 -4450 21370
rect -4380 21330 -4360 21370
rect -4290 21330 -4270 21370
rect -4200 21370 -4190 21400
rect -4200 21330 -4180 21370
rect -4110 21330 -4090 21370
rect -4020 21330 -4000 21370
rect -3930 21330 -3910 21400
rect -3840 21330 -3820 21370
rect -3750 21330 -3730 21370
rect -3660 21330 -3640 21370
rect -3570 21330 -3550 21400
rect -3290 21370 -3280 21400
rect -3480 21330 -3460 21370
rect -3390 21330 -3370 21370
rect -3300 21330 -3280 21370
rect -3210 21370 -3200 21400
rect -3210 21330 -3190 21370
rect -3120 21330 -3100 21370
rect -3030 21330 -3010 21370
rect -2940 21330 -2920 21400
rect -2850 21330 -2830 21370
rect -2760 21330 -2740 21370
rect -2670 21330 -2650 21370
rect -2580 21330 -2560 21400
rect -2300 21370 -2250 21400
rect -2490 21330 -2470 21370
rect -2400 21330 -2380 21370
rect -2310 21330 -2250 21370
rect -2180 21370 -2170 21400
rect -2180 21330 -2160 21370
rect -2090 21330 -2070 21370
rect -2000 21330 -1980 21370
rect -1910 21330 -1890 21400
rect -1820 21330 -1800 21370
rect -1730 21330 -1710 21370
rect -1640 21330 -1620 21370
rect -1550 21330 -1530 21400
rect -1270 21370 -1260 21400
rect -1460 21330 -1440 21370
rect -1370 21330 -1350 21370
rect -1280 21330 -1260 21370
rect -1190 21370 -1180 21400
rect -1190 21330 -1170 21370
rect -1100 21330 -1080 21370
rect -1010 21330 -990 21370
rect -920 21330 -900 21400
rect -830 21330 -810 21370
rect -740 21330 -720 21370
rect -650 21330 -630 21370
rect -560 21330 -540 21400
rect -280 21370 -270 21400
rect -470 21330 -450 21370
rect -380 21330 -360 21370
rect -290 21330 -270 21370
rect -200 21370 -190 21400
rect -200 21330 -180 21370
rect -110 21330 -90 21370
rect -20 21330 0 21370
rect 70 21330 90 21400
rect 160 21330 180 21370
rect 250 21330 270 21370
rect 340 21330 360 21370
rect 430 21330 450 21400
rect 710 21370 760 21400
rect 520 21330 540 21370
rect 610 21330 630 21370
rect 700 21330 760 21370
rect 830 21370 840 21400
rect 830 21330 850 21370
rect 920 21330 940 21370
rect 1010 21330 1030 21370
rect 1100 21330 1120 21400
rect 1190 21330 1210 21370
rect 1280 21330 1300 21370
rect 1370 21330 1390 21370
rect 1460 21330 1480 21400
rect 1740 21370 1750 21400
rect 1550 21330 1570 21370
rect 1640 21330 1660 21370
rect 1730 21330 1750 21370
rect 1820 21370 1830 21400
rect 1820 21330 1840 21370
rect 1910 21330 1930 21370
rect 2000 21330 2020 21370
rect 2090 21330 2110 21400
rect 2180 21330 2200 21370
rect 2270 21330 2290 21370
rect 2360 21330 2380 21370
rect 2450 21330 2470 21400
rect 2730 21370 2740 21400
rect 2540 21330 2560 21370
rect 2630 21330 2650 21370
rect 2720 21330 2740 21370
rect 2810 21370 2820 21400
rect 2810 21330 2830 21370
rect 2900 21330 2920 21370
rect 2990 21330 3010 21370
rect 3080 21330 3100 21400
rect 3170 21330 3190 21370
rect 3260 21330 3280 21370
rect 3350 21330 3370 21370
rect 3440 21330 3460 21400
rect 3720 21370 3770 21400
rect 3530 21330 3550 21370
rect 3620 21330 3640 21370
rect 3710 21330 3770 21370
rect 3840 21370 3850 21400
rect 3840 21330 3860 21370
rect 3930 21330 3950 21370
rect 4020 21330 4040 21370
rect 4110 21330 4130 21400
rect 4200 21330 4220 21370
rect 4290 21330 4310 21370
rect 4380 21330 4400 21370
rect 4470 21330 4490 21400
rect 4750 21370 4760 21400
rect 4560 21330 4580 21370
rect 4650 21330 4670 21370
rect 4740 21330 4760 21370
rect 4830 21370 4840 21400
rect 4830 21330 4850 21370
rect 4920 21330 4940 21370
rect 5010 21330 5030 21370
rect 5100 21330 5120 21400
rect 5190 21330 5210 21370
rect 5280 21330 5300 21370
rect 5370 21330 5390 21370
rect 5460 21330 5480 21400
rect 5740 21370 5750 21400
rect 5550 21330 5570 21370
rect 5640 21330 5660 21370
rect 5730 21330 5750 21370
rect 5820 21370 5830 21400
rect 5820 21330 5840 21370
rect 5910 21330 5930 21370
rect 6000 21330 6020 21370
rect 6090 21330 6110 21400
rect 6180 21330 6200 21370
rect 6270 21330 6290 21370
rect 6360 21330 6380 21370
rect 6450 21330 6470 21400
rect 6730 21370 6760 21610
rect 6540 21330 6560 21370
rect 6630 21330 6650 21370
rect 6720 21330 6760 21370
rect -5550 21320 6760 21330
rect 8140 21610 20450 21640
rect 8140 21370 8170 21610
rect 8410 21580 8500 21610
rect 8740 21580 8830 21610
rect 9070 21580 9160 21610
rect 9400 21580 9490 21610
rect 9730 21580 9820 21610
rect 10060 21580 10150 21610
rect 10390 21580 10480 21610
rect 10720 21580 10810 21610
rect 11050 21580 11180 21610
rect 11420 21580 11510 21610
rect 11750 21580 11840 21610
rect 12080 21580 12170 21610
rect 12410 21580 12500 21610
rect 12740 21580 12830 21610
rect 13070 21580 13160 21610
rect 13400 21580 13490 21610
rect 13730 21580 13820 21610
rect 14060 21580 14190 21610
rect 14430 21580 14520 21610
rect 14760 21580 14850 21610
rect 15090 21580 15180 21610
rect 15420 21580 15510 21610
rect 15750 21580 15840 21610
rect 16080 21580 16170 21610
rect 16410 21580 16500 21610
rect 16740 21580 16830 21610
rect 17070 21580 17200 21610
rect 17440 21580 17530 21610
rect 17770 21580 17860 21610
rect 18100 21580 18190 21610
rect 18430 21580 18520 21610
rect 18760 21580 18850 21610
rect 19090 21580 19180 21610
rect 19420 21580 19510 21610
rect 19750 21580 19840 21610
rect 20080 21580 20450 21610
rect 8430 21510 8450 21580
rect 8790 21510 8810 21580
rect 9070 21510 9080 21580
rect 9150 21510 9160 21580
rect 9420 21510 9440 21580
rect 9780 21510 9800 21580
rect 10060 21510 10070 21580
rect 10140 21510 10150 21580
rect 10410 21510 10430 21580
rect 10770 21510 10790 21580
rect 11050 21510 11060 21580
rect 11130 21510 11180 21580
rect 11440 21510 11460 21580
rect 11800 21510 11820 21580
rect 12080 21510 12090 21580
rect 12160 21510 12170 21580
rect 12430 21510 12450 21580
rect 12790 21510 12810 21580
rect 13070 21510 13080 21580
rect 13150 21510 13160 21580
rect 13420 21510 13440 21580
rect 13780 21510 13800 21580
rect 14060 21510 14070 21580
rect 14140 21510 14190 21580
rect 14450 21510 14470 21580
rect 14810 21510 14830 21580
rect 15090 21510 15100 21580
rect 15170 21510 15180 21580
rect 15440 21510 15460 21580
rect 15800 21510 15820 21580
rect 16080 21510 16090 21580
rect 16160 21510 16170 21580
rect 16430 21510 16450 21580
rect 16790 21510 16810 21580
rect 17070 21510 17080 21580
rect 17150 21510 17200 21580
rect 17460 21510 17480 21580
rect 17820 21510 17840 21580
rect 18100 21510 18110 21580
rect 18180 21510 18190 21580
rect 18450 21510 18470 21580
rect 18810 21510 18830 21580
rect 19090 21510 19100 21580
rect 19170 21510 19180 21580
rect 19440 21510 19460 21580
rect 19800 21510 19820 21580
rect 20080 21510 20090 21580
rect 20160 21510 20450 21580
rect 8410 21490 8500 21510
rect 8740 21490 8830 21510
rect 9070 21490 9160 21510
rect 9400 21490 9490 21510
rect 9730 21490 9820 21510
rect 10060 21490 10150 21510
rect 10390 21490 10480 21510
rect 10720 21490 10810 21510
rect 11050 21490 11180 21510
rect 11420 21490 11510 21510
rect 11750 21490 11840 21510
rect 12080 21490 12170 21510
rect 12410 21490 12500 21510
rect 12740 21490 12830 21510
rect 13070 21490 13160 21510
rect 13400 21490 13490 21510
rect 13730 21490 13820 21510
rect 14060 21490 14190 21510
rect 14430 21490 14520 21510
rect 14760 21490 14850 21510
rect 15090 21490 15180 21510
rect 15420 21490 15510 21510
rect 15750 21490 15840 21510
rect 16080 21490 16170 21510
rect 16410 21490 16500 21510
rect 16740 21490 16830 21510
rect 17070 21490 17200 21510
rect 17440 21490 17530 21510
rect 17770 21490 17860 21510
rect 18100 21490 18190 21510
rect 18430 21490 18520 21510
rect 18760 21490 18850 21510
rect 19090 21490 19180 21510
rect 19420 21490 19510 21510
rect 19750 21490 19840 21510
rect 20080 21490 20450 21510
rect 8430 21420 8450 21490
rect 8790 21420 8810 21490
rect 9070 21420 9080 21490
rect 9150 21420 9160 21490
rect 9420 21420 9440 21490
rect 9780 21420 9800 21490
rect 10060 21420 10070 21490
rect 10140 21420 10150 21490
rect 10410 21420 10430 21490
rect 10770 21420 10790 21490
rect 11050 21420 11060 21490
rect 11130 21420 11180 21490
rect 11440 21420 11460 21490
rect 11800 21420 11820 21490
rect 12080 21420 12090 21490
rect 12160 21420 12170 21490
rect 12430 21420 12450 21490
rect 12790 21420 12810 21490
rect 13070 21420 13080 21490
rect 13150 21420 13160 21490
rect 13420 21420 13440 21490
rect 13780 21420 13800 21490
rect 14060 21420 14070 21490
rect 14140 21420 14190 21490
rect 14450 21420 14470 21490
rect 14810 21420 14830 21490
rect 15090 21420 15100 21490
rect 15170 21420 15180 21490
rect 15440 21420 15460 21490
rect 15800 21420 15820 21490
rect 16080 21420 16090 21490
rect 16160 21420 16170 21490
rect 16430 21420 16450 21490
rect 16790 21420 16810 21490
rect 17070 21420 17080 21490
rect 17150 21420 17200 21490
rect 17460 21420 17480 21490
rect 17820 21420 17840 21490
rect 18100 21420 18110 21490
rect 18180 21420 18190 21490
rect 18450 21420 18470 21490
rect 18810 21420 18830 21490
rect 19090 21420 19100 21490
rect 19170 21420 19180 21490
rect 19440 21420 19460 21490
rect 19800 21420 19820 21490
rect 20080 21420 20090 21490
rect 20160 21420 20450 21490
rect 8410 21400 8500 21420
rect 8740 21400 8830 21420
rect 9070 21400 9160 21420
rect 9400 21400 9490 21420
rect 9730 21400 9820 21420
rect 10060 21400 10150 21420
rect 10390 21400 10480 21420
rect 10720 21400 10810 21420
rect 11050 21400 11180 21420
rect 11420 21400 11510 21420
rect 11750 21400 11840 21420
rect 12080 21400 12170 21420
rect 12410 21400 12500 21420
rect 12740 21400 12830 21420
rect 13070 21400 13160 21420
rect 13400 21400 13490 21420
rect 13730 21400 13820 21420
rect 14060 21400 14190 21420
rect 14430 21400 14520 21420
rect 14760 21400 14850 21420
rect 15090 21400 15180 21420
rect 15420 21400 15510 21420
rect 15750 21400 15840 21420
rect 16080 21400 16170 21420
rect 16410 21400 16500 21420
rect 16740 21400 16830 21420
rect 17070 21400 17200 21420
rect 17440 21400 17530 21420
rect 17770 21400 17860 21420
rect 18100 21400 18190 21420
rect 18430 21400 18520 21420
rect 18760 21400 18850 21420
rect 19090 21400 19180 21420
rect 19420 21400 19510 21420
rect 19750 21400 19840 21420
rect 20080 21400 20450 21420
rect 8140 21330 8180 21370
rect 8250 21330 8270 21370
rect 8340 21330 8360 21370
rect 8430 21330 8450 21400
rect 8520 21330 8540 21370
rect 8610 21330 8630 21370
rect 8700 21330 8720 21370
rect 8790 21330 8810 21400
rect 9070 21370 9080 21400
rect 8880 21330 8900 21370
rect 8970 21330 8990 21370
rect 9060 21330 9080 21370
rect 9150 21370 9160 21400
rect 9150 21330 9170 21370
rect 9240 21330 9260 21370
rect 9330 21330 9350 21370
rect 9420 21330 9440 21400
rect 9510 21330 9530 21370
rect 9600 21330 9620 21370
rect 9690 21330 9710 21370
rect 9780 21330 9800 21400
rect 10060 21370 10070 21400
rect 9870 21330 9890 21370
rect 9960 21330 9980 21370
rect 10050 21330 10070 21370
rect 10140 21370 10150 21400
rect 10140 21330 10160 21370
rect 10230 21330 10250 21370
rect 10320 21330 10340 21370
rect 10410 21330 10430 21400
rect 10500 21330 10520 21370
rect 10590 21330 10610 21370
rect 10680 21330 10700 21370
rect 10770 21330 10790 21400
rect 11050 21370 11060 21400
rect 10860 21330 10880 21370
rect 10950 21330 10970 21370
rect 11040 21330 11060 21370
rect 11130 21370 11180 21400
rect 11130 21330 11190 21370
rect 11260 21330 11280 21370
rect 11350 21330 11370 21370
rect 11440 21330 11460 21400
rect 11530 21330 11550 21370
rect 11620 21330 11640 21370
rect 11710 21330 11730 21370
rect 11800 21330 11820 21400
rect 12080 21370 12090 21400
rect 11890 21330 11910 21370
rect 11980 21330 12000 21370
rect 12070 21330 12090 21370
rect 12160 21370 12170 21400
rect 12160 21330 12180 21370
rect 12250 21330 12270 21370
rect 12340 21330 12360 21370
rect 12430 21330 12450 21400
rect 12520 21330 12540 21370
rect 12610 21330 12630 21370
rect 12700 21330 12720 21370
rect 12790 21330 12810 21400
rect 13070 21370 13080 21400
rect 12880 21330 12900 21370
rect 12970 21330 12990 21370
rect 13060 21330 13080 21370
rect 13150 21370 13160 21400
rect 13150 21330 13170 21370
rect 13240 21330 13260 21370
rect 13330 21330 13350 21370
rect 13420 21330 13440 21400
rect 13510 21330 13530 21370
rect 13600 21330 13620 21370
rect 13690 21330 13710 21370
rect 13780 21330 13800 21400
rect 14060 21370 14070 21400
rect 13870 21330 13890 21370
rect 13960 21330 13980 21370
rect 14050 21330 14070 21370
rect 14140 21370 14190 21400
rect 14140 21330 14200 21370
rect 14270 21330 14290 21370
rect 14360 21330 14380 21370
rect 14450 21330 14470 21400
rect 14540 21330 14560 21370
rect 14630 21330 14650 21370
rect 14720 21330 14740 21370
rect 14810 21330 14830 21400
rect 15090 21370 15100 21400
rect 14900 21330 14920 21370
rect 14990 21330 15010 21370
rect 15080 21330 15100 21370
rect 15170 21370 15180 21400
rect 15170 21330 15190 21370
rect 15260 21330 15280 21370
rect 15350 21330 15370 21370
rect 15440 21330 15460 21400
rect 15530 21330 15550 21370
rect 15620 21330 15640 21370
rect 15710 21330 15730 21370
rect 15800 21330 15820 21400
rect 16080 21370 16090 21400
rect 15890 21330 15910 21370
rect 15980 21330 16000 21370
rect 16070 21330 16090 21370
rect 16160 21370 16170 21400
rect 16160 21330 16180 21370
rect 16250 21330 16270 21370
rect 16340 21330 16360 21370
rect 16430 21330 16450 21400
rect 16520 21330 16540 21370
rect 16610 21330 16630 21370
rect 16700 21330 16720 21370
rect 16790 21330 16810 21400
rect 17070 21370 17080 21400
rect 16880 21330 16900 21370
rect 16970 21330 16990 21370
rect 17060 21330 17080 21370
rect 17150 21370 17200 21400
rect 17150 21330 17210 21370
rect 17280 21330 17300 21370
rect 17370 21330 17390 21370
rect 17460 21330 17480 21400
rect 17550 21330 17570 21370
rect 17640 21330 17660 21370
rect 17730 21330 17750 21370
rect 17820 21330 17840 21400
rect 18100 21370 18110 21400
rect 17910 21330 17930 21370
rect 18000 21330 18020 21370
rect 18090 21330 18110 21370
rect 18180 21370 18190 21400
rect 18180 21330 18200 21370
rect 18270 21330 18290 21370
rect 18360 21330 18380 21370
rect 18450 21330 18470 21400
rect 18540 21330 18560 21370
rect 18630 21330 18650 21370
rect 18720 21330 18740 21370
rect 18810 21330 18830 21400
rect 19090 21370 19100 21400
rect 18900 21330 18920 21370
rect 18990 21330 19010 21370
rect 19080 21330 19100 21370
rect 19170 21370 19180 21400
rect 19170 21330 19190 21370
rect 19260 21330 19280 21370
rect 19350 21330 19370 21370
rect 19440 21330 19460 21400
rect 19530 21330 19550 21370
rect 19620 21330 19640 21370
rect 19710 21330 19730 21370
rect 19800 21330 19820 21400
rect 20080 21370 20090 21400
rect 19890 21330 19910 21370
rect 19980 21330 20000 21370
rect 20070 21330 20090 21370
rect 20160 21330 20450 21400
rect 8140 21320 20450 21330
rect -5550 20830 6760 21000
rect -5550 20590 -5200 20830
rect -4960 20590 -4870 20830
rect -4630 20590 -4540 20830
rect -4300 20590 -4210 20830
rect -3970 20590 -3880 20830
rect -3640 20590 -3550 20830
rect -3310 20590 -3220 20830
rect -2980 20590 -2890 20830
rect -2650 20590 -2560 20830
rect -2320 20590 -2230 20830
rect -1990 20590 -1900 20830
rect -1660 20590 -1570 20830
rect -1330 20590 -1240 20830
rect -1000 20590 -910 20830
rect -670 20590 -580 20830
rect -340 20590 -250 20830
rect -10 20590 80 20830
rect 320 20590 410 20830
rect 650 20590 740 20830
rect 980 20590 1070 20830
rect 1310 20590 1400 20830
rect 1640 20590 1730 20830
rect 1970 20590 2060 20830
rect 2300 20590 2390 20830
rect 2630 20590 2720 20830
rect 2960 20590 3050 20830
rect 3290 20590 3380 20830
rect 3620 20590 3710 20830
rect 3950 20590 4040 20830
rect 4280 20590 4370 20830
rect 4610 20590 4700 20830
rect 4940 20590 5030 20830
rect 5270 20590 5360 20830
rect 5600 20590 5690 20830
rect 5930 20590 6020 20830
rect 6260 20590 6350 20830
rect 6590 20590 6760 20830
rect -5550 20500 6760 20590
rect -5550 20260 -5200 20500
rect -4960 20260 -4870 20500
rect -4630 20260 -4540 20500
rect -4300 20260 -4210 20500
rect -3970 20260 -3880 20500
rect -3640 20260 -3550 20500
rect -3310 20260 -3220 20500
rect -2980 20260 -2890 20500
rect -2650 20260 -2560 20500
rect -2320 20260 -2230 20500
rect -1990 20260 -1900 20500
rect -1660 20260 -1570 20500
rect -1330 20260 -1240 20500
rect -1000 20260 -910 20500
rect -670 20260 -580 20500
rect -340 20260 -250 20500
rect -10 20260 80 20500
rect 320 20260 410 20500
rect 650 20260 740 20500
rect 980 20260 1070 20500
rect 1310 20260 1400 20500
rect 1640 20260 1730 20500
rect 1970 20260 2060 20500
rect 2300 20260 2390 20500
rect 2630 20260 2720 20500
rect 2960 20260 3050 20500
rect 3290 20260 3380 20500
rect 3620 20260 3710 20500
rect 3950 20260 4040 20500
rect 4280 20260 4370 20500
rect 4610 20260 4700 20500
rect 4940 20260 5030 20500
rect 5270 20260 5360 20500
rect 5600 20260 5690 20500
rect 5930 20260 6020 20500
rect 6260 20260 6350 20500
rect 6590 20260 6760 20500
rect -5550 20170 6760 20260
rect -5550 19930 -5200 20170
rect -4960 19930 -4870 20170
rect -4630 19930 -4540 20170
rect -4300 19930 -4210 20170
rect -3970 19930 -3880 20170
rect -3640 19930 -3550 20170
rect -3310 19930 -3220 20170
rect -2980 19930 -2890 20170
rect -2650 19930 -2560 20170
rect -2320 19930 -2230 20170
rect -1990 19930 -1900 20170
rect -1660 19930 -1570 20170
rect -1330 19930 -1240 20170
rect -1000 19930 -910 20170
rect -670 19930 -580 20170
rect -340 19930 -250 20170
rect -10 19930 80 20170
rect 320 19930 410 20170
rect 650 19930 740 20170
rect 980 19930 1070 20170
rect 1310 19930 1400 20170
rect 1640 19930 1730 20170
rect 1970 19930 2060 20170
rect 2300 19930 2390 20170
rect 2630 19930 2720 20170
rect 2960 19930 3050 20170
rect 3290 19930 3380 20170
rect 3620 19930 3710 20170
rect 3950 19930 4040 20170
rect 4280 19930 4370 20170
rect 4610 19930 4700 20170
rect 4940 19930 5030 20170
rect 5270 19930 5360 20170
rect 5600 19930 5690 20170
rect 5930 19930 6020 20170
rect 6260 19930 6350 20170
rect 6590 19930 6760 20170
rect -5550 19840 6760 19930
rect -5550 19600 -5200 19840
rect -4960 19600 -4870 19840
rect -4630 19600 -4540 19840
rect -4300 19600 -4210 19840
rect -3970 19600 -3880 19840
rect -3640 19600 -3550 19840
rect -3310 19600 -3220 19840
rect -2980 19600 -2890 19840
rect -2650 19600 -2560 19840
rect -2320 19600 -2230 19840
rect -1990 19600 -1900 19840
rect -1660 19600 -1570 19840
rect -1330 19600 -1240 19840
rect -1000 19600 -910 19840
rect -670 19600 -580 19840
rect -340 19600 -250 19840
rect -10 19600 80 19840
rect 320 19600 410 19840
rect 650 19600 740 19840
rect 980 19600 1070 19840
rect 1310 19600 1400 19840
rect 1640 19600 1730 19840
rect 1970 19600 2060 19840
rect 2300 19600 2390 19840
rect 2630 19600 2720 19840
rect 2960 19600 3050 19840
rect 3290 19600 3380 19840
rect 3620 19600 3710 19840
rect 3950 19600 4040 19840
rect 4280 19600 4370 19840
rect 4610 19600 4700 19840
rect 4940 19600 5030 19840
rect 5270 19600 5360 19840
rect 5600 19600 5690 19840
rect 5930 19600 6020 19840
rect 6260 19600 6350 19840
rect 6590 19600 6760 19840
rect -5550 19510 6760 19600
rect -5550 19270 -5200 19510
rect -4960 19270 -4870 19510
rect -4630 19270 -4540 19510
rect -4300 19270 -4210 19510
rect -3970 19270 -3880 19510
rect -3640 19270 -3550 19510
rect -3310 19270 -3220 19510
rect -2980 19270 -2890 19510
rect -2650 19270 -2560 19510
rect -2320 19270 -2230 19510
rect -1990 19270 -1900 19510
rect -1660 19270 -1570 19510
rect -1330 19270 -1240 19510
rect -1000 19270 -910 19510
rect -670 19270 -580 19510
rect -340 19270 -250 19510
rect -10 19270 80 19510
rect 320 19270 410 19510
rect 650 19270 740 19510
rect 980 19270 1070 19510
rect 1310 19270 1400 19510
rect 1640 19270 1730 19510
rect 1970 19270 2060 19510
rect 2300 19270 2390 19510
rect 2630 19270 2720 19510
rect 2960 19270 3050 19510
rect 3290 19270 3380 19510
rect 3620 19270 3710 19510
rect 3950 19270 4040 19510
rect 4280 19270 4370 19510
rect 4610 19270 4700 19510
rect 4940 19270 5030 19510
rect 5270 19270 5360 19510
rect 5600 19270 5690 19510
rect 5930 19270 6020 19510
rect 6260 19270 6350 19510
rect 6590 19270 6760 19510
rect -5550 19180 6760 19270
rect -5550 18940 -5200 19180
rect -4960 18940 -4870 19180
rect -4630 18940 -4540 19180
rect -4300 18940 -4210 19180
rect -3970 18940 -3880 19180
rect -3640 18940 -3550 19180
rect -3310 18940 -3220 19180
rect -2980 18940 -2890 19180
rect -2650 18940 -2560 19180
rect -2320 18940 -2230 19180
rect -1990 18940 -1900 19180
rect -1660 18940 -1570 19180
rect -1330 18940 -1240 19180
rect -1000 18940 -910 19180
rect -670 18940 -580 19180
rect -340 18940 -250 19180
rect -10 18940 80 19180
rect 320 18940 410 19180
rect 650 18940 740 19180
rect 980 18940 1070 19180
rect 1310 18940 1400 19180
rect 1640 18940 1730 19180
rect 1970 18940 2060 19180
rect 2300 18940 2390 19180
rect 2630 18940 2720 19180
rect 2960 18940 3050 19180
rect 3290 18940 3380 19180
rect 3620 18940 3710 19180
rect 3950 18940 4040 19180
rect 4280 18940 4370 19180
rect 4610 18940 4700 19180
rect 4940 18940 5030 19180
rect 5270 18940 5360 19180
rect 5600 18940 5690 19180
rect 5930 18940 6020 19180
rect 6260 18940 6350 19180
rect 6590 18940 6760 19180
rect -5550 18850 6760 18940
rect -5550 18610 -5200 18850
rect -4960 18610 -4870 18850
rect -4630 18610 -4540 18850
rect -4300 18610 -4210 18850
rect -3970 18610 -3880 18850
rect -3640 18610 -3550 18850
rect -3310 18610 -3220 18850
rect -2980 18610 -2890 18850
rect -2650 18610 -2560 18850
rect -2320 18610 -2230 18850
rect -1990 18610 -1900 18850
rect -1660 18610 -1570 18850
rect -1330 18610 -1240 18850
rect -1000 18610 -910 18850
rect -670 18610 -580 18850
rect -340 18610 -250 18850
rect -10 18610 80 18850
rect 320 18610 410 18850
rect 650 18610 740 18850
rect 980 18610 1070 18850
rect 1310 18610 1400 18850
rect 1640 18610 1730 18850
rect 1970 18610 2060 18850
rect 2300 18610 2390 18850
rect 2630 18610 2720 18850
rect 2960 18610 3050 18850
rect 3290 18610 3380 18850
rect 3620 18610 3710 18850
rect 3950 18610 4040 18850
rect 4280 18610 4370 18850
rect 4610 18610 4700 18850
rect 4940 18610 5030 18850
rect 5270 18610 5360 18850
rect 5600 18610 5690 18850
rect 5930 18610 6020 18850
rect 6260 18610 6350 18850
rect 6590 18610 6760 18850
rect -5550 18520 6760 18610
rect -5550 18280 -5200 18520
rect -4960 18280 -4870 18520
rect -4630 18280 -4540 18520
rect -4300 18280 -4210 18520
rect -3970 18280 -3880 18520
rect -3640 18280 -3550 18520
rect -3310 18280 -3220 18520
rect -2980 18280 -2890 18520
rect -2650 18280 -2560 18520
rect -2320 18280 -2230 18520
rect -1990 18280 -1900 18520
rect -1660 18280 -1570 18520
rect -1330 18280 -1240 18520
rect -1000 18280 -910 18520
rect -670 18280 -580 18520
rect -340 18280 -250 18520
rect -10 18280 80 18520
rect 320 18280 410 18520
rect 650 18280 740 18520
rect 980 18280 1070 18520
rect 1310 18280 1400 18520
rect 1640 18280 1730 18520
rect 1970 18280 2060 18520
rect 2300 18280 2390 18520
rect 2630 18280 2720 18520
rect 2960 18280 3050 18520
rect 3290 18280 3380 18520
rect 3620 18280 3710 18520
rect 3950 18280 4040 18520
rect 4280 18280 4370 18520
rect 4610 18280 4700 18520
rect 4940 18280 5030 18520
rect 5270 18280 5360 18520
rect 5600 18280 5690 18520
rect 5930 18280 6020 18520
rect 6260 18280 6350 18520
rect 6590 18280 6760 18520
rect -5550 18190 6760 18280
rect -5550 17950 -5200 18190
rect -4960 17950 -4870 18190
rect -4630 17950 -4540 18190
rect -4300 17950 -4210 18190
rect -3970 17950 -3880 18190
rect -3640 17950 -3550 18190
rect -3310 17950 -3220 18190
rect -2980 17950 -2890 18190
rect -2650 17950 -2560 18190
rect -2320 17950 -2230 18190
rect -1990 17950 -1900 18190
rect -1660 17950 -1570 18190
rect -1330 17950 -1240 18190
rect -1000 17950 -910 18190
rect -670 17950 -580 18190
rect -340 17950 -250 18190
rect -10 17950 80 18190
rect 320 17950 410 18190
rect 650 17950 740 18190
rect 980 17950 1070 18190
rect 1310 17950 1400 18190
rect 1640 17950 1730 18190
rect 1970 17950 2060 18190
rect 2300 17950 2390 18190
rect 2630 17950 2720 18190
rect 2960 17950 3050 18190
rect 3290 17950 3380 18190
rect 3620 17950 3710 18190
rect 3950 17950 4040 18190
rect 4280 17950 4370 18190
rect 4610 17950 4700 18190
rect 4940 17950 5030 18190
rect 5270 17950 5360 18190
rect 5600 17950 5690 18190
rect 5930 17950 6020 18190
rect 6260 17950 6350 18190
rect 6590 17950 6760 18190
rect -5550 17860 6760 17950
rect -5550 17620 -5200 17860
rect -4960 17620 -4870 17860
rect -4630 17620 -4540 17860
rect -4300 17620 -4210 17860
rect -3970 17620 -3880 17860
rect -3640 17620 -3550 17860
rect -3310 17620 -3220 17860
rect -2980 17620 -2890 17860
rect -2650 17620 -2560 17860
rect -2320 17620 -2230 17860
rect -1990 17620 -1900 17860
rect -1660 17620 -1570 17860
rect -1330 17620 -1240 17860
rect -1000 17620 -910 17860
rect -670 17620 -580 17860
rect -340 17620 -250 17860
rect -10 17620 80 17860
rect 320 17620 410 17860
rect 650 17620 740 17860
rect 980 17620 1070 17860
rect 1310 17620 1400 17860
rect 1640 17620 1730 17860
rect 1970 17620 2060 17860
rect 2300 17620 2390 17860
rect 2630 17620 2720 17860
rect 2960 17620 3050 17860
rect 3290 17620 3380 17860
rect 3620 17620 3710 17860
rect 3950 17620 4040 17860
rect 4280 17620 4370 17860
rect 4610 17620 4700 17860
rect 4940 17620 5030 17860
rect 5270 17620 5360 17860
rect 5600 17620 5690 17860
rect 5930 17620 6020 17860
rect 6260 17620 6350 17860
rect 6590 17620 6760 17860
rect -5550 17530 6760 17620
rect -5550 17290 -5200 17530
rect -4960 17290 -4870 17530
rect -4630 17290 -4540 17530
rect -4300 17290 -4210 17530
rect -3970 17290 -3880 17530
rect -3640 17290 -3550 17530
rect -3310 17290 -3220 17530
rect -2980 17290 -2890 17530
rect -2650 17290 -2560 17530
rect -2320 17290 -2230 17530
rect -1990 17290 -1900 17530
rect -1660 17290 -1570 17530
rect -1330 17290 -1240 17530
rect -1000 17290 -910 17530
rect -670 17290 -580 17530
rect -340 17290 -250 17530
rect -10 17290 80 17530
rect 320 17290 410 17530
rect 650 17290 740 17530
rect 980 17290 1070 17530
rect 1310 17290 1400 17530
rect 1640 17290 1730 17530
rect 1970 17290 2060 17530
rect 2300 17290 2390 17530
rect 2630 17290 2720 17530
rect 2960 17290 3050 17530
rect 3290 17290 3380 17530
rect 3620 17290 3710 17530
rect 3950 17290 4040 17530
rect 4280 17290 4370 17530
rect 4610 17290 4700 17530
rect 4940 17290 5030 17530
rect 5270 17290 5360 17530
rect 5600 17290 5690 17530
rect 5930 17290 6020 17530
rect 6260 17290 6350 17530
rect 6590 17290 6760 17530
rect -5550 17200 6760 17290
rect -5550 16960 -5200 17200
rect -4960 16960 -4870 17200
rect -4630 16960 -4540 17200
rect -4300 16960 -4210 17200
rect -3970 16960 -3880 17200
rect -3640 16960 -3550 17200
rect -3310 16960 -3220 17200
rect -2980 16960 -2890 17200
rect -2650 16960 -2560 17200
rect -2320 16960 -2230 17200
rect -1990 16960 -1900 17200
rect -1660 16960 -1570 17200
rect -1330 16960 -1240 17200
rect -1000 16960 -910 17200
rect -670 16960 -580 17200
rect -340 16960 -250 17200
rect -10 16960 80 17200
rect 320 16960 410 17200
rect 650 16960 740 17200
rect 980 16960 1070 17200
rect 1310 16960 1400 17200
rect 1640 16960 1730 17200
rect 1970 16960 2060 17200
rect 2300 16960 2390 17200
rect 2630 16960 2720 17200
rect 2960 16960 3050 17200
rect 3290 16960 3380 17200
rect 3620 16960 3710 17200
rect 3950 16960 4040 17200
rect 4280 16960 4370 17200
rect 4610 16960 4700 17200
rect 4940 16960 5030 17200
rect 5270 16960 5360 17200
rect 5600 16960 5690 17200
rect 5930 16960 6020 17200
rect 6260 16960 6350 17200
rect 6590 16960 6760 17200
rect -5550 16870 6760 16960
rect -5550 16630 -5200 16870
rect -4960 16630 -4870 16870
rect -4630 16630 -4540 16870
rect -4300 16630 -4210 16870
rect -3970 16630 -3880 16870
rect -3640 16630 -3550 16870
rect -3310 16630 -3220 16870
rect -2980 16630 -2890 16870
rect -2650 16630 -2560 16870
rect -2320 16630 -2230 16870
rect -1990 16630 -1900 16870
rect -1660 16630 -1570 16870
rect -1330 16630 -1240 16870
rect -1000 16630 -910 16870
rect -670 16630 -580 16870
rect -340 16630 -250 16870
rect -10 16630 80 16870
rect 320 16630 410 16870
rect 650 16630 740 16870
rect 980 16630 1070 16870
rect 1310 16630 1400 16870
rect 1640 16630 1730 16870
rect 1970 16630 2060 16870
rect 2300 16630 2390 16870
rect 2630 16630 2720 16870
rect 2960 16630 3050 16870
rect 3290 16630 3380 16870
rect 3620 16630 3710 16870
rect 3950 16630 4040 16870
rect 4280 16630 4370 16870
rect 4610 16630 4700 16870
rect 4940 16630 5030 16870
rect 5270 16630 5360 16870
rect 5600 16630 5690 16870
rect 5930 16630 6020 16870
rect 6260 16630 6350 16870
rect 6590 16630 6760 16870
rect -5550 16540 6760 16630
rect -5550 16300 -5200 16540
rect -4960 16300 -4870 16540
rect -4630 16300 -4540 16540
rect -4300 16300 -4210 16540
rect -3970 16300 -3880 16540
rect -3640 16300 -3550 16540
rect -3310 16300 -3220 16540
rect -2980 16300 -2890 16540
rect -2650 16300 -2560 16540
rect -2320 16300 -2230 16540
rect -1990 16300 -1900 16540
rect -1660 16300 -1570 16540
rect -1330 16300 -1240 16540
rect -1000 16300 -910 16540
rect -670 16300 -580 16540
rect -340 16300 -250 16540
rect -10 16300 80 16540
rect 320 16300 410 16540
rect 650 16300 740 16540
rect 980 16300 1070 16540
rect 1310 16300 1400 16540
rect 1640 16300 1730 16540
rect 1970 16300 2060 16540
rect 2300 16300 2390 16540
rect 2630 16300 2720 16540
rect 2960 16300 3050 16540
rect 3290 16300 3380 16540
rect 3620 16300 3710 16540
rect 3950 16300 4040 16540
rect 4280 16300 4370 16540
rect 4610 16300 4700 16540
rect 4940 16300 5030 16540
rect 5270 16300 5360 16540
rect 5600 16300 5690 16540
rect 5930 16300 6020 16540
rect 6260 16300 6350 16540
rect 6590 16300 6760 16540
rect -5550 16210 6760 16300
rect -5550 15970 -5200 16210
rect -4960 15970 -4870 16210
rect -4630 15970 -4540 16210
rect -4300 15970 -4210 16210
rect -3970 15970 -3880 16210
rect -3640 15970 -3550 16210
rect -3310 15970 -3220 16210
rect -2980 15970 -2890 16210
rect -2650 15970 -2560 16210
rect -2320 15970 -2230 16210
rect -1990 15970 -1900 16210
rect -1660 15970 -1570 16210
rect -1330 15970 -1240 16210
rect -1000 15970 -910 16210
rect -670 15970 -580 16210
rect -340 15970 -250 16210
rect -10 15970 80 16210
rect 320 15970 410 16210
rect 650 15970 740 16210
rect 980 15970 1070 16210
rect 1310 15970 1400 16210
rect 1640 15970 1730 16210
rect 1970 15970 2060 16210
rect 2300 15970 2390 16210
rect 2630 15970 2720 16210
rect 2960 15970 3050 16210
rect 3290 15970 3380 16210
rect 3620 15970 3710 16210
rect 3950 15970 4040 16210
rect 4280 15970 4370 16210
rect 4610 15970 4700 16210
rect 4940 15970 5030 16210
rect 5270 15970 5360 16210
rect 5600 15970 5690 16210
rect 5930 15970 6020 16210
rect 6260 15970 6350 16210
rect 6590 15970 6760 16210
rect -5550 15880 6760 15970
rect -5550 15640 -5200 15880
rect -4960 15640 -4870 15880
rect -4630 15640 -4540 15880
rect -4300 15640 -4210 15880
rect -3970 15640 -3880 15880
rect -3640 15640 -3550 15880
rect -3310 15640 -3220 15880
rect -2980 15640 -2890 15880
rect -2650 15640 -2560 15880
rect -2320 15640 -2230 15880
rect -1990 15640 -1900 15880
rect -1660 15640 -1570 15880
rect -1330 15640 -1240 15880
rect -1000 15640 -910 15880
rect -670 15640 -580 15880
rect -340 15640 -250 15880
rect -10 15640 80 15880
rect 320 15640 410 15880
rect 650 15640 740 15880
rect 980 15640 1070 15880
rect 1310 15640 1400 15880
rect 1640 15640 1730 15880
rect 1970 15640 2060 15880
rect 2300 15640 2390 15880
rect 2630 15640 2720 15880
rect 2960 15640 3050 15880
rect 3290 15640 3380 15880
rect 3620 15640 3710 15880
rect 3950 15640 4040 15880
rect 4280 15640 4370 15880
rect 4610 15640 4700 15880
rect 4940 15640 5030 15880
rect 5270 15640 5360 15880
rect 5600 15640 5690 15880
rect 5930 15640 6020 15880
rect 6260 15640 6350 15880
rect 6590 15640 6760 15880
rect -5550 15550 6760 15640
rect -5550 15310 -5200 15550
rect -4960 15310 -4870 15550
rect -4630 15310 -4540 15550
rect -4300 15310 -4210 15550
rect -3970 15310 -3880 15550
rect -3640 15310 -3550 15550
rect -3310 15310 -3220 15550
rect -2980 15310 -2890 15550
rect -2650 15310 -2560 15550
rect -2320 15310 -2230 15550
rect -1990 15310 -1900 15550
rect -1660 15310 -1570 15550
rect -1330 15310 -1240 15550
rect -1000 15310 -910 15550
rect -670 15310 -580 15550
rect -340 15310 -250 15550
rect -10 15310 80 15550
rect 320 15310 410 15550
rect 650 15310 740 15550
rect 980 15310 1070 15550
rect 1310 15310 1400 15550
rect 1640 15310 1730 15550
rect 1970 15310 2060 15550
rect 2300 15310 2390 15550
rect 2630 15310 2720 15550
rect 2960 15310 3050 15550
rect 3290 15310 3380 15550
rect 3620 15310 3710 15550
rect 3950 15310 4040 15550
rect 4280 15310 4370 15550
rect 4610 15310 4700 15550
rect 4940 15310 5030 15550
rect 5270 15310 5360 15550
rect 5600 15310 5690 15550
rect 5930 15310 6020 15550
rect 6260 15310 6350 15550
rect 6590 15310 6760 15550
rect -5550 15220 6760 15310
rect -5550 14980 -5200 15220
rect -4960 14980 -4870 15220
rect -4630 14980 -4540 15220
rect -4300 14980 -4210 15220
rect -3970 14980 -3880 15220
rect -3640 14980 -3550 15220
rect -3310 14980 -3220 15220
rect -2980 14980 -2890 15220
rect -2650 14980 -2560 15220
rect -2320 14980 -2230 15220
rect -1990 14980 -1900 15220
rect -1660 14980 -1570 15220
rect -1330 14980 -1240 15220
rect -1000 14980 -910 15220
rect -670 14980 -580 15220
rect -340 14980 -250 15220
rect -10 14980 80 15220
rect 320 14980 410 15220
rect 650 14980 740 15220
rect 980 14980 1070 15220
rect 1310 14980 1400 15220
rect 1640 14980 1730 15220
rect 1970 14980 2060 15220
rect 2300 14980 2390 15220
rect 2630 14980 2720 15220
rect 2960 14980 3050 15220
rect 3290 14980 3380 15220
rect 3620 14980 3710 15220
rect 3950 14980 4040 15220
rect 4280 14980 4370 15220
rect 4610 14980 4700 15220
rect 4940 14980 5030 15220
rect 5270 14980 5360 15220
rect 5600 14980 5690 15220
rect 5930 14980 6020 15220
rect 6260 14980 6350 15220
rect 6590 14980 6760 15220
rect -5550 14890 6760 14980
rect -5550 14650 -5200 14890
rect -4960 14650 -4870 14890
rect -4630 14650 -4540 14890
rect -4300 14650 -4210 14890
rect -3970 14650 -3880 14890
rect -3640 14650 -3550 14890
rect -3310 14650 -3220 14890
rect -2980 14650 -2890 14890
rect -2650 14650 -2560 14890
rect -2320 14650 -2230 14890
rect -1990 14650 -1900 14890
rect -1660 14650 -1570 14890
rect -1330 14650 -1240 14890
rect -1000 14650 -910 14890
rect -670 14650 -580 14890
rect -340 14650 -250 14890
rect -10 14650 80 14890
rect 320 14650 410 14890
rect 650 14650 740 14890
rect 980 14650 1070 14890
rect 1310 14650 1400 14890
rect 1640 14650 1730 14890
rect 1970 14650 2060 14890
rect 2300 14650 2390 14890
rect 2630 14650 2720 14890
rect 2960 14650 3050 14890
rect 3290 14650 3380 14890
rect 3620 14650 3710 14890
rect 3950 14650 4040 14890
rect 4280 14650 4370 14890
rect 4610 14650 4700 14890
rect 4940 14650 5030 14890
rect 5270 14650 5360 14890
rect 5600 14650 5690 14890
rect 5930 14650 6020 14890
rect 6260 14650 6350 14890
rect 6590 14650 6760 14890
rect -5550 14560 6760 14650
rect -5550 14320 -5200 14560
rect -4960 14320 -4870 14560
rect -4630 14320 -4540 14560
rect -4300 14320 -4210 14560
rect -3970 14320 -3880 14560
rect -3640 14320 -3550 14560
rect -3310 14320 -3220 14560
rect -2980 14320 -2890 14560
rect -2650 14320 -2560 14560
rect -2320 14320 -2230 14560
rect -1990 14320 -1900 14560
rect -1660 14320 -1570 14560
rect -1330 14320 -1240 14560
rect -1000 14320 -910 14560
rect -670 14320 -580 14560
rect -340 14320 -250 14560
rect -10 14320 80 14560
rect 320 14320 410 14560
rect 650 14320 740 14560
rect 980 14320 1070 14560
rect 1310 14320 1400 14560
rect 1640 14320 1730 14560
rect 1970 14320 2060 14560
rect 2300 14320 2390 14560
rect 2630 14320 2720 14560
rect 2960 14320 3050 14560
rect 3290 14320 3380 14560
rect 3620 14320 3710 14560
rect 3950 14320 4040 14560
rect 4280 14320 4370 14560
rect 4610 14320 4700 14560
rect 4940 14320 5030 14560
rect 5270 14320 5360 14560
rect 5600 14320 5690 14560
rect 5930 14320 6020 14560
rect 6260 14320 6350 14560
rect 6590 14320 6760 14560
rect -5550 14230 6760 14320
rect -5550 13990 -5200 14230
rect -4960 13990 -4870 14230
rect -4630 13990 -4540 14230
rect -4300 13990 -4210 14230
rect -3970 13990 -3880 14230
rect -3640 13990 -3550 14230
rect -3310 13990 -3220 14230
rect -2980 13990 -2890 14230
rect -2650 13990 -2560 14230
rect -2320 13990 -2230 14230
rect -1990 13990 -1900 14230
rect -1660 13990 -1570 14230
rect -1330 13990 -1240 14230
rect -1000 13990 -910 14230
rect -670 13990 -580 14230
rect -340 13990 -250 14230
rect -10 13990 80 14230
rect 320 13990 410 14230
rect 650 13990 740 14230
rect 980 13990 1070 14230
rect 1310 13990 1400 14230
rect 1640 13990 1730 14230
rect 1970 13990 2060 14230
rect 2300 13990 2390 14230
rect 2630 13990 2720 14230
rect 2960 13990 3050 14230
rect 3290 13990 3380 14230
rect 3620 13990 3710 14230
rect 3950 13990 4040 14230
rect 4280 13990 4370 14230
rect 4610 13990 4700 14230
rect 4940 13990 5030 14230
rect 5270 13990 5360 14230
rect 5600 13990 5690 14230
rect 5930 13990 6020 14230
rect 6260 13990 6350 14230
rect 6590 13990 6760 14230
rect -5550 13900 6760 13990
rect -5550 13660 -5200 13900
rect -4960 13660 -4870 13900
rect -4630 13660 -4540 13900
rect -4300 13660 -4210 13900
rect -3970 13660 -3880 13900
rect -3640 13660 -3550 13900
rect -3310 13660 -3220 13900
rect -2980 13660 -2890 13900
rect -2650 13660 -2560 13900
rect -2320 13660 -2230 13900
rect -1990 13660 -1900 13900
rect -1660 13660 -1570 13900
rect -1330 13660 -1240 13900
rect -1000 13660 -910 13900
rect -670 13660 -580 13900
rect -340 13660 -250 13900
rect -10 13660 80 13900
rect 320 13660 410 13900
rect 650 13660 740 13900
rect 980 13660 1070 13900
rect 1310 13660 1400 13900
rect 1640 13660 1730 13900
rect 1970 13660 2060 13900
rect 2300 13660 2390 13900
rect 2630 13660 2720 13900
rect 2960 13660 3050 13900
rect 3290 13660 3380 13900
rect 3620 13660 3710 13900
rect 3950 13660 4040 13900
rect 4280 13660 4370 13900
rect 4610 13660 4700 13900
rect 4940 13660 5030 13900
rect 5270 13660 5360 13900
rect 5600 13660 5690 13900
rect 5930 13660 6020 13900
rect 6260 13660 6350 13900
rect 6590 13660 6760 13900
rect -5550 13570 6760 13660
rect -5550 13330 -5200 13570
rect -4960 13330 -4870 13570
rect -4630 13330 -4540 13570
rect -4300 13330 -4210 13570
rect -3970 13330 -3880 13570
rect -3640 13330 -3550 13570
rect -3310 13330 -3220 13570
rect -2980 13330 -2890 13570
rect -2650 13330 -2560 13570
rect -2320 13330 -2230 13570
rect -1990 13330 -1900 13570
rect -1660 13330 -1570 13570
rect -1330 13330 -1240 13570
rect -1000 13330 -910 13570
rect -670 13330 -580 13570
rect -340 13330 -250 13570
rect -10 13330 80 13570
rect 320 13330 410 13570
rect 650 13330 740 13570
rect 980 13330 1070 13570
rect 1310 13330 1400 13570
rect 1640 13330 1730 13570
rect 1970 13330 2060 13570
rect 2300 13330 2390 13570
rect 2630 13330 2720 13570
rect 2960 13330 3050 13570
rect 3290 13330 3380 13570
rect 3620 13330 3710 13570
rect 3950 13330 4040 13570
rect 4280 13330 4370 13570
rect 4610 13330 4700 13570
rect 4940 13330 5030 13570
rect 5270 13330 5360 13570
rect 5600 13330 5690 13570
rect 5930 13330 6020 13570
rect 6260 13330 6350 13570
rect 6590 13330 6760 13570
rect -5550 13240 6760 13330
rect -5550 13000 -5200 13240
rect -4960 13000 -4870 13240
rect -4630 13000 -4540 13240
rect -4300 13000 -4210 13240
rect -3970 13000 -3880 13240
rect -3640 13000 -3550 13240
rect -3310 13000 -3220 13240
rect -2980 13000 -2890 13240
rect -2650 13000 -2560 13240
rect -2320 13000 -2230 13240
rect -1990 13000 -1900 13240
rect -1660 13000 -1570 13240
rect -1330 13000 -1240 13240
rect -1000 13000 -910 13240
rect -670 13000 -580 13240
rect -340 13000 -250 13240
rect -10 13000 80 13240
rect 320 13000 410 13240
rect 650 13000 740 13240
rect 980 13000 1070 13240
rect 1310 13000 1400 13240
rect 1640 13000 1730 13240
rect 1970 13000 2060 13240
rect 2300 13000 2390 13240
rect 2630 13000 2720 13240
rect 2960 13000 3050 13240
rect 3290 13000 3380 13240
rect 3620 13000 3710 13240
rect 3950 13000 4040 13240
rect 4280 13000 4370 13240
rect 4610 13000 4700 13240
rect 4940 13000 5030 13240
rect 5270 13000 5360 13240
rect 5600 13000 5690 13240
rect 5930 13000 6020 13240
rect 6260 13000 6350 13240
rect 6590 13000 6760 13240
rect -5550 12910 6760 13000
rect -5550 12670 -5200 12910
rect -4960 12670 -4870 12910
rect -4630 12670 -4540 12910
rect -4300 12670 -4210 12910
rect -3970 12670 -3880 12910
rect -3640 12670 -3550 12910
rect -3310 12670 -3220 12910
rect -2980 12670 -2890 12910
rect -2650 12670 -2560 12910
rect -2320 12670 -2230 12910
rect -1990 12670 -1900 12910
rect -1660 12670 -1570 12910
rect -1330 12670 -1240 12910
rect -1000 12670 -910 12910
rect -670 12670 -580 12910
rect -340 12670 -250 12910
rect -10 12670 80 12910
rect 320 12670 410 12910
rect 650 12670 740 12910
rect 980 12670 1070 12910
rect 1310 12670 1400 12910
rect 1640 12670 1730 12910
rect 1970 12670 2060 12910
rect 2300 12670 2390 12910
rect 2630 12670 2720 12910
rect 2960 12670 3050 12910
rect 3290 12670 3380 12910
rect 3620 12670 3710 12910
rect 3950 12670 4040 12910
rect 4280 12670 4370 12910
rect 4610 12670 4700 12910
rect 4940 12670 5030 12910
rect 5270 12670 5360 12910
rect 5600 12670 5690 12910
rect 5930 12670 6020 12910
rect 6260 12670 6350 12910
rect 6590 12670 6760 12910
rect -5550 12580 6760 12670
rect -5550 12340 -5200 12580
rect -4960 12340 -4870 12580
rect -4630 12340 -4540 12580
rect -4300 12340 -4210 12580
rect -3970 12340 -3880 12580
rect -3640 12340 -3550 12580
rect -3310 12340 -3220 12580
rect -2980 12340 -2890 12580
rect -2650 12340 -2560 12580
rect -2320 12340 -2230 12580
rect -1990 12340 -1900 12580
rect -1660 12340 -1570 12580
rect -1330 12340 -1240 12580
rect -1000 12340 -910 12580
rect -670 12340 -580 12580
rect -340 12340 -250 12580
rect -10 12340 80 12580
rect 320 12340 410 12580
rect 650 12340 740 12580
rect 980 12340 1070 12580
rect 1310 12340 1400 12580
rect 1640 12340 1730 12580
rect 1970 12340 2060 12580
rect 2300 12340 2390 12580
rect 2630 12340 2720 12580
rect 2960 12340 3050 12580
rect 3290 12340 3380 12580
rect 3620 12340 3710 12580
rect 3950 12340 4040 12580
rect 4280 12340 4370 12580
rect 4610 12340 4700 12580
rect 4940 12340 5030 12580
rect 5270 12340 5360 12580
rect 5600 12340 5690 12580
rect 5930 12340 6020 12580
rect 6260 12340 6350 12580
rect 6590 12340 6760 12580
rect -5550 12250 6760 12340
rect -5550 12010 -5200 12250
rect -4960 12010 -4870 12250
rect -4630 12010 -4540 12250
rect -4300 12010 -4210 12250
rect -3970 12010 -3880 12250
rect -3640 12010 -3550 12250
rect -3310 12010 -3220 12250
rect -2980 12010 -2890 12250
rect -2650 12010 -2560 12250
rect -2320 12010 -2230 12250
rect -1990 12010 -1900 12250
rect -1660 12010 -1570 12250
rect -1330 12010 -1240 12250
rect -1000 12010 -910 12250
rect -670 12010 -580 12250
rect -340 12010 -250 12250
rect -10 12010 80 12250
rect 320 12010 410 12250
rect 650 12010 740 12250
rect 980 12010 1070 12250
rect 1310 12010 1400 12250
rect 1640 12010 1730 12250
rect 1970 12010 2060 12250
rect 2300 12010 2390 12250
rect 2630 12010 2720 12250
rect 2960 12010 3050 12250
rect 3290 12010 3380 12250
rect 3620 12010 3710 12250
rect 3950 12010 4040 12250
rect 4280 12010 4370 12250
rect 4610 12010 4700 12250
rect 4940 12010 5030 12250
rect 5270 12010 5360 12250
rect 5600 12010 5690 12250
rect 5930 12010 6020 12250
rect 6260 12010 6350 12250
rect 6590 12010 6760 12250
rect -5550 11920 6760 12010
rect -5550 11680 -5200 11920
rect -4960 11680 -4870 11920
rect -4630 11680 -4540 11920
rect -4300 11680 -4210 11920
rect -3970 11680 -3880 11920
rect -3640 11680 -3550 11920
rect -3310 11680 -3220 11920
rect -2980 11680 -2890 11920
rect -2650 11680 -2560 11920
rect -2320 11680 -2230 11920
rect -1990 11680 -1900 11920
rect -1660 11680 -1570 11920
rect -1330 11680 -1240 11920
rect -1000 11680 -910 11920
rect -670 11680 -580 11920
rect -340 11680 -250 11920
rect -10 11680 80 11920
rect 320 11680 410 11920
rect 650 11680 740 11920
rect 980 11680 1070 11920
rect 1310 11680 1400 11920
rect 1640 11680 1730 11920
rect 1970 11680 2060 11920
rect 2300 11680 2390 11920
rect 2630 11680 2720 11920
rect 2960 11680 3050 11920
rect 3290 11680 3380 11920
rect 3620 11680 3710 11920
rect 3950 11680 4040 11920
rect 4280 11680 4370 11920
rect 4610 11680 4700 11920
rect 4940 11680 5030 11920
rect 5270 11680 5360 11920
rect 5600 11680 5690 11920
rect 5930 11680 6020 11920
rect 6260 11680 6350 11920
rect 6590 11680 6760 11920
rect -5550 11590 6760 11680
rect -5550 11350 -5200 11590
rect -4960 11350 -4870 11590
rect -4630 11350 -4540 11590
rect -4300 11350 -4210 11590
rect -3970 11350 -3880 11590
rect -3640 11350 -3550 11590
rect -3310 11350 -3220 11590
rect -2980 11350 -2890 11590
rect -2650 11350 -2560 11590
rect -2320 11350 -2230 11590
rect -1990 11350 -1900 11590
rect -1660 11350 -1570 11590
rect -1330 11350 -1240 11590
rect -1000 11350 -910 11590
rect -670 11350 -580 11590
rect -340 11350 -250 11590
rect -10 11350 80 11590
rect 320 11350 410 11590
rect 650 11350 740 11590
rect 980 11350 1070 11590
rect 1310 11350 1400 11590
rect 1640 11350 1730 11590
rect 1970 11350 2060 11590
rect 2300 11350 2390 11590
rect 2630 11350 2720 11590
rect 2960 11350 3050 11590
rect 3290 11350 3380 11590
rect 3620 11350 3710 11590
rect 3950 11350 4040 11590
rect 4280 11350 4370 11590
rect 4610 11350 4700 11590
rect 4940 11350 5030 11590
rect 5270 11350 5360 11590
rect 5600 11350 5690 11590
rect 5930 11350 6020 11590
rect 6260 11350 6350 11590
rect 6590 11350 6760 11590
rect -5550 11260 6760 11350
rect -5550 11020 -5200 11260
rect -4960 11020 -4870 11260
rect -4630 11020 -4540 11260
rect -4300 11020 -4210 11260
rect -3970 11020 -3880 11260
rect -3640 11020 -3550 11260
rect -3310 11020 -3220 11260
rect -2980 11020 -2890 11260
rect -2650 11020 -2560 11260
rect -2320 11020 -2230 11260
rect -1990 11020 -1900 11260
rect -1660 11020 -1570 11260
rect -1330 11020 -1240 11260
rect -1000 11020 -910 11260
rect -670 11020 -580 11260
rect -340 11020 -250 11260
rect -10 11020 80 11260
rect 320 11020 410 11260
rect 650 11020 740 11260
rect 980 11020 1070 11260
rect 1310 11020 1400 11260
rect 1640 11020 1730 11260
rect 1970 11020 2060 11260
rect 2300 11020 2390 11260
rect 2630 11020 2720 11260
rect 2960 11020 3050 11260
rect 3290 11020 3380 11260
rect 3620 11020 3710 11260
rect 3950 11020 4040 11260
rect 4280 11020 4370 11260
rect 4610 11020 4700 11260
rect 4940 11020 5030 11260
rect 5270 11020 5360 11260
rect 5600 11020 5690 11260
rect 5930 11020 6020 11260
rect 6260 11020 6350 11260
rect 6590 11020 6760 11260
rect -5550 10930 6760 11020
rect -5550 10690 -5200 10930
rect -4960 10690 -4870 10930
rect -4630 10690 -4540 10930
rect -4300 10690 -4210 10930
rect -3970 10690 -3880 10930
rect -3640 10690 -3550 10930
rect -3310 10690 -3220 10930
rect -2980 10690 -2890 10930
rect -2650 10690 -2560 10930
rect -2320 10690 -2230 10930
rect -1990 10690 -1900 10930
rect -1660 10690 -1570 10930
rect -1330 10690 -1240 10930
rect -1000 10690 -910 10930
rect -670 10690 -580 10930
rect -340 10690 -250 10930
rect -10 10690 80 10930
rect 320 10690 410 10930
rect 650 10690 740 10930
rect 980 10690 1070 10930
rect 1310 10690 1400 10930
rect 1640 10690 1730 10930
rect 1970 10690 2060 10930
rect 2300 10690 2390 10930
rect 2630 10690 2720 10930
rect 2960 10690 3050 10930
rect 3290 10690 3380 10930
rect 3620 10690 3710 10930
rect 3950 10690 4040 10930
rect 4280 10690 4370 10930
rect 4610 10690 4700 10930
rect 4940 10690 5030 10930
rect 5270 10690 5360 10930
rect 5600 10690 5690 10930
rect 5930 10690 6020 10930
rect 6260 10690 6350 10930
rect 6590 10690 6760 10930
rect -5550 10600 6760 10690
rect -5550 10360 -5200 10600
rect -4960 10360 -4870 10600
rect -4630 10360 -4540 10600
rect -4300 10360 -4210 10600
rect -3970 10360 -3880 10600
rect -3640 10360 -3550 10600
rect -3310 10360 -3220 10600
rect -2980 10360 -2890 10600
rect -2650 10360 -2560 10600
rect -2320 10360 -2230 10600
rect -1990 10360 -1900 10600
rect -1660 10360 -1570 10600
rect -1330 10360 -1240 10600
rect -1000 10360 -910 10600
rect -670 10360 -580 10600
rect -340 10360 -250 10600
rect -10 10360 80 10600
rect 320 10360 410 10600
rect 650 10360 740 10600
rect 980 10360 1070 10600
rect 1310 10360 1400 10600
rect 1640 10360 1730 10600
rect 1970 10360 2060 10600
rect 2300 10360 2390 10600
rect 2630 10360 2720 10600
rect 2960 10360 3050 10600
rect 3290 10360 3380 10600
rect 3620 10360 3710 10600
rect 3950 10360 4040 10600
rect 4280 10360 4370 10600
rect 4610 10360 4700 10600
rect 4940 10360 5030 10600
rect 5270 10360 5360 10600
rect 5600 10360 5690 10600
rect 5930 10360 6020 10600
rect 6260 10360 6350 10600
rect 6590 10360 6760 10600
rect -5550 10270 6760 10360
rect -5550 10030 -5200 10270
rect -4960 10030 -4870 10270
rect -4630 10030 -4540 10270
rect -4300 10030 -4210 10270
rect -3970 10030 -3880 10270
rect -3640 10030 -3550 10270
rect -3310 10030 -3220 10270
rect -2980 10030 -2890 10270
rect -2650 10030 -2560 10270
rect -2320 10030 -2230 10270
rect -1990 10030 -1900 10270
rect -1660 10030 -1570 10270
rect -1330 10030 -1240 10270
rect -1000 10030 -910 10270
rect -670 10030 -580 10270
rect -340 10030 -250 10270
rect -10 10030 80 10270
rect 320 10030 410 10270
rect 650 10030 740 10270
rect 980 10030 1070 10270
rect 1310 10030 1400 10270
rect 1640 10030 1730 10270
rect 1970 10030 2060 10270
rect 2300 10030 2390 10270
rect 2630 10030 2720 10270
rect 2960 10030 3050 10270
rect 3290 10030 3380 10270
rect 3620 10030 3710 10270
rect 3950 10030 4040 10270
rect 4280 10030 4370 10270
rect 4610 10030 4700 10270
rect 4940 10030 5030 10270
rect 5270 10030 5360 10270
rect 5600 10030 5690 10270
rect 5930 10030 6020 10270
rect 6260 10030 6350 10270
rect 6590 10030 6760 10270
rect -5550 9940 6760 10030
rect -5550 9700 -5200 9940
rect -4960 9700 -4870 9940
rect -4630 9700 -4540 9940
rect -4300 9700 -4210 9940
rect -3970 9700 -3880 9940
rect -3640 9700 -3550 9940
rect -3310 9700 -3220 9940
rect -2980 9700 -2890 9940
rect -2650 9700 -2560 9940
rect -2320 9700 -2230 9940
rect -1990 9700 -1900 9940
rect -1660 9700 -1570 9940
rect -1330 9700 -1240 9940
rect -1000 9700 -910 9940
rect -670 9700 -580 9940
rect -340 9700 -250 9940
rect -10 9700 80 9940
rect 320 9700 410 9940
rect 650 9700 740 9940
rect 980 9700 1070 9940
rect 1310 9700 1400 9940
rect 1640 9700 1730 9940
rect 1970 9700 2060 9940
rect 2300 9700 2390 9940
rect 2630 9700 2720 9940
rect 2960 9700 3050 9940
rect 3290 9700 3380 9940
rect 3620 9700 3710 9940
rect 3950 9700 4040 9940
rect 4280 9700 4370 9940
rect 4610 9700 4700 9940
rect 4940 9700 5030 9940
rect 5270 9700 5360 9940
rect 5600 9700 5690 9940
rect 5930 9700 6020 9940
rect 6260 9700 6350 9940
rect 6590 9700 6760 9940
rect -5550 9610 6760 9700
rect -5550 9370 -5200 9610
rect -4960 9370 -4870 9610
rect -4630 9370 -4540 9610
rect -4300 9370 -4210 9610
rect -3970 9370 -3880 9610
rect -3640 9370 -3550 9610
rect -3310 9370 -3220 9610
rect -2980 9370 -2890 9610
rect -2650 9370 -2560 9610
rect -2320 9370 -2230 9610
rect -1990 9370 -1900 9610
rect -1660 9370 -1570 9610
rect -1330 9370 -1240 9610
rect -1000 9370 -910 9610
rect -670 9370 -580 9610
rect -340 9370 -250 9610
rect -10 9370 80 9610
rect 320 9370 410 9610
rect 650 9370 740 9610
rect 980 9370 1070 9610
rect 1310 9370 1400 9610
rect 1640 9370 1730 9610
rect 1970 9370 2060 9610
rect 2300 9370 2390 9610
rect 2630 9370 2720 9610
rect 2960 9370 3050 9610
rect 3290 9370 3380 9610
rect 3620 9370 3710 9610
rect 3950 9370 4040 9610
rect 4280 9370 4370 9610
rect 4610 9370 4700 9610
rect 4940 9370 5030 9610
rect 5270 9370 5360 9610
rect 5600 9370 5690 9610
rect 5930 9370 6020 9610
rect 6260 9370 6350 9610
rect 6590 9370 6760 9610
rect -5550 9280 6760 9370
rect -5550 9040 -5200 9280
rect -4960 9040 -4870 9280
rect -4630 9040 -4540 9280
rect -4300 9040 -4210 9280
rect -3970 9040 -3880 9280
rect -3640 9040 -3550 9280
rect -3310 9040 -3220 9280
rect -2980 9040 -2890 9280
rect -2650 9040 -2560 9280
rect -2320 9040 -2230 9280
rect -1990 9040 -1900 9280
rect -1660 9040 -1570 9280
rect -1330 9040 -1240 9280
rect -1000 9040 -910 9280
rect -670 9040 -580 9280
rect -340 9040 -250 9280
rect -10 9040 80 9280
rect 320 9040 410 9280
rect 650 9040 740 9280
rect 980 9040 1070 9280
rect 1310 9040 1400 9280
rect 1640 9040 1730 9280
rect 1970 9040 2060 9280
rect 2300 9040 2390 9280
rect 2630 9040 2720 9280
rect 2960 9040 3050 9280
rect 3290 9040 3380 9280
rect 3620 9040 3710 9280
rect 3950 9040 4040 9280
rect 4280 9040 4370 9280
rect 4610 9040 4700 9280
rect 4940 9040 5030 9280
rect 5270 9040 5360 9280
rect 5600 9040 5690 9280
rect 5930 9040 6020 9280
rect 6260 9040 6350 9280
rect 6590 9040 6760 9280
rect -5550 8690 6760 9040
rect 6440 8410 6760 8690
rect 6440 8340 6470 8410
rect 6540 8340 6560 8410
rect 6630 8340 6650 8410
rect 6720 8340 6760 8410
rect 6440 8320 6760 8340
rect 6440 8250 6470 8320
rect 6540 8250 6560 8320
rect 6630 8250 6650 8320
rect 6720 8250 6760 8320
rect 6440 8230 6760 8250
rect 8140 20830 20450 21000
rect 8140 20590 8310 20830
rect 8550 20590 8640 20830
rect 8880 20590 8970 20830
rect 9210 20590 9300 20830
rect 9540 20590 9630 20830
rect 9870 20590 9960 20830
rect 10200 20590 10290 20830
rect 10530 20590 10620 20830
rect 10860 20590 10950 20830
rect 11190 20590 11280 20830
rect 11520 20590 11610 20830
rect 11850 20590 11940 20830
rect 12180 20590 12270 20830
rect 12510 20590 12600 20830
rect 12840 20590 12930 20830
rect 13170 20590 13260 20830
rect 13500 20590 13590 20830
rect 13830 20590 13920 20830
rect 14160 20590 14250 20830
rect 14490 20590 14580 20830
rect 14820 20590 14910 20830
rect 15150 20590 15240 20830
rect 15480 20590 15570 20830
rect 15810 20590 15900 20830
rect 16140 20590 16230 20830
rect 16470 20590 16560 20830
rect 16800 20590 16890 20830
rect 17130 20590 17220 20830
rect 17460 20590 17550 20830
rect 17790 20590 17880 20830
rect 18120 20590 18210 20830
rect 18450 20590 18540 20830
rect 18780 20590 18870 20830
rect 19110 20590 19200 20830
rect 19440 20590 19530 20830
rect 19770 20590 19860 20830
rect 20100 20590 20450 20830
rect 8140 20500 20450 20590
rect 8140 20260 8310 20500
rect 8550 20260 8640 20500
rect 8880 20260 8970 20500
rect 9210 20260 9300 20500
rect 9540 20260 9630 20500
rect 9870 20260 9960 20500
rect 10200 20260 10290 20500
rect 10530 20260 10620 20500
rect 10860 20260 10950 20500
rect 11190 20260 11280 20500
rect 11520 20260 11610 20500
rect 11850 20260 11940 20500
rect 12180 20260 12270 20500
rect 12510 20260 12600 20500
rect 12840 20260 12930 20500
rect 13170 20260 13260 20500
rect 13500 20260 13590 20500
rect 13830 20260 13920 20500
rect 14160 20260 14250 20500
rect 14490 20260 14580 20500
rect 14820 20260 14910 20500
rect 15150 20260 15240 20500
rect 15480 20260 15570 20500
rect 15810 20260 15900 20500
rect 16140 20260 16230 20500
rect 16470 20260 16560 20500
rect 16800 20260 16890 20500
rect 17130 20260 17220 20500
rect 17460 20260 17550 20500
rect 17790 20260 17880 20500
rect 18120 20260 18210 20500
rect 18450 20260 18540 20500
rect 18780 20260 18870 20500
rect 19110 20260 19200 20500
rect 19440 20260 19530 20500
rect 19770 20260 19860 20500
rect 20100 20260 20450 20500
rect 8140 20170 20450 20260
rect 8140 19930 8310 20170
rect 8550 19930 8640 20170
rect 8880 19930 8970 20170
rect 9210 19930 9300 20170
rect 9540 19930 9630 20170
rect 9870 19930 9960 20170
rect 10200 19930 10290 20170
rect 10530 19930 10620 20170
rect 10860 19930 10950 20170
rect 11190 19930 11280 20170
rect 11520 19930 11610 20170
rect 11850 19930 11940 20170
rect 12180 19930 12270 20170
rect 12510 19930 12600 20170
rect 12840 19930 12930 20170
rect 13170 19930 13260 20170
rect 13500 19930 13590 20170
rect 13830 19930 13920 20170
rect 14160 19930 14250 20170
rect 14490 19930 14580 20170
rect 14820 19930 14910 20170
rect 15150 19930 15240 20170
rect 15480 19930 15570 20170
rect 15810 19930 15900 20170
rect 16140 19930 16230 20170
rect 16470 19930 16560 20170
rect 16800 19930 16890 20170
rect 17130 19930 17220 20170
rect 17460 19930 17550 20170
rect 17790 19930 17880 20170
rect 18120 19930 18210 20170
rect 18450 19930 18540 20170
rect 18780 19930 18870 20170
rect 19110 19930 19200 20170
rect 19440 19930 19530 20170
rect 19770 19930 19860 20170
rect 20100 19930 20450 20170
rect 8140 19840 20450 19930
rect 8140 19600 8310 19840
rect 8550 19600 8640 19840
rect 8880 19600 8970 19840
rect 9210 19600 9300 19840
rect 9540 19600 9630 19840
rect 9870 19600 9960 19840
rect 10200 19600 10290 19840
rect 10530 19600 10620 19840
rect 10860 19600 10950 19840
rect 11190 19600 11280 19840
rect 11520 19600 11610 19840
rect 11850 19600 11940 19840
rect 12180 19600 12270 19840
rect 12510 19600 12600 19840
rect 12840 19600 12930 19840
rect 13170 19600 13260 19840
rect 13500 19600 13590 19840
rect 13830 19600 13920 19840
rect 14160 19600 14250 19840
rect 14490 19600 14580 19840
rect 14820 19600 14910 19840
rect 15150 19600 15240 19840
rect 15480 19600 15570 19840
rect 15810 19600 15900 19840
rect 16140 19600 16230 19840
rect 16470 19600 16560 19840
rect 16800 19600 16890 19840
rect 17130 19600 17220 19840
rect 17460 19600 17550 19840
rect 17790 19600 17880 19840
rect 18120 19600 18210 19840
rect 18450 19600 18540 19840
rect 18780 19600 18870 19840
rect 19110 19600 19200 19840
rect 19440 19600 19530 19840
rect 19770 19600 19860 19840
rect 20100 19600 20450 19840
rect 8140 19510 20450 19600
rect 8140 19270 8310 19510
rect 8550 19270 8640 19510
rect 8880 19270 8970 19510
rect 9210 19270 9300 19510
rect 9540 19270 9630 19510
rect 9870 19270 9960 19510
rect 10200 19270 10290 19510
rect 10530 19270 10620 19510
rect 10860 19270 10950 19510
rect 11190 19270 11280 19510
rect 11520 19270 11610 19510
rect 11850 19270 11940 19510
rect 12180 19270 12270 19510
rect 12510 19270 12600 19510
rect 12840 19270 12930 19510
rect 13170 19270 13260 19510
rect 13500 19270 13590 19510
rect 13830 19270 13920 19510
rect 14160 19270 14250 19510
rect 14490 19270 14580 19510
rect 14820 19270 14910 19510
rect 15150 19270 15240 19510
rect 15480 19270 15570 19510
rect 15810 19270 15900 19510
rect 16140 19270 16230 19510
rect 16470 19270 16560 19510
rect 16800 19270 16890 19510
rect 17130 19270 17220 19510
rect 17460 19270 17550 19510
rect 17790 19270 17880 19510
rect 18120 19270 18210 19510
rect 18450 19270 18540 19510
rect 18780 19270 18870 19510
rect 19110 19270 19200 19510
rect 19440 19270 19530 19510
rect 19770 19270 19860 19510
rect 20100 19270 20450 19510
rect 8140 19180 20450 19270
rect 8140 18940 8310 19180
rect 8550 18940 8640 19180
rect 8880 18940 8970 19180
rect 9210 18940 9300 19180
rect 9540 18940 9630 19180
rect 9870 18940 9960 19180
rect 10200 18940 10290 19180
rect 10530 18940 10620 19180
rect 10860 18940 10950 19180
rect 11190 18940 11280 19180
rect 11520 18940 11610 19180
rect 11850 18940 11940 19180
rect 12180 18940 12270 19180
rect 12510 18940 12600 19180
rect 12840 18940 12930 19180
rect 13170 18940 13260 19180
rect 13500 18940 13590 19180
rect 13830 18940 13920 19180
rect 14160 18940 14250 19180
rect 14490 18940 14580 19180
rect 14820 18940 14910 19180
rect 15150 18940 15240 19180
rect 15480 18940 15570 19180
rect 15810 18940 15900 19180
rect 16140 18940 16230 19180
rect 16470 18940 16560 19180
rect 16800 18940 16890 19180
rect 17130 18940 17220 19180
rect 17460 18940 17550 19180
rect 17790 18940 17880 19180
rect 18120 18940 18210 19180
rect 18450 18940 18540 19180
rect 18780 18940 18870 19180
rect 19110 18940 19200 19180
rect 19440 18940 19530 19180
rect 19770 18940 19860 19180
rect 20100 18940 20450 19180
rect 8140 18850 20450 18940
rect 8140 18610 8310 18850
rect 8550 18610 8640 18850
rect 8880 18610 8970 18850
rect 9210 18610 9300 18850
rect 9540 18610 9630 18850
rect 9870 18610 9960 18850
rect 10200 18610 10290 18850
rect 10530 18610 10620 18850
rect 10860 18610 10950 18850
rect 11190 18610 11280 18850
rect 11520 18610 11610 18850
rect 11850 18610 11940 18850
rect 12180 18610 12270 18850
rect 12510 18610 12600 18850
rect 12840 18610 12930 18850
rect 13170 18610 13260 18850
rect 13500 18610 13590 18850
rect 13830 18610 13920 18850
rect 14160 18610 14250 18850
rect 14490 18610 14580 18850
rect 14820 18610 14910 18850
rect 15150 18610 15240 18850
rect 15480 18610 15570 18850
rect 15810 18610 15900 18850
rect 16140 18610 16230 18850
rect 16470 18610 16560 18850
rect 16800 18610 16890 18850
rect 17130 18610 17220 18850
rect 17460 18610 17550 18850
rect 17790 18610 17880 18850
rect 18120 18610 18210 18850
rect 18450 18610 18540 18850
rect 18780 18610 18870 18850
rect 19110 18610 19200 18850
rect 19440 18610 19530 18850
rect 19770 18610 19860 18850
rect 20100 18610 20450 18850
rect 8140 18520 20450 18610
rect 8140 18280 8310 18520
rect 8550 18280 8640 18520
rect 8880 18280 8970 18520
rect 9210 18280 9300 18520
rect 9540 18280 9630 18520
rect 9870 18280 9960 18520
rect 10200 18280 10290 18520
rect 10530 18280 10620 18520
rect 10860 18280 10950 18520
rect 11190 18280 11280 18520
rect 11520 18280 11610 18520
rect 11850 18280 11940 18520
rect 12180 18280 12270 18520
rect 12510 18280 12600 18520
rect 12840 18280 12930 18520
rect 13170 18280 13260 18520
rect 13500 18280 13590 18520
rect 13830 18280 13920 18520
rect 14160 18280 14250 18520
rect 14490 18280 14580 18520
rect 14820 18280 14910 18520
rect 15150 18280 15240 18520
rect 15480 18280 15570 18520
rect 15810 18280 15900 18520
rect 16140 18280 16230 18520
rect 16470 18280 16560 18520
rect 16800 18280 16890 18520
rect 17130 18280 17220 18520
rect 17460 18280 17550 18520
rect 17790 18280 17880 18520
rect 18120 18280 18210 18520
rect 18450 18280 18540 18520
rect 18780 18280 18870 18520
rect 19110 18280 19200 18520
rect 19440 18280 19530 18520
rect 19770 18280 19860 18520
rect 20100 18280 20450 18520
rect 8140 18190 20450 18280
rect 8140 17950 8310 18190
rect 8550 17950 8640 18190
rect 8880 17950 8970 18190
rect 9210 17950 9300 18190
rect 9540 17950 9630 18190
rect 9870 17950 9960 18190
rect 10200 17950 10290 18190
rect 10530 17950 10620 18190
rect 10860 17950 10950 18190
rect 11190 17950 11280 18190
rect 11520 17950 11610 18190
rect 11850 17950 11940 18190
rect 12180 17950 12270 18190
rect 12510 17950 12600 18190
rect 12840 17950 12930 18190
rect 13170 17950 13260 18190
rect 13500 17950 13590 18190
rect 13830 17950 13920 18190
rect 14160 17950 14250 18190
rect 14490 17950 14580 18190
rect 14820 17950 14910 18190
rect 15150 17950 15240 18190
rect 15480 17950 15570 18190
rect 15810 17950 15900 18190
rect 16140 17950 16230 18190
rect 16470 17950 16560 18190
rect 16800 17950 16890 18190
rect 17130 17950 17220 18190
rect 17460 17950 17550 18190
rect 17790 17950 17880 18190
rect 18120 17950 18210 18190
rect 18450 17950 18540 18190
rect 18780 17950 18870 18190
rect 19110 17950 19200 18190
rect 19440 17950 19530 18190
rect 19770 17950 19860 18190
rect 20100 17950 20450 18190
rect 8140 17860 20450 17950
rect 8140 17620 8310 17860
rect 8550 17620 8640 17860
rect 8880 17620 8970 17860
rect 9210 17620 9300 17860
rect 9540 17620 9630 17860
rect 9870 17620 9960 17860
rect 10200 17620 10290 17860
rect 10530 17620 10620 17860
rect 10860 17620 10950 17860
rect 11190 17620 11280 17860
rect 11520 17620 11610 17860
rect 11850 17620 11940 17860
rect 12180 17620 12270 17860
rect 12510 17620 12600 17860
rect 12840 17620 12930 17860
rect 13170 17620 13260 17860
rect 13500 17620 13590 17860
rect 13830 17620 13920 17860
rect 14160 17620 14250 17860
rect 14490 17620 14580 17860
rect 14820 17620 14910 17860
rect 15150 17620 15240 17860
rect 15480 17620 15570 17860
rect 15810 17620 15900 17860
rect 16140 17620 16230 17860
rect 16470 17620 16560 17860
rect 16800 17620 16890 17860
rect 17130 17620 17220 17860
rect 17460 17620 17550 17860
rect 17790 17620 17880 17860
rect 18120 17620 18210 17860
rect 18450 17620 18540 17860
rect 18780 17620 18870 17860
rect 19110 17620 19200 17860
rect 19440 17620 19530 17860
rect 19770 17620 19860 17860
rect 20100 17620 20450 17860
rect 8140 17530 20450 17620
rect 8140 17290 8310 17530
rect 8550 17290 8640 17530
rect 8880 17290 8970 17530
rect 9210 17290 9300 17530
rect 9540 17290 9630 17530
rect 9870 17290 9960 17530
rect 10200 17290 10290 17530
rect 10530 17290 10620 17530
rect 10860 17290 10950 17530
rect 11190 17290 11280 17530
rect 11520 17290 11610 17530
rect 11850 17290 11940 17530
rect 12180 17290 12270 17530
rect 12510 17290 12600 17530
rect 12840 17290 12930 17530
rect 13170 17290 13260 17530
rect 13500 17290 13590 17530
rect 13830 17290 13920 17530
rect 14160 17290 14250 17530
rect 14490 17290 14580 17530
rect 14820 17290 14910 17530
rect 15150 17290 15240 17530
rect 15480 17290 15570 17530
rect 15810 17290 15900 17530
rect 16140 17290 16230 17530
rect 16470 17290 16560 17530
rect 16800 17290 16890 17530
rect 17130 17290 17220 17530
rect 17460 17290 17550 17530
rect 17790 17290 17880 17530
rect 18120 17290 18210 17530
rect 18450 17290 18540 17530
rect 18780 17290 18870 17530
rect 19110 17290 19200 17530
rect 19440 17290 19530 17530
rect 19770 17290 19860 17530
rect 20100 17290 20450 17530
rect 8140 17200 20450 17290
rect 8140 16960 8310 17200
rect 8550 16960 8640 17200
rect 8880 16960 8970 17200
rect 9210 16960 9300 17200
rect 9540 16960 9630 17200
rect 9870 16960 9960 17200
rect 10200 16960 10290 17200
rect 10530 16960 10620 17200
rect 10860 16960 10950 17200
rect 11190 16960 11280 17200
rect 11520 16960 11610 17200
rect 11850 16960 11940 17200
rect 12180 16960 12270 17200
rect 12510 16960 12600 17200
rect 12840 16960 12930 17200
rect 13170 16960 13260 17200
rect 13500 16960 13590 17200
rect 13830 16960 13920 17200
rect 14160 16960 14250 17200
rect 14490 16960 14580 17200
rect 14820 16960 14910 17200
rect 15150 16960 15240 17200
rect 15480 16960 15570 17200
rect 15810 16960 15900 17200
rect 16140 16960 16230 17200
rect 16470 16960 16560 17200
rect 16800 16960 16890 17200
rect 17130 16960 17220 17200
rect 17460 16960 17550 17200
rect 17790 16960 17880 17200
rect 18120 16960 18210 17200
rect 18450 16960 18540 17200
rect 18780 16960 18870 17200
rect 19110 16960 19200 17200
rect 19440 16960 19530 17200
rect 19770 16960 19860 17200
rect 20100 16960 20450 17200
rect 8140 16870 20450 16960
rect 8140 16630 8310 16870
rect 8550 16630 8640 16870
rect 8880 16630 8970 16870
rect 9210 16630 9300 16870
rect 9540 16630 9630 16870
rect 9870 16630 9960 16870
rect 10200 16630 10290 16870
rect 10530 16630 10620 16870
rect 10860 16630 10950 16870
rect 11190 16630 11280 16870
rect 11520 16630 11610 16870
rect 11850 16630 11940 16870
rect 12180 16630 12270 16870
rect 12510 16630 12600 16870
rect 12840 16630 12930 16870
rect 13170 16630 13260 16870
rect 13500 16630 13590 16870
rect 13830 16630 13920 16870
rect 14160 16630 14250 16870
rect 14490 16630 14580 16870
rect 14820 16630 14910 16870
rect 15150 16630 15240 16870
rect 15480 16630 15570 16870
rect 15810 16630 15900 16870
rect 16140 16630 16230 16870
rect 16470 16630 16560 16870
rect 16800 16630 16890 16870
rect 17130 16630 17220 16870
rect 17460 16630 17550 16870
rect 17790 16630 17880 16870
rect 18120 16630 18210 16870
rect 18450 16630 18540 16870
rect 18780 16630 18870 16870
rect 19110 16630 19200 16870
rect 19440 16630 19530 16870
rect 19770 16630 19860 16870
rect 20100 16630 20450 16870
rect 8140 16540 20450 16630
rect 8140 16300 8310 16540
rect 8550 16300 8640 16540
rect 8880 16300 8970 16540
rect 9210 16300 9300 16540
rect 9540 16300 9630 16540
rect 9870 16300 9960 16540
rect 10200 16300 10290 16540
rect 10530 16300 10620 16540
rect 10860 16300 10950 16540
rect 11190 16300 11280 16540
rect 11520 16300 11610 16540
rect 11850 16300 11940 16540
rect 12180 16300 12270 16540
rect 12510 16300 12600 16540
rect 12840 16300 12930 16540
rect 13170 16300 13260 16540
rect 13500 16300 13590 16540
rect 13830 16300 13920 16540
rect 14160 16300 14250 16540
rect 14490 16300 14580 16540
rect 14820 16300 14910 16540
rect 15150 16300 15240 16540
rect 15480 16300 15570 16540
rect 15810 16300 15900 16540
rect 16140 16300 16230 16540
rect 16470 16300 16560 16540
rect 16800 16300 16890 16540
rect 17130 16300 17220 16540
rect 17460 16300 17550 16540
rect 17790 16300 17880 16540
rect 18120 16300 18210 16540
rect 18450 16300 18540 16540
rect 18780 16300 18870 16540
rect 19110 16300 19200 16540
rect 19440 16300 19530 16540
rect 19770 16300 19860 16540
rect 20100 16300 20450 16540
rect 8140 16210 20450 16300
rect 8140 15970 8310 16210
rect 8550 15970 8640 16210
rect 8880 15970 8970 16210
rect 9210 15970 9300 16210
rect 9540 15970 9630 16210
rect 9870 15970 9960 16210
rect 10200 15970 10290 16210
rect 10530 15970 10620 16210
rect 10860 15970 10950 16210
rect 11190 15970 11280 16210
rect 11520 15970 11610 16210
rect 11850 15970 11940 16210
rect 12180 15970 12270 16210
rect 12510 15970 12600 16210
rect 12840 15970 12930 16210
rect 13170 15970 13260 16210
rect 13500 15970 13590 16210
rect 13830 15970 13920 16210
rect 14160 15970 14250 16210
rect 14490 15970 14580 16210
rect 14820 15970 14910 16210
rect 15150 15970 15240 16210
rect 15480 15970 15570 16210
rect 15810 15970 15900 16210
rect 16140 15970 16230 16210
rect 16470 15970 16560 16210
rect 16800 15970 16890 16210
rect 17130 15970 17220 16210
rect 17460 15970 17550 16210
rect 17790 15970 17880 16210
rect 18120 15970 18210 16210
rect 18450 15970 18540 16210
rect 18780 15970 18870 16210
rect 19110 15970 19200 16210
rect 19440 15970 19530 16210
rect 19770 15970 19860 16210
rect 20100 15970 20450 16210
rect 8140 15880 20450 15970
rect 8140 15640 8310 15880
rect 8550 15640 8640 15880
rect 8880 15640 8970 15880
rect 9210 15640 9300 15880
rect 9540 15640 9630 15880
rect 9870 15640 9960 15880
rect 10200 15640 10290 15880
rect 10530 15640 10620 15880
rect 10860 15640 10950 15880
rect 11190 15640 11280 15880
rect 11520 15640 11610 15880
rect 11850 15640 11940 15880
rect 12180 15640 12270 15880
rect 12510 15640 12600 15880
rect 12840 15640 12930 15880
rect 13170 15640 13260 15880
rect 13500 15640 13590 15880
rect 13830 15640 13920 15880
rect 14160 15640 14250 15880
rect 14490 15640 14580 15880
rect 14820 15640 14910 15880
rect 15150 15640 15240 15880
rect 15480 15640 15570 15880
rect 15810 15640 15900 15880
rect 16140 15640 16230 15880
rect 16470 15640 16560 15880
rect 16800 15640 16890 15880
rect 17130 15640 17220 15880
rect 17460 15640 17550 15880
rect 17790 15640 17880 15880
rect 18120 15640 18210 15880
rect 18450 15640 18540 15880
rect 18780 15640 18870 15880
rect 19110 15640 19200 15880
rect 19440 15640 19530 15880
rect 19770 15640 19860 15880
rect 20100 15640 20450 15880
rect 8140 15550 20450 15640
rect 8140 15310 8310 15550
rect 8550 15310 8640 15550
rect 8880 15310 8970 15550
rect 9210 15310 9300 15550
rect 9540 15310 9630 15550
rect 9870 15310 9960 15550
rect 10200 15310 10290 15550
rect 10530 15310 10620 15550
rect 10860 15310 10950 15550
rect 11190 15310 11280 15550
rect 11520 15310 11610 15550
rect 11850 15310 11940 15550
rect 12180 15310 12270 15550
rect 12510 15310 12600 15550
rect 12840 15310 12930 15550
rect 13170 15310 13260 15550
rect 13500 15310 13590 15550
rect 13830 15310 13920 15550
rect 14160 15310 14250 15550
rect 14490 15310 14580 15550
rect 14820 15310 14910 15550
rect 15150 15310 15240 15550
rect 15480 15310 15570 15550
rect 15810 15310 15900 15550
rect 16140 15310 16230 15550
rect 16470 15310 16560 15550
rect 16800 15310 16890 15550
rect 17130 15310 17220 15550
rect 17460 15310 17550 15550
rect 17790 15310 17880 15550
rect 18120 15310 18210 15550
rect 18450 15310 18540 15550
rect 18780 15310 18870 15550
rect 19110 15310 19200 15550
rect 19440 15310 19530 15550
rect 19770 15310 19860 15550
rect 20100 15310 20450 15550
rect 8140 15220 20450 15310
rect 8140 14980 8310 15220
rect 8550 14980 8640 15220
rect 8880 14980 8970 15220
rect 9210 14980 9300 15220
rect 9540 14980 9630 15220
rect 9870 14980 9960 15220
rect 10200 14980 10290 15220
rect 10530 14980 10620 15220
rect 10860 14980 10950 15220
rect 11190 14980 11280 15220
rect 11520 14980 11610 15220
rect 11850 14980 11940 15220
rect 12180 14980 12270 15220
rect 12510 14980 12600 15220
rect 12840 14980 12930 15220
rect 13170 14980 13260 15220
rect 13500 14980 13590 15220
rect 13830 14980 13920 15220
rect 14160 14980 14250 15220
rect 14490 14980 14580 15220
rect 14820 14980 14910 15220
rect 15150 14980 15240 15220
rect 15480 14980 15570 15220
rect 15810 14980 15900 15220
rect 16140 14980 16230 15220
rect 16470 14980 16560 15220
rect 16800 14980 16890 15220
rect 17130 14980 17220 15220
rect 17460 14980 17550 15220
rect 17790 14980 17880 15220
rect 18120 14980 18210 15220
rect 18450 14980 18540 15220
rect 18780 14980 18870 15220
rect 19110 14980 19200 15220
rect 19440 14980 19530 15220
rect 19770 14980 19860 15220
rect 20100 14980 20450 15220
rect 8140 14890 20450 14980
rect 8140 14650 8310 14890
rect 8550 14650 8640 14890
rect 8880 14650 8970 14890
rect 9210 14650 9300 14890
rect 9540 14650 9630 14890
rect 9870 14650 9960 14890
rect 10200 14650 10290 14890
rect 10530 14650 10620 14890
rect 10860 14650 10950 14890
rect 11190 14650 11280 14890
rect 11520 14650 11610 14890
rect 11850 14650 11940 14890
rect 12180 14650 12270 14890
rect 12510 14650 12600 14890
rect 12840 14650 12930 14890
rect 13170 14650 13260 14890
rect 13500 14650 13590 14890
rect 13830 14650 13920 14890
rect 14160 14650 14250 14890
rect 14490 14650 14580 14890
rect 14820 14650 14910 14890
rect 15150 14650 15240 14890
rect 15480 14650 15570 14890
rect 15810 14650 15900 14890
rect 16140 14650 16230 14890
rect 16470 14650 16560 14890
rect 16800 14650 16890 14890
rect 17130 14650 17220 14890
rect 17460 14650 17550 14890
rect 17790 14650 17880 14890
rect 18120 14650 18210 14890
rect 18450 14650 18540 14890
rect 18780 14650 18870 14890
rect 19110 14650 19200 14890
rect 19440 14650 19530 14890
rect 19770 14650 19860 14890
rect 20100 14650 20450 14890
rect 8140 14560 20450 14650
rect 8140 14320 8310 14560
rect 8550 14320 8640 14560
rect 8880 14320 8970 14560
rect 9210 14320 9300 14560
rect 9540 14320 9630 14560
rect 9870 14320 9960 14560
rect 10200 14320 10290 14560
rect 10530 14320 10620 14560
rect 10860 14320 10950 14560
rect 11190 14320 11280 14560
rect 11520 14320 11610 14560
rect 11850 14320 11940 14560
rect 12180 14320 12270 14560
rect 12510 14320 12600 14560
rect 12840 14320 12930 14560
rect 13170 14320 13260 14560
rect 13500 14320 13590 14560
rect 13830 14320 13920 14560
rect 14160 14320 14250 14560
rect 14490 14320 14580 14560
rect 14820 14320 14910 14560
rect 15150 14320 15240 14560
rect 15480 14320 15570 14560
rect 15810 14320 15900 14560
rect 16140 14320 16230 14560
rect 16470 14320 16560 14560
rect 16800 14320 16890 14560
rect 17130 14320 17220 14560
rect 17460 14320 17550 14560
rect 17790 14320 17880 14560
rect 18120 14320 18210 14560
rect 18450 14320 18540 14560
rect 18780 14320 18870 14560
rect 19110 14320 19200 14560
rect 19440 14320 19530 14560
rect 19770 14320 19860 14560
rect 20100 14320 20450 14560
rect 8140 14230 20450 14320
rect 8140 13990 8310 14230
rect 8550 13990 8640 14230
rect 8880 13990 8970 14230
rect 9210 13990 9300 14230
rect 9540 13990 9630 14230
rect 9870 13990 9960 14230
rect 10200 13990 10290 14230
rect 10530 13990 10620 14230
rect 10860 13990 10950 14230
rect 11190 13990 11280 14230
rect 11520 13990 11610 14230
rect 11850 13990 11940 14230
rect 12180 13990 12270 14230
rect 12510 13990 12600 14230
rect 12840 13990 12930 14230
rect 13170 13990 13260 14230
rect 13500 13990 13590 14230
rect 13830 13990 13920 14230
rect 14160 13990 14250 14230
rect 14490 13990 14580 14230
rect 14820 13990 14910 14230
rect 15150 13990 15240 14230
rect 15480 13990 15570 14230
rect 15810 13990 15900 14230
rect 16140 13990 16230 14230
rect 16470 13990 16560 14230
rect 16800 13990 16890 14230
rect 17130 13990 17220 14230
rect 17460 13990 17550 14230
rect 17790 13990 17880 14230
rect 18120 13990 18210 14230
rect 18450 13990 18540 14230
rect 18780 13990 18870 14230
rect 19110 13990 19200 14230
rect 19440 13990 19530 14230
rect 19770 13990 19860 14230
rect 20100 13990 20450 14230
rect 8140 13900 20450 13990
rect 8140 13660 8310 13900
rect 8550 13660 8640 13900
rect 8880 13660 8970 13900
rect 9210 13660 9300 13900
rect 9540 13660 9630 13900
rect 9870 13660 9960 13900
rect 10200 13660 10290 13900
rect 10530 13660 10620 13900
rect 10860 13660 10950 13900
rect 11190 13660 11280 13900
rect 11520 13660 11610 13900
rect 11850 13660 11940 13900
rect 12180 13660 12270 13900
rect 12510 13660 12600 13900
rect 12840 13660 12930 13900
rect 13170 13660 13260 13900
rect 13500 13660 13590 13900
rect 13830 13660 13920 13900
rect 14160 13660 14250 13900
rect 14490 13660 14580 13900
rect 14820 13660 14910 13900
rect 15150 13660 15240 13900
rect 15480 13660 15570 13900
rect 15810 13660 15900 13900
rect 16140 13660 16230 13900
rect 16470 13660 16560 13900
rect 16800 13660 16890 13900
rect 17130 13660 17220 13900
rect 17460 13660 17550 13900
rect 17790 13660 17880 13900
rect 18120 13660 18210 13900
rect 18450 13660 18540 13900
rect 18780 13660 18870 13900
rect 19110 13660 19200 13900
rect 19440 13660 19530 13900
rect 19770 13660 19860 13900
rect 20100 13660 20450 13900
rect 8140 13570 20450 13660
rect 8140 13330 8310 13570
rect 8550 13330 8640 13570
rect 8880 13330 8970 13570
rect 9210 13330 9300 13570
rect 9540 13330 9630 13570
rect 9870 13330 9960 13570
rect 10200 13330 10290 13570
rect 10530 13330 10620 13570
rect 10860 13330 10950 13570
rect 11190 13330 11280 13570
rect 11520 13330 11610 13570
rect 11850 13330 11940 13570
rect 12180 13330 12270 13570
rect 12510 13330 12600 13570
rect 12840 13330 12930 13570
rect 13170 13330 13260 13570
rect 13500 13330 13590 13570
rect 13830 13330 13920 13570
rect 14160 13330 14250 13570
rect 14490 13330 14580 13570
rect 14820 13330 14910 13570
rect 15150 13330 15240 13570
rect 15480 13330 15570 13570
rect 15810 13330 15900 13570
rect 16140 13330 16230 13570
rect 16470 13330 16560 13570
rect 16800 13330 16890 13570
rect 17130 13330 17220 13570
rect 17460 13330 17550 13570
rect 17790 13330 17880 13570
rect 18120 13330 18210 13570
rect 18450 13330 18540 13570
rect 18780 13330 18870 13570
rect 19110 13330 19200 13570
rect 19440 13330 19530 13570
rect 19770 13330 19860 13570
rect 20100 13330 20450 13570
rect 8140 13240 20450 13330
rect 8140 13000 8310 13240
rect 8550 13000 8640 13240
rect 8880 13000 8970 13240
rect 9210 13000 9300 13240
rect 9540 13000 9630 13240
rect 9870 13000 9960 13240
rect 10200 13000 10290 13240
rect 10530 13000 10620 13240
rect 10860 13000 10950 13240
rect 11190 13000 11280 13240
rect 11520 13000 11610 13240
rect 11850 13000 11940 13240
rect 12180 13000 12270 13240
rect 12510 13000 12600 13240
rect 12840 13000 12930 13240
rect 13170 13000 13260 13240
rect 13500 13000 13590 13240
rect 13830 13000 13920 13240
rect 14160 13000 14250 13240
rect 14490 13000 14580 13240
rect 14820 13000 14910 13240
rect 15150 13000 15240 13240
rect 15480 13000 15570 13240
rect 15810 13000 15900 13240
rect 16140 13000 16230 13240
rect 16470 13000 16560 13240
rect 16800 13000 16890 13240
rect 17130 13000 17220 13240
rect 17460 13000 17550 13240
rect 17790 13000 17880 13240
rect 18120 13000 18210 13240
rect 18450 13000 18540 13240
rect 18780 13000 18870 13240
rect 19110 13000 19200 13240
rect 19440 13000 19530 13240
rect 19770 13000 19860 13240
rect 20100 13000 20450 13240
rect 8140 12910 20450 13000
rect 8140 12670 8310 12910
rect 8550 12670 8640 12910
rect 8880 12670 8970 12910
rect 9210 12670 9300 12910
rect 9540 12670 9630 12910
rect 9870 12670 9960 12910
rect 10200 12670 10290 12910
rect 10530 12670 10620 12910
rect 10860 12670 10950 12910
rect 11190 12670 11280 12910
rect 11520 12670 11610 12910
rect 11850 12670 11940 12910
rect 12180 12670 12270 12910
rect 12510 12670 12600 12910
rect 12840 12670 12930 12910
rect 13170 12670 13260 12910
rect 13500 12670 13590 12910
rect 13830 12670 13920 12910
rect 14160 12670 14250 12910
rect 14490 12670 14580 12910
rect 14820 12670 14910 12910
rect 15150 12670 15240 12910
rect 15480 12670 15570 12910
rect 15810 12670 15900 12910
rect 16140 12670 16230 12910
rect 16470 12670 16560 12910
rect 16800 12670 16890 12910
rect 17130 12670 17220 12910
rect 17460 12670 17550 12910
rect 17790 12670 17880 12910
rect 18120 12670 18210 12910
rect 18450 12670 18540 12910
rect 18780 12670 18870 12910
rect 19110 12670 19200 12910
rect 19440 12670 19530 12910
rect 19770 12670 19860 12910
rect 20100 12670 20450 12910
rect 8140 12580 20450 12670
rect 8140 12340 8310 12580
rect 8550 12340 8640 12580
rect 8880 12340 8970 12580
rect 9210 12340 9300 12580
rect 9540 12340 9630 12580
rect 9870 12340 9960 12580
rect 10200 12340 10290 12580
rect 10530 12340 10620 12580
rect 10860 12340 10950 12580
rect 11190 12340 11280 12580
rect 11520 12340 11610 12580
rect 11850 12340 11940 12580
rect 12180 12340 12270 12580
rect 12510 12340 12600 12580
rect 12840 12340 12930 12580
rect 13170 12340 13260 12580
rect 13500 12340 13590 12580
rect 13830 12340 13920 12580
rect 14160 12340 14250 12580
rect 14490 12340 14580 12580
rect 14820 12340 14910 12580
rect 15150 12340 15240 12580
rect 15480 12340 15570 12580
rect 15810 12340 15900 12580
rect 16140 12340 16230 12580
rect 16470 12340 16560 12580
rect 16800 12340 16890 12580
rect 17130 12340 17220 12580
rect 17460 12340 17550 12580
rect 17790 12340 17880 12580
rect 18120 12340 18210 12580
rect 18450 12340 18540 12580
rect 18780 12340 18870 12580
rect 19110 12340 19200 12580
rect 19440 12340 19530 12580
rect 19770 12340 19860 12580
rect 20100 12340 20450 12580
rect 8140 12250 20450 12340
rect 8140 12010 8310 12250
rect 8550 12010 8640 12250
rect 8880 12010 8970 12250
rect 9210 12010 9300 12250
rect 9540 12010 9630 12250
rect 9870 12010 9960 12250
rect 10200 12010 10290 12250
rect 10530 12010 10620 12250
rect 10860 12010 10950 12250
rect 11190 12010 11280 12250
rect 11520 12010 11610 12250
rect 11850 12010 11940 12250
rect 12180 12010 12270 12250
rect 12510 12010 12600 12250
rect 12840 12010 12930 12250
rect 13170 12010 13260 12250
rect 13500 12010 13590 12250
rect 13830 12010 13920 12250
rect 14160 12010 14250 12250
rect 14490 12010 14580 12250
rect 14820 12010 14910 12250
rect 15150 12010 15240 12250
rect 15480 12010 15570 12250
rect 15810 12010 15900 12250
rect 16140 12010 16230 12250
rect 16470 12010 16560 12250
rect 16800 12010 16890 12250
rect 17130 12010 17220 12250
rect 17460 12010 17550 12250
rect 17790 12010 17880 12250
rect 18120 12010 18210 12250
rect 18450 12010 18540 12250
rect 18780 12010 18870 12250
rect 19110 12010 19200 12250
rect 19440 12010 19530 12250
rect 19770 12010 19860 12250
rect 20100 12010 20450 12250
rect 8140 11920 20450 12010
rect 8140 11680 8310 11920
rect 8550 11680 8640 11920
rect 8880 11680 8970 11920
rect 9210 11680 9300 11920
rect 9540 11680 9630 11920
rect 9870 11680 9960 11920
rect 10200 11680 10290 11920
rect 10530 11680 10620 11920
rect 10860 11680 10950 11920
rect 11190 11680 11280 11920
rect 11520 11680 11610 11920
rect 11850 11680 11940 11920
rect 12180 11680 12270 11920
rect 12510 11680 12600 11920
rect 12840 11680 12930 11920
rect 13170 11680 13260 11920
rect 13500 11680 13590 11920
rect 13830 11680 13920 11920
rect 14160 11680 14250 11920
rect 14490 11680 14580 11920
rect 14820 11680 14910 11920
rect 15150 11680 15240 11920
rect 15480 11680 15570 11920
rect 15810 11680 15900 11920
rect 16140 11680 16230 11920
rect 16470 11680 16560 11920
rect 16800 11680 16890 11920
rect 17130 11680 17220 11920
rect 17460 11680 17550 11920
rect 17790 11680 17880 11920
rect 18120 11680 18210 11920
rect 18450 11680 18540 11920
rect 18780 11680 18870 11920
rect 19110 11680 19200 11920
rect 19440 11680 19530 11920
rect 19770 11680 19860 11920
rect 20100 11680 20450 11920
rect 8140 11590 20450 11680
rect 8140 11350 8310 11590
rect 8550 11350 8640 11590
rect 8880 11350 8970 11590
rect 9210 11350 9300 11590
rect 9540 11350 9630 11590
rect 9870 11350 9960 11590
rect 10200 11350 10290 11590
rect 10530 11350 10620 11590
rect 10860 11350 10950 11590
rect 11190 11350 11280 11590
rect 11520 11350 11610 11590
rect 11850 11350 11940 11590
rect 12180 11350 12270 11590
rect 12510 11350 12600 11590
rect 12840 11350 12930 11590
rect 13170 11350 13260 11590
rect 13500 11350 13590 11590
rect 13830 11350 13920 11590
rect 14160 11350 14250 11590
rect 14490 11350 14580 11590
rect 14820 11350 14910 11590
rect 15150 11350 15240 11590
rect 15480 11350 15570 11590
rect 15810 11350 15900 11590
rect 16140 11350 16230 11590
rect 16470 11350 16560 11590
rect 16800 11350 16890 11590
rect 17130 11350 17220 11590
rect 17460 11350 17550 11590
rect 17790 11350 17880 11590
rect 18120 11350 18210 11590
rect 18450 11350 18540 11590
rect 18780 11350 18870 11590
rect 19110 11350 19200 11590
rect 19440 11350 19530 11590
rect 19770 11350 19860 11590
rect 20100 11350 20450 11590
rect 8140 11260 20450 11350
rect 8140 11020 8310 11260
rect 8550 11020 8640 11260
rect 8880 11020 8970 11260
rect 9210 11020 9300 11260
rect 9540 11020 9630 11260
rect 9870 11020 9960 11260
rect 10200 11020 10290 11260
rect 10530 11020 10620 11260
rect 10860 11020 10950 11260
rect 11190 11020 11280 11260
rect 11520 11020 11610 11260
rect 11850 11020 11940 11260
rect 12180 11020 12270 11260
rect 12510 11020 12600 11260
rect 12840 11020 12930 11260
rect 13170 11020 13260 11260
rect 13500 11020 13590 11260
rect 13830 11020 13920 11260
rect 14160 11020 14250 11260
rect 14490 11020 14580 11260
rect 14820 11020 14910 11260
rect 15150 11020 15240 11260
rect 15480 11020 15570 11260
rect 15810 11020 15900 11260
rect 16140 11020 16230 11260
rect 16470 11020 16560 11260
rect 16800 11020 16890 11260
rect 17130 11020 17220 11260
rect 17460 11020 17550 11260
rect 17790 11020 17880 11260
rect 18120 11020 18210 11260
rect 18450 11020 18540 11260
rect 18780 11020 18870 11260
rect 19110 11020 19200 11260
rect 19440 11020 19530 11260
rect 19770 11020 19860 11260
rect 20100 11020 20450 11260
rect 8140 10930 20450 11020
rect 8140 10690 8310 10930
rect 8550 10690 8640 10930
rect 8880 10690 8970 10930
rect 9210 10690 9300 10930
rect 9540 10690 9630 10930
rect 9870 10690 9960 10930
rect 10200 10690 10290 10930
rect 10530 10690 10620 10930
rect 10860 10690 10950 10930
rect 11190 10690 11280 10930
rect 11520 10690 11610 10930
rect 11850 10690 11940 10930
rect 12180 10690 12270 10930
rect 12510 10690 12600 10930
rect 12840 10690 12930 10930
rect 13170 10690 13260 10930
rect 13500 10690 13590 10930
rect 13830 10690 13920 10930
rect 14160 10690 14250 10930
rect 14490 10690 14580 10930
rect 14820 10690 14910 10930
rect 15150 10690 15240 10930
rect 15480 10690 15570 10930
rect 15810 10690 15900 10930
rect 16140 10690 16230 10930
rect 16470 10690 16560 10930
rect 16800 10690 16890 10930
rect 17130 10690 17220 10930
rect 17460 10690 17550 10930
rect 17790 10690 17880 10930
rect 18120 10690 18210 10930
rect 18450 10690 18540 10930
rect 18780 10690 18870 10930
rect 19110 10690 19200 10930
rect 19440 10690 19530 10930
rect 19770 10690 19860 10930
rect 20100 10690 20450 10930
rect 8140 10600 20450 10690
rect 8140 10360 8310 10600
rect 8550 10360 8640 10600
rect 8880 10360 8970 10600
rect 9210 10360 9300 10600
rect 9540 10360 9630 10600
rect 9870 10360 9960 10600
rect 10200 10360 10290 10600
rect 10530 10360 10620 10600
rect 10860 10360 10950 10600
rect 11190 10360 11280 10600
rect 11520 10360 11610 10600
rect 11850 10360 11940 10600
rect 12180 10360 12270 10600
rect 12510 10360 12600 10600
rect 12840 10360 12930 10600
rect 13170 10360 13260 10600
rect 13500 10360 13590 10600
rect 13830 10360 13920 10600
rect 14160 10360 14250 10600
rect 14490 10360 14580 10600
rect 14820 10360 14910 10600
rect 15150 10360 15240 10600
rect 15480 10360 15570 10600
rect 15810 10360 15900 10600
rect 16140 10360 16230 10600
rect 16470 10360 16560 10600
rect 16800 10360 16890 10600
rect 17130 10360 17220 10600
rect 17460 10360 17550 10600
rect 17790 10360 17880 10600
rect 18120 10360 18210 10600
rect 18450 10360 18540 10600
rect 18780 10360 18870 10600
rect 19110 10360 19200 10600
rect 19440 10360 19530 10600
rect 19770 10360 19860 10600
rect 20100 10360 20450 10600
rect 8140 10270 20450 10360
rect 8140 10030 8310 10270
rect 8550 10030 8640 10270
rect 8880 10030 8970 10270
rect 9210 10030 9300 10270
rect 9540 10030 9630 10270
rect 9870 10030 9960 10270
rect 10200 10030 10290 10270
rect 10530 10030 10620 10270
rect 10860 10030 10950 10270
rect 11190 10030 11280 10270
rect 11520 10030 11610 10270
rect 11850 10030 11940 10270
rect 12180 10030 12270 10270
rect 12510 10030 12600 10270
rect 12840 10030 12930 10270
rect 13170 10030 13260 10270
rect 13500 10030 13590 10270
rect 13830 10030 13920 10270
rect 14160 10030 14250 10270
rect 14490 10030 14580 10270
rect 14820 10030 14910 10270
rect 15150 10030 15240 10270
rect 15480 10030 15570 10270
rect 15810 10030 15900 10270
rect 16140 10030 16230 10270
rect 16470 10030 16560 10270
rect 16800 10030 16890 10270
rect 17130 10030 17220 10270
rect 17460 10030 17550 10270
rect 17790 10030 17880 10270
rect 18120 10030 18210 10270
rect 18450 10030 18540 10270
rect 18780 10030 18870 10270
rect 19110 10030 19200 10270
rect 19440 10030 19530 10270
rect 19770 10030 19860 10270
rect 20100 10030 20450 10270
rect 8140 9940 20450 10030
rect 8140 9700 8310 9940
rect 8550 9700 8640 9940
rect 8880 9700 8970 9940
rect 9210 9700 9300 9940
rect 9540 9700 9630 9940
rect 9870 9700 9960 9940
rect 10200 9700 10290 9940
rect 10530 9700 10620 9940
rect 10860 9700 10950 9940
rect 11190 9700 11280 9940
rect 11520 9700 11610 9940
rect 11850 9700 11940 9940
rect 12180 9700 12270 9940
rect 12510 9700 12600 9940
rect 12840 9700 12930 9940
rect 13170 9700 13260 9940
rect 13500 9700 13590 9940
rect 13830 9700 13920 9940
rect 14160 9700 14250 9940
rect 14490 9700 14580 9940
rect 14820 9700 14910 9940
rect 15150 9700 15240 9940
rect 15480 9700 15570 9940
rect 15810 9700 15900 9940
rect 16140 9700 16230 9940
rect 16470 9700 16560 9940
rect 16800 9700 16890 9940
rect 17130 9700 17220 9940
rect 17460 9700 17550 9940
rect 17790 9700 17880 9940
rect 18120 9700 18210 9940
rect 18450 9700 18540 9940
rect 18780 9700 18870 9940
rect 19110 9700 19200 9940
rect 19440 9700 19530 9940
rect 19770 9700 19860 9940
rect 20100 9700 20450 9940
rect 8140 9610 20450 9700
rect 8140 9370 8310 9610
rect 8550 9370 8640 9610
rect 8880 9370 8970 9610
rect 9210 9370 9300 9610
rect 9540 9370 9630 9610
rect 9870 9370 9960 9610
rect 10200 9370 10290 9610
rect 10530 9370 10620 9610
rect 10860 9370 10950 9610
rect 11190 9370 11280 9610
rect 11520 9370 11610 9610
rect 11850 9370 11940 9610
rect 12180 9370 12270 9610
rect 12510 9370 12600 9610
rect 12840 9370 12930 9610
rect 13170 9370 13260 9610
rect 13500 9370 13590 9610
rect 13830 9370 13920 9610
rect 14160 9370 14250 9610
rect 14490 9370 14580 9610
rect 14820 9370 14910 9610
rect 15150 9370 15240 9610
rect 15480 9370 15570 9610
rect 15810 9370 15900 9610
rect 16140 9370 16230 9610
rect 16470 9370 16560 9610
rect 16800 9370 16890 9610
rect 17130 9370 17220 9610
rect 17460 9370 17550 9610
rect 17790 9370 17880 9610
rect 18120 9370 18210 9610
rect 18450 9370 18540 9610
rect 18780 9370 18870 9610
rect 19110 9370 19200 9610
rect 19440 9370 19530 9610
rect 19770 9370 19860 9610
rect 20100 9370 20450 9610
rect 8140 9280 20450 9370
rect 8140 9040 8310 9280
rect 8550 9040 8640 9280
rect 8880 9040 8970 9280
rect 9210 9040 9300 9280
rect 9540 9040 9630 9280
rect 9870 9040 9960 9280
rect 10200 9040 10290 9280
rect 10530 9040 10620 9280
rect 10860 9040 10950 9280
rect 11190 9040 11280 9280
rect 11520 9040 11610 9280
rect 11850 9040 11940 9280
rect 12180 9040 12270 9280
rect 12510 9040 12600 9280
rect 12840 9040 12930 9280
rect 13170 9040 13260 9280
rect 13500 9040 13590 9280
rect 13830 9040 13920 9280
rect 14160 9040 14250 9280
rect 14490 9040 14580 9280
rect 14820 9040 14910 9280
rect 15150 9040 15240 9280
rect 15480 9040 15570 9280
rect 15810 9040 15900 9280
rect 16140 9040 16230 9280
rect 16470 9040 16560 9280
rect 16800 9040 16890 9280
rect 17130 9040 17220 9280
rect 17460 9040 17550 9280
rect 17790 9040 17880 9280
rect 18120 9040 18210 9280
rect 18450 9040 18540 9280
rect 18780 9040 18870 9280
rect 19110 9040 19200 9280
rect 19440 9040 19530 9280
rect 19770 9040 19860 9280
rect 20100 9040 20450 9280
rect 8140 8690 20450 9040
rect 8140 8410 8460 8690
rect 8140 8340 8180 8410
rect 8250 8340 8270 8410
rect 8340 8340 8360 8410
rect 8430 8340 8460 8410
rect 8140 8320 8460 8340
rect 8140 8250 8180 8320
rect 8250 8250 8270 8320
rect 8340 8250 8360 8320
rect 8430 8250 8460 8320
rect 8140 8230 8460 8250
rect 11760 6940 13360 6960
rect 1540 6910 3140 6930
rect 1540 6850 1720 6910
rect 1960 6850 2050 6910
rect 2290 6850 2390 6910
rect 2630 6850 2720 6910
rect 2960 6850 3140 6910
rect 1540 6780 1570 6850
rect 1640 6780 1680 6850
rect 1970 6780 2010 6850
rect 2300 6780 2340 6850
rect 2630 6780 2670 6850
rect 2960 6780 3000 6850
rect 3070 6780 3140 6850
rect 1540 6740 1720 6780
rect 1960 6740 2050 6780
rect 2290 6740 2390 6780
rect 2630 6740 2720 6780
rect 2960 6740 3140 6780
rect 1540 6670 1570 6740
rect 1640 6670 1680 6740
rect 1970 6670 2010 6740
rect 2300 6670 2340 6740
rect 2630 6670 2670 6740
rect 2960 6670 3000 6740
rect 3070 6670 3140 6740
rect 11760 6880 11940 6940
rect 12180 6880 12270 6940
rect 12510 6880 12610 6940
rect 12850 6880 12940 6940
rect 13180 6880 13360 6940
rect 11760 6810 11790 6880
rect 11860 6810 11900 6880
rect 12190 6810 12230 6880
rect 12520 6810 12560 6880
rect 12850 6810 12890 6880
rect 13180 6810 13220 6880
rect 13290 6810 13360 6880
rect 11760 6770 11940 6810
rect 12180 6770 12270 6810
rect 12510 6770 12610 6810
rect 12850 6770 12940 6810
rect 13180 6770 13360 6810
rect 11760 6700 11790 6770
rect 11860 6700 11900 6770
rect 12190 6700 12230 6770
rect 12520 6700 12560 6770
rect 12850 6700 12890 6770
rect 13180 6700 13220 6770
rect 13290 6700 13360 6770
rect 11760 6670 13360 6700
rect 1540 6640 3140 6670
rect 7400 5390 7490 5410
rect 7400 5320 7410 5390
rect 7480 5320 7490 5390
rect 7400 5280 7490 5320
rect 7400 5240 7410 5280
rect -2870 5210 7410 5240
rect 7480 5240 7490 5280
rect 21120 5240 21280 8880
rect 7480 5210 21280 5240
rect -2870 5170 21280 5210
rect -2870 5100 7410 5170
rect 7480 5100 21280 5170
rect -2870 5080 21280 5100
rect 21800 8230 39650 8490
rect 21800 5670 22060 8230
rect 31100 7830 37860 7910
rect 31100 7590 31180 7830
rect 31420 7590 31510 7830
rect 31750 7590 31840 7830
rect 32080 7590 32170 7830
rect 32410 7590 32500 7830
rect 32740 7590 32830 7830
rect 33070 7590 33160 7830
rect 33400 7590 33490 7830
rect 33730 7590 33820 7830
rect 34060 7590 34150 7830
rect 34390 7590 34480 7830
rect 34720 7590 34810 7830
rect 35050 7590 35140 7830
rect 35380 7590 35470 7830
rect 35710 7590 35800 7830
rect 36040 7590 36130 7830
rect 36370 7590 36460 7830
rect 36700 7590 36790 7830
rect 37030 7590 37120 7830
rect 37360 7590 37450 7830
rect 37690 7590 37860 7830
rect 31100 7500 37860 7590
rect 23460 7270 23940 7290
rect 23460 7210 23510 7270
rect 23880 7210 23940 7270
rect 23460 7140 23490 7210
rect 23890 7140 23940 7210
rect 23460 7100 23510 7140
rect 23880 7100 23940 7140
rect 23460 7030 23490 7100
rect 23890 7030 23940 7100
rect 23460 7000 23940 7030
rect 25860 7270 26340 7290
rect 25860 7210 25910 7270
rect 26280 7210 26340 7270
rect 25860 7140 25890 7210
rect 26290 7140 26340 7210
rect 25860 7100 25910 7140
rect 26280 7100 26340 7140
rect 25860 7030 25890 7100
rect 26290 7030 26340 7100
rect 25860 7000 26340 7030
rect 31100 7260 31180 7500
rect 31420 7260 31510 7500
rect 31750 7260 31840 7500
rect 32080 7260 32170 7500
rect 32410 7260 32500 7500
rect 32740 7260 32830 7500
rect 33070 7260 33160 7500
rect 33400 7260 33490 7500
rect 33730 7260 33820 7500
rect 34060 7260 34150 7500
rect 34390 7260 34480 7500
rect 34720 7260 34810 7500
rect 35050 7260 35140 7500
rect 35380 7260 35470 7500
rect 35710 7260 35800 7500
rect 36040 7260 36130 7500
rect 36370 7260 36460 7500
rect 36700 7260 36790 7500
rect 37030 7260 37120 7500
rect 37360 7260 37450 7500
rect 37690 7260 37860 7500
rect 31100 7170 37860 7260
rect 31100 6930 31180 7170
rect 31420 6930 31510 7170
rect 31750 6930 31840 7170
rect 32080 6930 32170 7170
rect 32410 6930 32500 7170
rect 32740 6930 32830 7170
rect 33070 6930 33160 7170
rect 33400 6930 33490 7170
rect 33730 6930 33820 7170
rect 34060 6930 34150 7170
rect 34390 6930 34480 7170
rect 34720 6930 34810 7170
rect 35050 6930 35140 7170
rect 35380 6930 35470 7170
rect 35710 6930 35800 7170
rect 36040 6930 36130 7170
rect 36370 6930 36460 7170
rect 36700 6930 36790 7170
rect 37030 6930 37120 7170
rect 37360 6930 37450 7170
rect 37690 6930 37860 7170
rect 31100 6840 37860 6930
rect 31100 6600 31180 6840
rect 31420 6600 31510 6840
rect 31750 6600 31840 6840
rect 32080 6600 32170 6840
rect 32410 6600 32500 6840
rect 32740 6600 32830 6840
rect 33070 6600 33160 6840
rect 33400 6600 33490 6840
rect 33730 6600 33820 6840
rect 34060 6600 34150 6840
rect 34390 6600 34480 6840
rect 34720 6600 34810 6840
rect 35050 6600 35140 6840
rect 35380 6600 35470 6840
rect 35710 6600 35800 6840
rect 36040 6600 36130 6840
rect 36370 6600 36460 6840
rect 36700 6600 36790 6840
rect 37030 6600 37120 6840
rect 37360 6600 37450 6840
rect 37690 6600 37860 6840
rect 31100 6510 37860 6600
rect 31100 6320 31180 6510
rect 30720 6300 31180 6320
rect 30720 6230 30740 6300
rect 30810 6230 30850 6300
rect 30920 6270 31180 6300
rect 31420 6270 31510 6510
rect 31750 6270 31840 6510
rect 32080 6270 32170 6510
rect 32410 6270 32500 6510
rect 32740 6270 32830 6510
rect 33070 6270 33160 6510
rect 33400 6270 33490 6510
rect 33730 6270 33820 6510
rect 34060 6270 34150 6510
rect 34390 6270 34480 6510
rect 34720 6270 34810 6510
rect 35050 6270 35140 6510
rect 35380 6270 35470 6510
rect 35710 6270 35800 6510
rect 36040 6270 36130 6510
rect 36370 6270 36460 6510
rect 36700 6270 36790 6510
rect 37030 6270 37120 6510
rect 37360 6270 37450 6510
rect 37690 6270 37860 6510
rect 30920 6230 37860 6270
rect 30720 6180 37860 6230
rect 30720 6170 31180 6180
rect 30720 6100 30740 6170
rect 30810 6100 30850 6170
rect 30920 6100 31180 6170
rect 30720 6040 31180 6100
rect 30720 5970 30740 6040
rect 30810 5970 30850 6040
rect 30920 5970 31180 6040
rect 30720 5950 31180 5970
rect 21800 5600 21820 5670
rect 21890 5600 21930 5670
rect 22000 5600 22060 5670
rect 21800 5560 22060 5600
rect 21800 5490 21820 5560
rect 21890 5490 21930 5560
rect 22000 5490 22060 5560
rect 21800 5450 22060 5490
rect 21800 5380 21820 5450
rect 21890 5380 21930 5450
rect 22000 5380 22060 5450
rect 21800 5340 22060 5380
rect 21800 5270 21820 5340
rect 21890 5270 21930 5340
rect 22000 5270 22060 5340
rect 21800 5230 22060 5270
rect 21800 5160 21820 5230
rect 21890 5160 21930 5230
rect 22000 5160 22060 5230
rect 21800 5120 22060 5160
rect 7400 5060 7490 5080
rect 7400 4990 7410 5060
rect 7480 4990 7490 5060
rect 7400 4950 7490 4990
rect 7400 4880 7410 4950
rect 7480 4880 7490 4950
rect 7400 4860 7490 4880
rect 1080 -790 2680 -760
rect 1080 -860 1150 -790
rect 1220 -860 1260 -790
rect 1550 -860 1590 -790
rect 1880 -860 1920 -790
rect 2210 -860 2250 -790
rect 2540 -860 2580 -790
rect 2650 -860 2680 -790
rect 1080 -900 1260 -860
rect 1500 -900 1590 -860
rect 1830 -900 1930 -860
rect 2170 -900 2260 -860
rect 2500 -900 2680 -860
rect 1080 -970 1150 -900
rect 1220 -970 1260 -900
rect 1550 -970 1590 -900
rect 1880 -970 1920 -900
rect 2210 -970 2250 -900
rect 2540 -970 2580 -900
rect 2650 -970 2680 -900
rect 1080 -1030 1260 -970
rect 1500 -1030 1590 -970
rect 1830 -1030 1930 -970
rect 2170 -1030 2260 -970
rect 2500 -1030 2680 -970
rect 1080 -1050 2680 -1030
rect 12220 -790 13820 -760
rect 12220 -860 12250 -790
rect 12320 -860 12360 -790
rect 12650 -860 12690 -790
rect 12980 -860 13020 -790
rect 13310 -860 13350 -790
rect 13640 -860 13680 -790
rect 13750 -860 13820 -790
rect 12220 -900 12400 -860
rect 12640 -900 12730 -860
rect 12970 -900 13070 -860
rect 13310 -900 13400 -860
rect 13640 -900 13820 -860
rect 12220 -970 12250 -900
rect 12320 -970 12360 -900
rect 12650 -970 12690 -900
rect 12980 -970 13020 -900
rect 13310 -970 13350 -900
rect 13640 -970 13680 -900
rect 13750 -970 13820 -900
rect 12220 -1030 12400 -970
rect 12640 -1030 12730 -970
rect 12970 -1030 13070 -970
rect 13310 -1030 13400 -970
rect 13640 -1030 13820 -970
rect 12220 -1050 13820 -1030
rect 1540 -2720 3140 -2700
rect 1540 -2780 1720 -2720
rect 1960 -2780 2050 -2720
rect 2290 -2780 2390 -2720
rect 2630 -2780 2720 -2720
rect 2960 -2780 3140 -2720
rect 1540 -2850 1570 -2780
rect 1640 -2850 1680 -2780
rect 1970 -2850 2010 -2780
rect 2300 -2850 2340 -2780
rect 2630 -2850 2670 -2780
rect 2960 -2850 3000 -2780
rect 3070 -2850 3140 -2780
rect 1540 -2890 1720 -2850
rect 1960 -2890 2050 -2850
rect 2290 -2890 2390 -2850
rect 2630 -2890 2720 -2850
rect 2960 -2890 3140 -2850
rect 1540 -2960 1570 -2890
rect 1640 -2960 1680 -2890
rect 1970 -2960 2010 -2890
rect 2300 -2960 2340 -2890
rect 2630 -2960 2670 -2890
rect 2960 -2960 3000 -2890
rect 3070 -2960 3140 -2890
rect 1540 -2990 3140 -2960
rect 11760 -2720 13360 -2700
rect 11760 -2780 11940 -2720
rect 12180 -2780 12270 -2720
rect 12510 -2780 12610 -2720
rect 12850 -2780 12940 -2720
rect 13180 -2780 13360 -2720
rect 11760 -2850 11790 -2780
rect 11860 -2850 11900 -2780
rect 12190 -2850 12230 -2780
rect 12520 -2850 12560 -2780
rect 12850 -2850 12890 -2780
rect 13180 -2850 13220 -2780
rect 13290 -2850 13360 -2780
rect 11760 -2890 11940 -2850
rect 12180 -2890 12270 -2850
rect 12510 -2890 12610 -2850
rect 12850 -2890 12940 -2850
rect 13180 -2890 13360 -2850
rect 11760 -2960 11790 -2890
rect 11860 -2960 11900 -2890
rect 12190 -2960 12230 -2890
rect 12520 -2960 12560 -2890
rect 12850 -2960 12890 -2890
rect 13180 -2960 13220 -2890
rect 13290 -2960 13360 -2890
rect 11760 -2990 13360 -2960
rect 7290 -3880 7620 -3860
rect 7290 -3920 7310 -3880
rect -2570 -3950 7310 -3920
rect 7380 -3950 7420 -3880
rect 7490 -3950 7530 -3880
rect 7600 -3920 7620 -3880
rect 18500 -3920 18660 5080
rect 21800 5050 21820 5120
rect 21890 5050 21930 5120
rect 22000 5050 22060 5120
rect 21800 5010 22060 5050
rect 21800 4940 21820 5010
rect 21890 4940 21930 5010
rect 22000 4940 22060 5010
rect 21800 4900 22060 4940
rect 21800 4830 21820 4900
rect 21890 4830 21930 4900
rect 22000 4830 22060 4900
rect 21800 4790 22060 4830
rect 21800 4720 21820 4790
rect 21890 4720 21930 4790
rect 22000 4720 22060 4790
rect 21800 4680 22060 4720
rect 21800 4610 21820 4680
rect 21890 4610 21930 4680
rect 22000 4610 22060 4680
rect 21800 4570 22060 4610
rect 21800 4500 21820 4570
rect 21890 4500 21930 4570
rect 22000 4500 22060 4570
rect 7600 -3950 18660 -3920
rect -2570 -3990 18660 -3950
rect -2570 -4060 7310 -3990
rect 7380 -4060 7420 -3990
rect 7490 -4060 7530 -3990
rect 7600 -4060 18660 -3990
rect -2570 -4080 18660 -4060
rect 18975 1160 19085 1180
rect 18975 1090 18995 1160
rect 19065 1090 19085 1160
rect 18975 1050 19085 1090
rect 18975 980 18995 1050
rect 19065 980 19085 1050
rect 18975 940 19085 980
rect 18975 870 18995 940
rect 19065 870 19085 940
rect 7290 -4100 7620 -4080
rect 7290 -4170 7310 -4100
rect 7380 -4170 7420 -4100
rect 7490 -4170 7530 -4100
rect 7600 -4170 7620 -4100
rect 7290 -4190 7620 -4170
rect -1350 -4350 -870 -4270
rect -1350 -4420 -1330 -4350
rect -1260 -4420 -1220 -4350
rect -1150 -4420 -1110 -4350
rect -1040 -4420 -1000 -4350
rect -930 -4420 -870 -4350
rect -1350 -4460 -870 -4420
rect -1350 -4530 -1330 -4460
rect -1260 -4530 -1220 -4460
rect -1150 -4530 -1110 -4460
rect -1040 -4530 -1000 -4460
rect -930 -4530 -870 -4460
rect -1350 -4630 -870 -4530
rect 15650 -4350 16130 -4270
rect 15650 -4420 15710 -4350
rect 15780 -4420 15820 -4350
rect 15890 -4420 15930 -4350
rect 16000 -4420 16040 -4350
rect 16110 -4420 16130 -4350
rect 15650 -4460 16130 -4420
rect 15650 -4530 15710 -4460
rect 15780 -4530 15820 -4460
rect 15890 -4530 15930 -4460
rect 16000 -4530 16040 -4460
rect 16110 -4530 16130 -4460
rect 15650 -4630 16130 -4530
rect -1350 -4840 260 -4630
rect -1350 -5080 -1180 -4840
rect -940 -5080 -850 -4840
rect -610 -5080 -520 -4840
rect -280 -5080 -190 -4840
rect 50 -5080 260 -4840
rect -1350 -5170 260 -5080
rect -1350 -5410 -1180 -5170
rect -940 -5410 -850 -5170
rect -610 -5410 -520 -5170
rect -280 -5410 -190 -5170
rect 50 -5410 260 -5170
rect -1350 -5500 260 -5410
rect -1350 -5740 -1180 -5500
rect -940 -5740 -850 -5500
rect -610 -5740 -520 -5500
rect -280 -5740 -190 -5500
rect 50 -5740 260 -5500
rect -1350 -5830 260 -5740
rect -1350 -6070 -1180 -5830
rect -940 -6070 -850 -5830
rect -610 -6070 -520 -5830
rect -280 -6070 -190 -5830
rect 50 -6070 260 -5830
rect -1350 -6240 260 -6070
rect 14520 -4840 16130 -4630
rect 14520 -5080 14730 -4840
rect 14970 -5080 15060 -4840
rect 15300 -5080 15390 -4840
rect 15630 -5080 15720 -4840
rect 15960 -5080 16130 -4840
rect 14520 -5170 16130 -5080
rect 14520 -5410 14730 -5170
rect 14970 -5410 15060 -5170
rect 15300 -5410 15390 -5170
rect 15630 -5410 15720 -5170
rect 15960 -5410 16130 -5170
rect 14520 -5500 16130 -5410
rect 14520 -5740 14730 -5500
rect 14970 -5740 15060 -5500
rect 15300 -5740 15390 -5500
rect 15630 -5740 15720 -5500
rect 15960 -5740 16130 -5500
rect 14520 -5830 16130 -5740
rect 14520 -6070 14730 -5830
rect 14970 -6070 15060 -5830
rect 15300 -6070 15390 -5830
rect 15630 -6070 15720 -5830
rect 15960 -6070 16130 -5830
rect 14520 -6240 16130 -6070
rect 18975 -5915 19085 870
rect 21800 -850 22060 4500
rect 31100 5940 31180 5950
rect 31420 5940 31510 6180
rect 31750 5940 31840 6180
rect 32080 5940 32170 6180
rect 32410 5940 32500 6180
rect 32740 5940 32830 6180
rect 33070 5940 33160 6180
rect 33400 5940 33490 6180
rect 33730 5940 33820 6180
rect 34060 5940 34150 6180
rect 34390 5940 34480 6180
rect 34720 5940 34810 6180
rect 35050 5940 35140 6180
rect 35380 5940 35470 6180
rect 35710 5940 35800 6180
rect 36040 5940 36130 6180
rect 36370 5940 36460 6180
rect 36700 5940 36790 6180
rect 37030 5940 37120 6180
rect 37360 5940 37450 6180
rect 37690 5940 37860 6180
rect 31100 5850 37860 5940
rect 31100 5610 31180 5850
rect 31420 5610 31510 5850
rect 31750 5610 31840 5850
rect 32080 5610 32170 5850
rect 32410 5610 32500 5850
rect 32740 5610 32830 5850
rect 33070 5610 33160 5850
rect 33400 5610 33490 5850
rect 33730 5610 33820 5850
rect 34060 5610 34150 5850
rect 34390 5610 34480 5850
rect 34720 5610 34810 5850
rect 35050 5610 35140 5850
rect 35380 5610 35470 5850
rect 35710 5610 35800 5850
rect 36040 5610 36130 5850
rect 36370 5610 36460 5850
rect 36700 5610 36790 5850
rect 37030 5610 37120 5850
rect 37360 5610 37450 5850
rect 37690 5610 37860 5850
rect 31100 5520 37860 5610
rect 31100 5280 31180 5520
rect 31420 5280 31510 5520
rect 31750 5280 31840 5520
rect 32080 5280 32170 5520
rect 32410 5280 32500 5520
rect 32740 5280 32830 5520
rect 33070 5280 33160 5520
rect 33400 5280 33490 5520
rect 33730 5280 33820 5520
rect 34060 5280 34150 5520
rect 34390 5280 34480 5520
rect 34720 5280 34810 5520
rect 35050 5280 35140 5520
rect 35380 5280 35470 5520
rect 35710 5280 35800 5520
rect 36040 5280 36130 5520
rect 36370 5280 36460 5520
rect 36700 5280 36790 5520
rect 37030 5280 37120 5520
rect 37360 5280 37450 5520
rect 37690 5280 37860 5520
rect 31100 5190 37860 5280
rect 31100 4950 31180 5190
rect 31420 4950 31510 5190
rect 31750 4950 31840 5190
rect 32080 4950 32170 5190
rect 32410 4950 32500 5190
rect 32740 4950 32830 5190
rect 33070 4950 33160 5190
rect 33400 4950 33490 5190
rect 33730 4950 33820 5190
rect 34060 4950 34150 5190
rect 34390 4950 34480 5190
rect 34720 4950 34810 5190
rect 35050 4950 35140 5190
rect 35380 4950 35470 5190
rect 35710 4950 35800 5190
rect 36040 4950 36130 5190
rect 36370 4950 36460 5190
rect 36700 4950 36790 5190
rect 37030 4950 37120 5190
rect 37360 4950 37450 5190
rect 37690 4950 37860 5190
rect 31100 4860 37860 4950
rect 31100 4620 31180 4860
rect 31420 4620 31510 4860
rect 31750 4620 31840 4860
rect 32080 4620 32170 4860
rect 32410 4620 32500 4860
rect 32740 4620 32830 4860
rect 33070 4620 33160 4860
rect 33400 4620 33490 4860
rect 33730 4620 33820 4860
rect 34060 4620 34150 4860
rect 34390 4620 34480 4860
rect 34720 4620 34810 4860
rect 35050 4620 35140 4860
rect 35380 4620 35470 4860
rect 35710 4620 35800 4860
rect 36040 4620 36130 4860
rect 36370 4620 36460 4860
rect 36700 4620 36790 4860
rect 37030 4620 37120 4860
rect 37360 4620 37450 4860
rect 37690 4620 37860 4860
rect 31100 4530 37860 4620
rect 31100 4290 31180 4530
rect 31420 4290 31510 4530
rect 31750 4290 31840 4530
rect 32080 4290 32170 4530
rect 32410 4290 32500 4530
rect 32740 4290 32830 4530
rect 33070 4290 33160 4530
rect 33400 4290 33490 4530
rect 33730 4290 33820 4530
rect 34060 4290 34150 4530
rect 34390 4290 34480 4530
rect 34720 4290 34810 4530
rect 35050 4290 35140 4530
rect 35380 4290 35470 4530
rect 35710 4290 35800 4530
rect 36040 4290 36130 4530
rect 36370 4290 36460 4530
rect 36700 4290 36790 4530
rect 37030 4290 37120 4530
rect 37360 4290 37450 4530
rect 37690 4290 37860 4530
rect 31100 4200 37860 4290
rect 31100 3960 31180 4200
rect 31420 3960 31510 4200
rect 31750 3960 31840 4200
rect 32080 3960 32170 4200
rect 32410 3960 32500 4200
rect 32740 3960 32830 4200
rect 33070 3960 33160 4200
rect 33400 3960 33490 4200
rect 33730 3960 33820 4200
rect 34060 3960 34150 4200
rect 34390 3960 34480 4200
rect 34720 3960 34810 4200
rect 35050 3960 35140 4200
rect 35380 3960 35470 4200
rect 35710 3960 35800 4200
rect 36040 3960 36130 4200
rect 36370 3960 36460 4200
rect 36700 3960 36790 4200
rect 37030 3960 37120 4200
rect 37360 3960 37450 4200
rect 37690 3960 37860 4200
rect 31100 3870 37860 3960
rect 31100 3630 31180 3870
rect 31420 3630 31510 3870
rect 31750 3630 31840 3870
rect 32080 3630 32170 3870
rect 32410 3630 32500 3870
rect 32740 3630 32830 3870
rect 33070 3630 33160 3870
rect 33400 3630 33490 3870
rect 33730 3630 33820 3870
rect 34060 3630 34150 3870
rect 34390 3630 34480 3870
rect 34720 3630 34810 3870
rect 35050 3630 35140 3870
rect 35380 3630 35470 3870
rect 35710 3630 35800 3870
rect 36040 3630 36130 3870
rect 36370 3630 36460 3870
rect 36700 3630 36790 3870
rect 37030 3630 37120 3870
rect 37360 3630 37450 3870
rect 37690 3630 37860 3870
rect 31100 3540 37860 3630
rect 24700 3360 25030 3380
rect 24700 3290 24720 3360
rect 24790 3290 24830 3360
rect 24900 3290 24940 3360
rect 25010 3290 25030 3360
rect 24700 3250 25030 3290
rect 24700 3236 24720 3250
rect 24684 3180 24720 3236
rect 24790 3180 24830 3250
rect 24900 3180 24940 3250
rect 25010 3236 25030 3250
rect 31100 3300 31180 3540
rect 31420 3300 31510 3540
rect 31750 3300 31840 3540
rect 32080 3300 32170 3540
rect 32410 3300 32500 3540
rect 32740 3300 32830 3540
rect 33070 3300 33160 3540
rect 33400 3300 33490 3540
rect 33730 3300 33820 3540
rect 34060 3300 34150 3540
rect 34390 3300 34480 3540
rect 34720 3300 34810 3540
rect 35050 3300 35140 3540
rect 35380 3300 35470 3540
rect 35710 3300 35800 3540
rect 36040 3300 36130 3540
rect 36370 3300 36460 3540
rect 36700 3300 36790 3540
rect 37030 3300 37120 3540
rect 37360 3300 37450 3540
rect 37690 3300 37860 3540
rect 25010 3180 30477 3236
rect 24684 3140 30477 3180
rect 24684 3103 24720 3140
rect 24700 3070 24720 3103
rect 24790 3070 24830 3140
rect 24900 3070 24940 3140
rect 25010 3103 30477 3140
rect 25010 3070 25030 3103
rect 24700 3050 25030 3070
rect 22420 2600 22900 2630
rect 22420 2530 22470 2600
rect 22870 2530 22900 2600
rect 22420 2490 22480 2530
rect 22850 2490 22900 2530
rect 22420 2420 22470 2490
rect 22870 2420 22900 2490
rect 22420 2360 22480 2420
rect 22850 2360 22900 2420
rect 22420 2340 22900 2360
rect 26900 2600 27380 2630
rect 26900 2530 26950 2600
rect 27350 2530 27380 2600
rect 26900 2490 26960 2530
rect 27330 2490 27380 2530
rect 26900 2420 26950 2490
rect 27350 2420 27380 2490
rect 26900 2360 26960 2420
rect 27330 2360 27380 2420
rect 26900 2340 27380 2360
rect 23460 980 23940 1000
rect 23460 920 23510 980
rect 23880 920 23940 980
rect 23460 850 23490 920
rect 23890 850 23940 920
rect 23460 810 23510 850
rect 23880 810 23940 850
rect 23460 740 23490 810
rect 23890 740 23940 810
rect 23460 710 23940 740
rect 25860 980 26340 1000
rect 25860 920 25910 980
rect 26280 920 26340 980
rect 25860 850 25890 920
rect 26290 850 26340 920
rect 25860 810 25910 850
rect 26280 810 26340 850
rect 25860 740 25890 810
rect 26290 740 26340 810
rect 25860 710 26340 740
rect 21800 -920 21820 -850
rect 21890 -920 21930 -850
rect 22000 -920 22060 -850
rect 21800 -960 22060 -920
rect 21800 -1030 21820 -960
rect 21890 -1030 21930 -960
rect 22000 -1030 22060 -960
rect 21800 -1070 22060 -1030
rect 21800 -1140 21820 -1070
rect 21890 -1140 21930 -1070
rect 22000 -1140 22060 -1070
rect 21800 -1180 22060 -1140
rect 21800 -1250 21820 -1180
rect 21890 -1250 21930 -1180
rect 22000 -1250 22060 -1180
rect 21800 -1290 22060 -1250
rect 21800 -1360 21820 -1290
rect 21890 -1360 21930 -1290
rect 22000 -1360 22060 -1290
rect 21800 -1400 22060 -1360
rect 21800 -1470 21820 -1400
rect 21890 -1470 21930 -1400
rect 22000 -1470 22060 -1400
rect 21800 -1510 22060 -1470
rect 21800 -1580 21820 -1510
rect 21890 -1580 21930 -1510
rect 22000 -1580 22060 -1510
rect 21800 -1620 22060 -1580
rect 21800 -1690 21820 -1620
rect 21890 -1690 21930 -1620
rect 22000 -1690 22060 -1620
rect 21800 -1730 22060 -1690
rect 21800 -1800 21820 -1730
rect 21890 -1800 21930 -1730
rect 22000 -1800 22060 -1730
rect 21800 -1840 22060 -1800
rect 21800 -1910 21820 -1840
rect 21890 -1910 21930 -1840
rect 22000 -1910 22060 -1840
rect 21800 -1950 22060 -1910
rect 21800 -2020 21820 -1950
rect 21890 -2020 21930 -1950
rect 22000 -2020 22060 -1950
rect 21800 -2040 22060 -2020
rect 24720 -3050 25050 -3030
rect 24720 -3120 24740 -3050
rect 24810 -3120 24850 -3050
rect 24920 -3120 24960 -3050
rect 25030 -3120 25050 -3050
rect 24720 -3125 25050 -3120
rect 30344 -3125 30477 3103
rect 31100 3210 37860 3300
rect 31100 2970 31180 3210
rect 31420 2970 31510 3210
rect 31750 2970 31840 3210
rect 32080 2970 32170 3210
rect 32410 2970 32500 3210
rect 32740 2970 32830 3210
rect 33070 2970 33160 3210
rect 33400 2970 33490 3210
rect 33730 2970 33820 3210
rect 34060 2970 34150 3210
rect 34390 2970 34480 3210
rect 34720 2970 34810 3210
rect 35050 2970 35140 3210
rect 35380 2970 35470 3210
rect 35710 2970 35800 3210
rect 36040 2970 36130 3210
rect 36370 2970 36460 3210
rect 36700 2970 36790 3210
rect 37030 2970 37120 3210
rect 37360 2970 37450 3210
rect 37690 2970 37860 3210
rect 31100 2880 37860 2970
rect 31100 2640 31180 2880
rect 31420 2640 31510 2880
rect 31750 2640 31840 2880
rect 32080 2640 32170 2880
rect 32410 2640 32500 2880
rect 32740 2640 32830 2880
rect 33070 2640 33160 2880
rect 33400 2640 33490 2880
rect 33730 2640 33820 2880
rect 34060 2640 34150 2880
rect 34390 2640 34480 2880
rect 34720 2640 34810 2880
rect 35050 2640 35140 2880
rect 35380 2640 35470 2880
rect 35710 2640 35800 2880
rect 36040 2640 36130 2880
rect 36370 2640 36460 2880
rect 36700 2640 36790 2880
rect 37030 2640 37120 2880
rect 37360 2640 37450 2880
rect 37690 2640 37860 2880
rect 31100 2550 37860 2640
rect 31100 2310 31180 2550
rect 31420 2310 31510 2550
rect 31750 2310 31840 2550
rect 32080 2310 32170 2550
rect 32410 2310 32500 2550
rect 32740 2310 32830 2550
rect 33070 2310 33160 2550
rect 33400 2310 33490 2550
rect 33730 2310 33820 2550
rect 34060 2310 34150 2550
rect 34390 2310 34480 2550
rect 34720 2310 34810 2550
rect 35050 2310 35140 2550
rect 35380 2310 35470 2550
rect 35710 2310 35800 2550
rect 36040 2310 36130 2550
rect 36370 2310 36460 2550
rect 36700 2310 36790 2550
rect 37030 2310 37120 2550
rect 37360 2310 37450 2550
rect 37690 2310 37860 2550
rect 31100 2220 37860 2310
rect 31100 1980 31180 2220
rect 31420 1980 31510 2220
rect 31750 1980 31840 2220
rect 32080 1980 32170 2220
rect 32410 1980 32500 2220
rect 32740 1980 32830 2220
rect 33070 1980 33160 2220
rect 33400 1980 33490 2220
rect 33730 1980 33820 2220
rect 34060 1980 34150 2220
rect 34390 1980 34480 2220
rect 34720 1980 34810 2220
rect 35050 1980 35140 2220
rect 35380 1980 35470 2220
rect 35710 1980 35800 2220
rect 36040 1980 36130 2220
rect 36370 1980 36460 2220
rect 36700 1980 36790 2220
rect 37030 1980 37120 2220
rect 37360 1980 37450 2220
rect 37690 1980 37860 2220
rect 31100 1890 37860 1980
rect 31100 1650 31180 1890
rect 31420 1650 31510 1890
rect 31750 1650 31840 1890
rect 32080 1650 32170 1890
rect 32410 1650 32500 1890
rect 32740 1650 32830 1890
rect 33070 1650 33160 1890
rect 33400 1650 33490 1890
rect 33730 1650 33820 1890
rect 34060 1650 34150 1890
rect 34390 1650 34480 1890
rect 34720 1650 34810 1890
rect 35050 1650 35140 1890
rect 35380 1650 35470 1890
rect 35710 1650 35800 1890
rect 36040 1650 36130 1890
rect 36370 1650 36460 1890
rect 36700 1650 36790 1890
rect 37030 1650 37120 1890
rect 37360 1650 37450 1890
rect 37690 1650 37860 1890
rect 31100 1560 37860 1650
rect 31100 1320 31180 1560
rect 31420 1320 31510 1560
rect 31750 1320 31840 1560
rect 32080 1320 32170 1560
rect 32410 1320 32500 1560
rect 32740 1320 32830 1560
rect 33070 1320 33160 1560
rect 33400 1320 33490 1560
rect 33730 1320 33820 1560
rect 34060 1320 34150 1560
rect 34390 1320 34480 1560
rect 34720 1320 34810 1560
rect 35050 1320 35140 1560
rect 35380 1320 35470 1560
rect 35710 1320 35800 1560
rect 36040 1320 36130 1560
rect 36370 1320 36460 1560
rect 36700 1320 36790 1560
rect 37030 1320 37120 1560
rect 37360 1320 37450 1560
rect 37690 1320 37860 1560
rect 31100 1150 37860 1320
rect 38180 7820 38500 7910
rect 38180 7750 38190 7820
rect 38260 7770 38280 7820
rect 38350 7770 38370 7820
rect 38440 7770 38500 7820
rect 38180 7730 38230 7750
rect 38180 7660 38190 7730
rect 38180 7640 38230 7660
rect 38180 7570 38190 7640
rect 38180 7550 38230 7570
rect 38180 7480 38190 7550
rect 38470 7530 38500 7770
rect 38260 7480 38280 7530
rect 38350 7480 38370 7530
rect 38440 7480 38500 7530
rect 38180 7460 38500 7480
rect 38180 7390 38190 7460
rect 38260 7440 38280 7460
rect 38350 7440 38370 7460
rect 38440 7440 38500 7460
rect 38180 7370 38230 7390
rect 38180 7300 38190 7370
rect 38180 7280 38230 7300
rect 38180 7210 38190 7280
rect 38180 7200 38230 7210
rect 38470 7200 38500 7440
rect 38180 7150 38500 7200
rect 38180 7080 38190 7150
rect 38260 7080 38280 7150
rect 38350 7080 38370 7150
rect 38440 7080 38500 7150
rect 38180 7070 38500 7080
rect 38180 7060 38230 7070
rect 38180 6990 38190 7060
rect 38180 6970 38230 6990
rect 38180 6900 38190 6970
rect 38180 6880 38230 6900
rect 38180 6810 38190 6880
rect 38470 6830 38500 7070
rect 38260 6810 38280 6830
rect 38350 6810 38370 6830
rect 38440 6810 38500 6830
rect 38180 6790 38500 6810
rect 38180 6720 38190 6790
rect 38260 6740 38280 6790
rect 38350 6740 38370 6790
rect 38440 6740 38500 6790
rect 38180 6700 38230 6720
rect 38180 6630 38190 6700
rect 38180 6610 38230 6630
rect 38180 6540 38190 6610
rect 38180 6520 38230 6540
rect 38180 6450 38190 6520
rect 38470 6500 38500 6740
rect 38260 6450 38280 6500
rect 38350 6450 38370 6500
rect 38440 6450 38500 6500
rect 38180 6430 38500 6450
rect 38180 6360 38190 6430
rect 38260 6410 38280 6430
rect 38350 6410 38370 6430
rect 38440 6410 38500 6430
rect 38180 6340 38230 6360
rect 38180 6270 38190 6340
rect 38180 6250 38230 6270
rect 38180 6180 38190 6250
rect 38180 6170 38230 6180
rect 38470 6170 38500 6410
rect 38180 6160 38500 6170
rect 38180 6090 38190 6160
rect 38260 6090 38280 6160
rect 38350 6090 38370 6160
rect 38440 6090 38500 6160
rect 38180 6080 38500 6090
rect 38180 6070 38230 6080
rect 38180 6000 38190 6070
rect 38180 5980 38230 6000
rect 38180 5910 38190 5980
rect 38180 5890 38230 5910
rect 38180 5820 38190 5890
rect 38470 5840 38500 6080
rect 38260 5820 38280 5840
rect 38350 5820 38370 5840
rect 38440 5820 38500 5840
rect 38180 5800 38500 5820
rect 38180 5730 38190 5800
rect 38260 5750 38280 5800
rect 38350 5750 38370 5800
rect 38440 5750 38500 5800
rect 38180 5710 38230 5730
rect 38180 5640 38190 5710
rect 38180 5620 38230 5640
rect 38180 5550 38190 5620
rect 38180 5530 38230 5550
rect 38180 5460 38190 5530
rect 38470 5510 38500 5750
rect 38260 5460 38280 5510
rect 38350 5460 38370 5510
rect 38440 5460 38500 5510
rect 38180 5440 38500 5460
rect 38180 5370 38190 5440
rect 38260 5420 38280 5440
rect 38350 5420 38370 5440
rect 38440 5420 38500 5440
rect 38180 5350 38230 5370
rect 38180 5280 38190 5350
rect 38180 5260 38230 5280
rect 38180 5190 38190 5260
rect 38180 5180 38230 5190
rect 38470 5180 38500 5420
rect 38180 5170 38500 5180
rect 38180 5100 38190 5170
rect 38260 5100 38280 5170
rect 38350 5100 38370 5170
rect 38440 5100 38500 5170
rect 38180 5090 38500 5100
rect 38180 5080 38230 5090
rect 38180 5010 38190 5080
rect 38180 4990 38230 5010
rect 38180 4920 38190 4990
rect 38180 4900 38230 4920
rect 38180 4830 38190 4900
rect 38470 4850 38500 5090
rect 38260 4830 38280 4850
rect 38350 4830 38370 4850
rect 38440 4830 38500 4850
rect 38180 4810 38500 4830
rect 38180 4740 38190 4810
rect 38260 4760 38280 4810
rect 38350 4760 38370 4810
rect 38440 4760 38500 4810
rect 38180 4720 38230 4740
rect 38180 4650 38190 4720
rect 38180 4630 38230 4650
rect 38180 4560 38190 4630
rect 38180 4540 38230 4560
rect 38180 4470 38190 4540
rect 38470 4520 38500 4760
rect 38260 4470 38280 4520
rect 38350 4470 38370 4520
rect 38440 4470 38500 4520
rect 38180 4450 38500 4470
rect 38180 4380 38190 4450
rect 38260 4430 38280 4450
rect 38350 4430 38370 4450
rect 38440 4430 38500 4450
rect 38180 4360 38230 4380
rect 38180 4290 38190 4360
rect 38180 4270 38230 4290
rect 38180 4200 38190 4270
rect 38180 4190 38230 4200
rect 38470 4190 38500 4430
rect 38180 4140 38500 4190
rect 38180 4070 38190 4140
rect 38260 4070 38280 4140
rect 38350 4070 38370 4140
rect 38440 4070 38500 4140
rect 38180 4060 38500 4070
rect 38180 4050 38230 4060
rect 38180 3980 38190 4050
rect 38180 3960 38230 3980
rect 38180 3890 38190 3960
rect 38180 3870 38230 3890
rect 38180 3800 38190 3870
rect 38470 3820 38500 4060
rect 38260 3800 38280 3820
rect 38350 3800 38370 3820
rect 38440 3800 38500 3820
rect 38180 3780 38500 3800
rect 38180 3710 38190 3780
rect 38260 3730 38280 3780
rect 38350 3730 38370 3780
rect 38440 3730 38500 3780
rect 38180 3690 38230 3710
rect 38180 3620 38190 3690
rect 38180 3600 38230 3620
rect 38180 3530 38190 3600
rect 38180 3510 38230 3530
rect 38180 3440 38190 3510
rect 38470 3490 38500 3730
rect 38260 3440 38280 3490
rect 38350 3440 38370 3490
rect 38440 3440 38500 3490
rect 38180 3420 38500 3440
rect 38180 3350 38190 3420
rect 38260 3400 38280 3420
rect 38350 3400 38370 3420
rect 38440 3400 38500 3420
rect 38180 3330 38230 3350
rect 38180 3260 38190 3330
rect 38180 3240 38230 3260
rect 38180 3170 38190 3240
rect 38180 3160 38230 3170
rect 38470 3160 38500 3400
rect 38180 3150 38500 3160
rect 38180 3080 38190 3150
rect 38260 3080 38280 3150
rect 38350 3080 38370 3150
rect 38440 3080 38500 3150
rect 38180 3070 38500 3080
rect 38180 3060 38230 3070
rect 38180 2990 38190 3060
rect 38180 2970 38230 2990
rect 38180 2900 38190 2970
rect 38180 2880 38230 2900
rect 38180 2810 38190 2880
rect 38470 2830 38500 3070
rect 38260 2810 38280 2830
rect 38350 2810 38370 2830
rect 38440 2810 38500 2830
rect 38180 2790 38500 2810
rect 38180 2720 38190 2790
rect 38260 2740 38280 2790
rect 38350 2740 38370 2790
rect 38440 2740 38500 2790
rect 38180 2700 38230 2720
rect 38180 2630 38190 2700
rect 38180 2610 38230 2630
rect 38180 2540 38190 2610
rect 38180 2520 38230 2540
rect 38180 2450 38190 2520
rect 38470 2500 38500 2740
rect 38260 2450 38280 2500
rect 38350 2450 38370 2500
rect 38440 2450 38500 2500
rect 38180 2430 38500 2450
rect 38180 2360 38190 2430
rect 38260 2410 38280 2430
rect 38350 2410 38370 2430
rect 38440 2410 38500 2430
rect 38180 2340 38230 2360
rect 38180 2270 38190 2340
rect 38180 2250 38230 2270
rect 38180 2180 38190 2250
rect 38180 2170 38230 2180
rect 38470 2170 38500 2410
rect 38180 2160 38500 2170
rect 38180 2090 38190 2160
rect 38260 2090 38280 2160
rect 38350 2090 38370 2160
rect 38440 2090 38500 2160
rect 38180 2080 38500 2090
rect 38180 2070 38230 2080
rect 38180 2000 38190 2070
rect 38180 1980 38230 2000
rect 38180 1910 38190 1980
rect 38180 1890 38230 1910
rect 38180 1820 38190 1890
rect 38470 1840 38500 2080
rect 38260 1820 38280 1840
rect 38350 1820 38370 1840
rect 38440 1820 38500 1840
rect 38180 1800 38500 1820
rect 38180 1730 38190 1800
rect 38260 1750 38280 1800
rect 38350 1750 38370 1800
rect 38440 1750 38500 1800
rect 38180 1710 38230 1730
rect 38180 1640 38190 1710
rect 38180 1620 38230 1640
rect 38180 1550 38190 1620
rect 38180 1530 38230 1550
rect 38180 1460 38190 1530
rect 38470 1510 38500 1750
rect 38260 1460 38280 1510
rect 38350 1460 38370 1510
rect 38440 1460 38500 1510
rect 38180 1440 38500 1460
rect 38180 1370 38190 1440
rect 38260 1420 38280 1440
rect 38350 1420 38370 1440
rect 38440 1420 38500 1440
rect 38180 1350 38230 1370
rect 38180 1280 38190 1350
rect 38180 1260 38230 1280
rect 38180 1190 38190 1260
rect 38180 1180 38230 1190
rect 38470 1180 38500 1420
rect 38180 1150 38500 1180
rect 31100 230 37860 310
rect 31100 20 31180 230
rect 30720 0 31180 20
rect 30720 -70 30740 0
rect 30810 -70 30850 0
rect 30920 -10 31180 0
rect 31420 -10 31510 230
rect 31750 -10 31840 230
rect 32080 -10 32170 230
rect 32410 -10 32500 230
rect 32740 -10 32830 230
rect 33070 -10 33160 230
rect 33400 -10 33490 230
rect 33730 -10 33820 230
rect 34060 -10 34150 230
rect 34390 -10 34480 230
rect 34720 -10 34810 230
rect 35050 -10 35140 230
rect 35380 -10 35470 230
rect 35710 -10 35800 230
rect 36040 -10 36130 230
rect 36370 -10 36460 230
rect 36700 -10 36790 230
rect 37030 -10 37120 230
rect 37360 -10 37450 230
rect 37690 -10 37860 230
rect 30920 -70 37860 -10
rect 30720 -100 37860 -70
rect 30720 -130 31180 -100
rect 30720 -200 30740 -130
rect 30810 -200 30850 -130
rect 30920 -200 31180 -130
rect 30720 -260 31180 -200
rect 30720 -330 30740 -260
rect 30810 -330 30850 -260
rect 30920 -330 31180 -260
rect 30720 -340 31180 -330
rect 31420 -340 31510 -100
rect 31750 -340 31840 -100
rect 32080 -340 32170 -100
rect 32410 -340 32500 -100
rect 32740 -340 32830 -100
rect 33070 -340 33160 -100
rect 33400 -340 33490 -100
rect 33730 -340 33820 -100
rect 34060 -340 34150 -100
rect 34390 -340 34480 -100
rect 34720 -340 34810 -100
rect 35050 -340 35140 -100
rect 35380 -340 35470 -100
rect 35710 -340 35800 -100
rect 36040 -340 36130 -100
rect 36370 -340 36460 -100
rect 36700 -340 36790 -100
rect 37030 -340 37120 -100
rect 37360 -340 37450 -100
rect 37690 -340 37860 -100
rect 30720 -350 37860 -340
rect 24720 -3160 30477 -3125
rect 24720 -3230 24740 -3160
rect 24810 -3230 24850 -3160
rect 24920 -3230 24960 -3160
rect 25030 -3230 30477 -3160
rect 24720 -3258 30477 -3230
rect 24720 -3270 25050 -3258
rect 24720 -3340 24740 -3270
rect 24810 -3340 24850 -3270
rect 24920 -3340 24960 -3270
rect 25030 -3340 25050 -3270
rect 24720 -3360 25050 -3340
rect 22420 -3690 22900 -3660
rect 22420 -3760 22470 -3690
rect 22870 -3760 22900 -3690
rect 22420 -3800 22480 -3760
rect 22850 -3800 22900 -3760
rect 22420 -3870 22470 -3800
rect 22870 -3870 22900 -3800
rect 22420 -3930 22480 -3870
rect 22850 -3930 22900 -3870
rect 22420 -3950 22900 -3930
rect 26900 -3690 27380 -3660
rect 26900 -3760 26950 -3690
rect 27350 -3760 27380 -3690
rect 26900 -3800 26960 -3760
rect 27330 -3800 27380 -3760
rect 26900 -3870 26950 -3800
rect 27350 -3870 27380 -3800
rect 26900 -3930 26960 -3870
rect 27330 -3930 27380 -3870
rect 26900 -3950 27380 -3930
rect 26400 -5890 26880 -5780
rect 26400 -5915 26510 -5890
rect 18975 -6025 26510 -5915
rect -1200 -6330 90 -6320
rect -1200 -6370 -1160 -6330
rect -1090 -6370 -1070 -6330
rect -1000 -6370 -980 -6330
rect -1200 -6610 -1170 -6370
rect -910 -6400 -890 -6330
rect -820 -6370 -800 -6330
rect -730 -6370 -710 -6330
rect -640 -6370 -620 -6330
rect -550 -6400 -530 -6330
rect -460 -6370 -440 -6330
rect -370 -6370 -350 -6330
rect -280 -6370 -260 -6330
rect -270 -6400 -260 -6370
rect -190 -6370 -170 -6330
rect -100 -6370 -80 -6330
rect -10 -6370 10 -6330
rect -190 -6400 -180 -6370
rect 80 -6400 90 -6330
rect -930 -6420 -840 -6400
rect -600 -6420 -510 -6400
rect -270 -6420 -180 -6400
rect 60 -6420 90 -6400
rect -910 -6490 -890 -6420
rect -550 -6490 -530 -6420
rect -270 -6490 -260 -6420
rect -190 -6490 -180 -6420
rect 80 -6490 90 -6420
rect -930 -6510 -840 -6490
rect -600 -6510 -510 -6490
rect -270 -6510 -180 -6490
rect 60 -6510 90 -6490
rect -910 -6580 -890 -6510
rect -550 -6580 -530 -6510
rect -270 -6580 -260 -6510
rect -190 -6580 -180 -6510
rect 80 -6580 90 -6510
rect -930 -6610 -840 -6580
rect -600 -6610 -510 -6580
rect -270 -6610 -180 -6580
rect 60 -6610 90 -6580
rect -1200 -6640 90 -6610
rect 14690 -6330 15980 -6320
rect 14690 -6400 14700 -6330
rect 14770 -6370 14790 -6330
rect 14860 -6370 14880 -6330
rect 14950 -6370 14970 -6330
rect 14960 -6400 14970 -6370
rect 15040 -6370 15060 -6330
rect 15130 -6370 15150 -6330
rect 15220 -6370 15240 -6330
rect 15040 -6400 15050 -6370
rect 15310 -6400 15330 -6330
rect 15400 -6370 15420 -6330
rect 15490 -6370 15510 -6330
rect 15580 -6370 15600 -6330
rect 15670 -6400 15690 -6330
rect 15760 -6370 15780 -6330
rect 15850 -6370 15870 -6330
rect 15940 -6370 15980 -6330
rect 14690 -6420 14720 -6400
rect 14960 -6420 15050 -6400
rect 15290 -6420 15380 -6400
rect 15620 -6420 15710 -6400
rect 14690 -6490 14700 -6420
rect 14960 -6490 14970 -6420
rect 15040 -6490 15050 -6420
rect 15310 -6490 15330 -6420
rect 15670 -6490 15690 -6420
rect 14690 -6510 14720 -6490
rect 14960 -6510 15050 -6490
rect 15290 -6510 15380 -6490
rect 15620 -6510 15710 -6490
rect 14690 -6580 14700 -6510
rect 14960 -6580 14970 -6510
rect 15040 -6580 15050 -6510
rect 15310 -6580 15330 -6510
rect 15670 -6580 15690 -6510
rect 14690 -6610 14720 -6580
rect 14960 -6610 15050 -6580
rect 15290 -6610 15380 -6580
rect 15620 -6610 15710 -6580
rect 15950 -6610 15980 -6370
rect 14690 -6640 15980 -6610
rect 0 -8140 310 -8120
rect 0 -8210 20 -8140
rect 90 -8210 130 -8140
rect 200 -8210 230 -8140
rect 300 -8210 310 -8140
rect 0 -8235 310 -8210
rect -2710 -8250 310 -8235
rect -2710 -8320 20 -8250
rect 90 -8320 130 -8250
rect 200 -8320 230 -8250
rect 300 -8320 310 -8250
rect -2710 -8345 310 -8320
rect 0 -8360 310 -8345
rect 0 -8430 20 -8360
rect 90 -8430 130 -8360
rect 200 -8430 230 -8360
rect 300 -8430 310 -8360
rect 0 -8450 310 -8430
rect 14590 -8230 14900 -8210
rect 14590 -8300 14600 -8230
rect 14670 -8300 14700 -8230
rect 14770 -8300 14810 -8230
rect 14880 -8300 14900 -8230
rect 14590 -8325 14900 -8300
rect 18975 -8325 19085 -6025
rect 14590 -8340 19085 -8325
rect 14590 -8410 14600 -8340
rect 14670 -8410 14700 -8340
rect 14770 -8410 14810 -8340
rect 14880 -8410 19085 -8340
rect 14590 -8435 19085 -8410
rect 21610 -8360 21930 -8330
rect 21610 -8430 21630 -8360
rect 21700 -8370 21730 -8360
rect 21800 -8370 21830 -8360
rect 21900 -8430 21930 -8360
rect 14590 -8450 14900 -8435
rect 14590 -8520 14600 -8450
rect 14670 -8520 14700 -8450
rect 14770 -8520 14810 -8450
rect 14880 -8520 14900 -8450
rect 14590 -8540 14900 -8520
rect 21610 -8460 21650 -8430
rect 21890 -8460 21930 -8430
rect 21610 -8530 21630 -8460
rect 21900 -8530 21930 -8460
rect 21610 -8560 21650 -8530
rect 21890 -8560 21930 -8530
rect 21610 -8630 21630 -8560
rect 21700 -8630 21730 -8610
rect 21800 -8630 21830 -8610
rect 21900 -8630 21930 -8560
rect 21610 -8650 21930 -8630
rect 22630 -9010 22950 -8980
rect 22630 -9080 22650 -9010
rect 22720 -9080 22750 -9010
rect 22820 -9080 22850 -9010
rect 22920 -9080 22950 -9010
rect 22630 -9110 22950 -9080
rect 22630 -9180 22650 -9110
rect 22720 -9180 22750 -9110
rect 22820 -9180 22850 -9110
rect 22920 -9180 22950 -9110
rect 22630 -9210 22950 -9180
rect 22630 -9280 22650 -9210
rect 22720 -9280 22750 -9210
rect 22820 -9280 22850 -9210
rect 22920 -9280 22950 -9210
rect 1080 -10340 2680 -10310
rect 1080 -10410 1150 -10340
rect 1220 -10410 1260 -10340
rect 1550 -10410 1590 -10340
rect 1880 -10410 1920 -10340
rect 2210 -10410 2250 -10340
rect 2540 -10410 2580 -10340
rect 2650 -10410 2680 -10340
rect 1080 -10450 1260 -10410
rect 1500 -10450 1590 -10410
rect 1830 -10450 1930 -10410
rect 2170 -10450 2260 -10410
rect 2500 -10450 2680 -10410
rect 1080 -10520 1150 -10450
rect 1220 -10520 1260 -10450
rect 1550 -10520 1590 -10450
rect 1880 -10520 1920 -10450
rect 2210 -10520 2250 -10450
rect 2540 -10520 2580 -10450
rect 2650 -10520 2680 -10450
rect 1080 -10580 1260 -10520
rect 1500 -10580 1590 -10520
rect 1830 -10580 1930 -10520
rect 2170 -10580 2260 -10520
rect 2500 -10580 2680 -10520
rect 1080 -10600 2680 -10580
rect 12220 -10370 13820 -10340
rect 12220 -10440 12290 -10370
rect 12360 -10440 12400 -10370
rect 12690 -10440 12730 -10370
rect 13020 -10440 13060 -10370
rect 13350 -10440 13390 -10370
rect 13680 -10440 13720 -10370
rect 13790 -10440 13820 -10370
rect 12220 -10480 12400 -10440
rect 12640 -10480 12730 -10440
rect 12970 -10480 13070 -10440
rect 13310 -10480 13400 -10440
rect 13640 -10480 13820 -10440
rect 12220 -10550 12290 -10480
rect 12360 -10550 12400 -10480
rect 12690 -10550 12730 -10480
rect 13020 -10550 13060 -10480
rect 13350 -10550 13390 -10480
rect 13680 -10550 13720 -10480
rect 13790 -10550 13820 -10480
rect 12220 -10610 12400 -10550
rect 12640 -10610 12730 -10550
rect 12970 -10610 13070 -10550
rect 13310 -10610 13400 -10550
rect 13640 -10610 13820 -10550
rect 12220 -10620 13820 -10610
rect 22630 -10510 22950 -9280
rect 22630 -10520 30080 -10510
rect 22630 -10590 29990 -10520
rect 30060 -10590 30080 -10520
rect 22630 -10630 30080 -10590
rect 22630 -10700 29990 -10630
rect 30060 -10700 30080 -10630
rect 22630 -10740 30080 -10700
rect 22630 -10810 29990 -10740
rect 30060 -10810 30080 -10740
rect 22630 -10830 30080 -10810
rect 30344 -10995 30477 -3258
rect 31100 -430 37860 -350
rect 31100 -670 31180 -430
rect 31420 -670 31510 -430
rect 31750 -670 31840 -430
rect 32080 -670 32170 -430
rect 32410 -670 32500 -430
rect 32740 -670 32830 -430
rect 33070 -670 33160 -430
rect 33400 -670 33490 -430
rect 33730 -670 33820 -430
rect 34060 -670 34150 -430
rect 34390 -670 34480 -430
rect 34720 -670 34810 -430
rect 35050 -670 35140 -430
rect 35380 -670 35470 -430
rect 35710 -670 35800 -430
rect 36040 -670 36130 -430
rect 36370 -670 36460 -430
rect 36700 -670 36790 -430
rect 37030 -670 37120 -430
rect 37360 -670 37450 -430
rect 37690 -670 37860 -430
rect 31100 -760 37860 -670
rect 31100 -1000 31180 -760
rect 31420 -1000 31510 -760
rect 31750 -1000 31840 -760
rect 32080 -1000 32170 -760
rect 32410 -1000 32500 -760
rect 32740 -1000 32830 -760
rect 33070 -1000 33160 -760
rect 33400 -1000 33490 -760
rect 33730 -1000 33820 -760
rect 34060 -1000 34150 -760
rect 34390 -1000 34480 -760
rect 34720 -1000 34810 -760
rect 35050 -1000 35140 -760
rect 35380 -1000 35470 -760
rect 35710 -1000 35800 -760
rect 36040 -1000 36130 -760
rect 36370 -1000 36460 -760
rect 36700 -1000 36790 -760
rect 37030 -1000 37120 -760
rect 37360 -1000 37450 -760
rect 37690 -1000 37860 -760
rect 31100 -1090 37860 -1000
rect 31100 -1330 31180 -1090
rect 31420 -1330 31510 -1090
rect 31750 -1330 31840 -1090
rect 32080 -1330 32170 -1090
rect 32410 -1330 32500 -1090
rect 32740 -1330 32830 -1090
rect 33070 -1330 33160 -1090
rect 33400 -1330 33490 -1090
rect 33730 -1330 33820 -1090
rect 34060 -1330 34150 -1090
rect 34390 -1330 34480 -1090
rect 34720 -1330 34810 -1090
rect 35050 -1330 35140 -1090
rect 35380 -1330 35470 -1090
rect 35710 -1330 35800 -1090
rect 36040 -1330 36130 -1090
rect 36370 -1330 36460 -1090
rect 36700 -1330 36790 -1090
rect 37030 -1330 37120 -1090
rect 37360 -1330 37450 -1090
rect 37690 -1330 37860 -1090
rect 31100 -1420 37860 -1330
rect 31100 -1660 31180 -1420
rect 31420 -1660 31510 -1420
rect 31750 -1660 31840 -1420
rect 32080 -1660 32170 -1420
rect 32410 -1660 32500 -1420
rect 32740 -1660 32830 -1420
rect 33070 -1660 33160 -1420
rect 33400 -1660 33490 -1420
rect 33730 -1660 33820 -1420
rect 34060 -1660 34150 -1420
rect 34390 -1660 34480 -1420
rect 34720 -1660 34810 -1420
rect 35050 -1660 35140 -1420
rect 35380 -1660 35470 -1420
rect 35710 -1660 35800 -1420
rect 36040 -1660 36130 -1420
rect 36370 -1660 36460 -1420
rect 36700 -1660 36790 -1420
rect 37030 -1660 37120 -1420
rect 37360 -1660 37450 -1420
rect 37690 -1660 37860 -1420
rect 31100 -1750 37860 -1660
rect 31100 -1990 31180 -1750
rect 31420 -1990 31510 -1750
rect 31750 -1990 31840 -1750
rect 32080 -1990 32170 -1750
rect 32410 -1990 32500 -1750
rect 32740 -1990 32830 -1750
rect 33070 -1990 33160 -1750
rect 33400 -1990 33490 -1750
rect 33730 -1990 33820 -1750
rect 34060 -1990 34150 -1750
rect 34390 -1990 34480 -1750
rect 34720 -1990 34810 -1750
rect 35050 -1990 35140 -1750
rect 35380 -1990 35470 -1750
rect 35710 -1990 35800 -1750
rect 36040 -1990 36130 -1750
rect 36370 -1990 36460 -1750
rect 36700 -1990 36790 -1750
rect 37030 -1990 37120 -1750
rect 37360 -1990 37450 -1750
rect 37690 -1990 37860 -1750
rect 31100 -2080 37860 -1990
rect 31100 -2320 31180 -2080
rect 31420 -2320 31510 -2080
rect 31750 -2320 31840 -2080
rect 32080 -2320 32170 -2080
rect 32410 -2320 32500 -2080
rect 32740 -2320 32830 -2080
rect 33070 -2320 33160 -2080
rect 33400 -2320 33490 -2080
rect 33730 -2320 33820 -2080
rect 34060 -2320 34150 -2080
rect 34390 -2320 34480 -2080
rect 34720 -2320 34810 -2080
rect 35050 -2320 35140 -2080
rect 35380 -2320 35470 -2080
rect 35710 -2320 35800 -2080
rect 36040 -2320 36130 -2080
rect 36370 -2320 36460 -2080
rect 36700 -2320 36790 -2080
rect 37030 -2320 37120 -2080
rect 37360 -2320 37450 -2080
rect 37690 -2320 37860 -2080
rect 31100 -2410 37860 -2320
rect 31100 -2650 31180 -2410
rect 31420 -2650 31510 -2410
rect 31750 -2650 31840 -2410
rect 32080 -2650 32170 -2410
rect 32410 -2650 32500 -2410
rect 32740 -2650 32830 -2410
rect 33070 -2650 33160 -2410
rect 33400 -2650 33490 -2410
rect 33730 -2650 33820 -2410
rect 34060 -2650 34150 -2410
rect 34390 -2650 34480 -2410
rect 34720 -2650 34810 -2410
rect 35050 -2650 35140 -2410
rect 35380 -2650 35470 -2410
rect 35710 -2650 35800 -2410
rect 36040 -2650 36130 -2410
rect 36370 -2650 36460 -2410
rect 36700 -2650 36790 -2410
rect 37030 -2650 37120 -2410
rect 37360 -2650 37450 -2410
rect 37690 -2650 37860 -2410
rect 31100 -2740 37860 -2650
rect 31100 -2980 31180 -2740
rect 31420 -2980 31510 -2740
rect 31750 -2980 31840 -2740
rect 32080 -2980 32170 -2740
rect 32410 -2980 32500 -2740
rect 32740 -2980 32830 -2740
rect 33070 -2980 33160 -2740
rect 33400 -2980 33490 -2740
rect 33730 -2980 33820 -2740
rect 34060 -2980 34150 -2740
rect 34390 -2980 34480 -2740
rect 34720 -2980 34810 -2740
rect 35050 -2980 35140 -2740
rect 35380 -2980 35470 -2740
rect 35710 -2980 35800 -2740
rect 36040 -2980 36130 -2740
rect 36370 -2980 36460 -2740
rect 36700 -2980 36790 -2740
rect 37030 -2980 37120 -2740
rect 37360 -2980 37450 -2740
rect 37690 -2980 37860 -2740
rect 31100 -3070 37860 -2980
rect 31100 -3310 31180 -3070
rect 31420 -3310 31510 -3070
rect 31750 -3310 31840 -3070
rect 32080 -3310 32170 -3070
rect 32410 -3310 32500 -3070
rect 32740 -3310 32830 -3070
rect 33070 -3310 33160 -3070
rect 33400 -3310 33490 -3070
rect 33730 -3310 33820 -3070
rect 34060 -3310 34150 -3070
rect 34390 -3310 34480 -3070
rect 34720 -3310 34810 -3070
rect 35050 -3310 35140 -3070
rect 35380 -3310 35470 -3070
rect 35710 -3310 35800 -3070
rect 36040 -3310 36130 -3070
rect 36370 -3310 36460 -3070
rect 36700 -3310 36790 -3070
rect 37030 -3310 37120 -3070
rect 37360 -3310 37450 -3070
rect 37690 -3310 37860 -3070
rect 31100 -3400 37860 -3310
rect 31100 -3640 31180 -3400
rect 31420 -3640 31510 -3400
rect 31750 -3640 31840 -3400
rect 32080 -3640 32170 -3400
rect 32410 -3640 32500 -3400
rect 32740 -3640 32830 -3400
rect 33070 -3640 33160 -3400
rect 33400 -3640 33490 -3400
rect 33730 -3640 33820 -3400
rect 34060 -3640 34150 -3400
rect 34390 -3640 34480 -3400
rect 34720 -3640 34810 -3400
rect 35050 -3640 35140 -3400
rect 35380 -3640 35470 -3400
rect 35710 -3640 35800 -3400
rect 36040 -3640 36130 -3400
rect 36370 -3640 36460 -3400
rect 36700 -3640 36790 -3400
rect 37030 -3640 37120 -3400
rect 37360 -3640 37450 -3400
rect 37690 -3640 37860 -3400
rect 31100 -3730 37860 -3640
rect 31100 -3970 31180 -3730
rect 31420 -3970 31510 -3730
rect 31750 -3970 31840 -3730
rect 32080 -3970 32170 -3730
rect 32410 -3970 32500 -3730
rect 32740 -3970 32830 -3730
rect 33070 -3970 33160 -3730
rect 33400 -3970 33490 -3730
rect 33730 -3970 33820 -3730
rect 34060 -3970 34150 -3730
rect 34390 -3970 34480 -3730
rect 34720 -3970 34810 -3730
rect 35050 -3970 35140 -3730
rect 35380 -3970 35470 -3730
rect 35710 -3970 35800 -3730
rect 36040 -3970 36130 -3730
rect 36370 -3970 36460 -3730
rect 36700 -3970 36790 -3730
rect 37030 -3970 37120 -3730
rect 37360 -3970 37450 -3730
rect 37690 -3970 37860 -3730
rect 31100 -4060 37860 -3970
rect 31100 -4300 31180 -4060
rect 31420 -4300 31510 -4060
rect 31750 -4300 31840 -4060
rect 32080 -4300 32170 -4060
rect 32410 -4300 32500 -4060
rect 32740 -4300 32830 -4060
rect 33070 -4300 33160 -4060
rect 33400 -4300 33490 -4060
rect 33730 -4300 33820 -4060
rect 34060 -4300 34150 -4060
rect 34390 -4300 34480 -4060
rect 34720 -4300 34810 -4060
rect 35050 -4300 35140 -4060
rect 35380 -4300 35470 -4060
rect 35710 -4300 35800 -4060
rect 36040 -4300 36130 -4060
rect 36370 -4300 36460 -4060
rect 36700 -4300 36790 -4060
rect 37030 -4300 37120 -4060
rect 37360 -4300 37450 -4060
rect 37690 -4300 37860 -4060
rect 31100 -4390 37860 -4300
rect 31100 -4630 31180 -4390
rect 31420 -4630 31510 -4390
rect 31750 -4630 31840 -4390
rect 32080 -4630 32170 -4390
rect 32410 -4630 32500 -4390
rect 32740 -4630 32830 -4390
rect 33070 -4630 33160 -4390
rect 33400 -4630 33490 -4390
rect 33730 -4630 33820 -4390
rect 34060 -4630 34150 -4390
rect 34390 -4630 34480 -4390
rect 34720 -4630 34810 -4390
rect 35050 -4630 35140 -4390
rect 35380 -4630 35470 -4390
rect 35710 -4630 35800 -4390
rect 36040 -4630 36130 -4390
rect 36370 -4630 36460 -4390
rect 36700 -4630 36790 -4390
rect 37030 -4630 37120 -4390
rect 37360 -4630 37450 -4390
rect 37690 -4630 37860 -4390
rect 31100 -4720 37860 -4630
rect 31100 -4960 31180 -4720
rect 31420 -4960 31510 -4720
rect 31750 -4960 31840 -4720
rect 32080 -4960 32170 -4720
rect 32410 -4960 32500 -4720
rect 32740 -4960 32830 -4720
rect 33070 -4960 33160 -4720
rect 33400 -4960 33490 -4720
rect 33730 -4960 33820 -4720
rect 34060 -4960 34150 -4720
rect 34390 -4960 34480 -4720
rect 34720 -4960 34810 -4720
rect 35050 -4960 35140 -4720
rect 35380 -4960 35470 -4720
rect 35710 -4960 35800 -4720
rect 36040 -4960 36130 -4720
rect 36370 -4960 36460 -4720
rect 36700 -4960 36790 -4720
rect 37030 -4960 37120 -4720
rect 37360 -4960 37450 -4720
rect 37690 -4960 37860 -4720
rect 31100 -5050 37860 -4960
rect 31100 -5290 31180 -5050
rect 31420 -5290 31510 -5050
rect 31750 -5290 31840 -5050
rect 32080 -5290 32170 -5050
rect 32410 -5290 32500 -5050
rect 32740 -5290 32830 -5050
rect 33070 -5290 33160 -5050
rect 33400 -5290 33490 -5050
rect 33730 -5290 33820 -5050
rect 34060 -5290 34150 -5050
rect 34390 -5290 34480 -5050
rect 34720 -5290 34810 -5050
rect 35050 -5290 35140 -5050
rect 35380 -5290 35470 -5050
rect 35710 -5290 35800 -5050
rect 36040 -5290 36130 -5050
rect 36370 -5290 36460 -5050
rect 36700 -5290 36790 -5050
rect 37030 -5290 37120 -5050
rect 37360 -5290 37450 -5050
rect 37690 -5290 37860 -5050
rect 31100 -5380 37860 -5290
rect 31100 -5620 31180 -5380
rect 31420 -5620 31510 -5380
rect 31750 -5620 31840 -5380
rect 32080 -5620 32170 -5380
rect 32410 -5620 32500 -5380
rect 32740 -5620 32830 -5380
rect 33070 -5620 33160 -5380
rect 33400 -5620 33490 -5380
rect 33730 -5620 33820 -5380
rect 34060 -5620 34150 -5380
rect 34390 -5620 34480 -5380
rect 34720 -5620 34810 -5380
rect 35050 -5620 35140 -5380
rect 35380 -5620 35470 -5380
rect 35710 -5620 35800 -5380
rect 36040 -5620 36130 -5380
rect 36370 -5620 36460 -5380
rect 36700 -5620 36790 -5380
rect 37030 -5620 37120 -5380
rect 37360 -5620 37450 -5380
rect 37690 -5620 37860 -5380
rect 31100 -5710 37860 -5620
rect 31100 -5950 31180 -5710
rect 31420 -5950 31510 -5710
rect 31750 -5950 31840 -5710
rect 32080 -5950 32170 -5710
rect 32410 -5950 32500 -5710
rect 32740 -5950 32830 -5710
rect 33070 -5950 33160 -5710
rect 33400 -5950 33490 -5710
rect 33730 -5950 33820 -5710
rect 34060 -5950 34150 -5710
rect 34390 -5950 34480 -5710
rect 34720 -5950 34810 -5710
rect 35050 -5950 35140 -5710
rect 35380 -5950 35470 -5710
rect 35710 -5950 35800 -5710
rect 36040 -5950 36130 -5710
rect 36370 -5950 36460 -5710
rect 36700 -5950 36790 -5710
rect 37030 -5950 37120 -5710
rect 37360 -5950 37450 -5710
rect 37690 -5950 37860 -5710
rect 31100 -6040 37860 -5950
rect 31100 -6280 31180 -6040
rect 31420 -6280 31510 -6040
rect 31750 -6280 31840 -6040
rect 32080 -6280 32170 -6040
rect 32410 -6280 32500 -6040
rect 32740 -6280 32830 -6040
rect 33070 -6280 33160 -6040
rect 33400 -6280 33490 -6040
rect 33730 -6280 33820 -6040
rect 34060 -6280 34150 -6040
rect 34390 -6280 34480 -6040
rect 34720 -6280 34810 -6040
rect 35050 -6280 35140 -6040
rect 35380 -6280 35470 -6040
rect 35710 -6280 35800 -6040
rect 36040 -6280 36130 -6040
rect 36370 -6280 36460 -6040
rect 36700 -6280 36790 -6040
rect 37030 -6280 37120 -6040
rect 37360 -6280 37450 -6040
rect 37690 -6280 37860 -6040
rect 31100 -6450 37860 -6280
rect 38180 220 38500 310
rect 38180 150 38190 220
rect 38260 170 38280 220
rect 38350 170 38370 220
rect 38440 170 38500 220
rect 38180 130 38230 150
rect 38180 60 38190 130
rect 38180 40 38230 60
rect 38180 -30 38190 40
rect 38180 -50 38230 -30
rect 38180 -120 38190 -50
rect 38470 -70 38500 170
rect 38260 -120 38280 -70
rect 38350 -120 38370 -70
rect 38440 -120 38500 -70
rect 38180 -140 38500 -120
rect 38180 -210 38190 -140
rect 38260 -160 38280 -140
rect 38350 -160 38370 -140
rect 38440 -160 38500 -140
rect 38180 -230 38230 -210
rect 38180 -300 38190 -230
rect 38180 -320 38230 -300
rect 38180 -390 38190 -320
rect 38180 -400 38230 -390
rect 38470 -400 38500 -160
rect 38180 -450 38500 -400
rect 38180 -520 38190 -450
rect 38260 -520 38280 -450
rect 38350 -520 38370 -450
rect 38440 -520 38500 -450
rect 38180 -530 38500 -520
rect 38180 -540 38230 -530
rect 38180 -610 38190 -540
rect 38180 -630 38230 -610
rect 38180 -700 38190 -630
rect 38180 -720 38230 -700
rect 38180 -790 38190 -720
rect 38470 -770 38500 -530
rect 38260 -790 38280 -770
rect 38350 -790 38370 -770
rect 38440 -790 38500 -770
rect 38180 -810 38500 -790
rect 38180 -880 38190 -810
rect 38260 -860 38280 -810
rect 38350 -860 38370 -810
rect 38440 -860 38500 -810
rect 38180 -900 38230 -880
rect 38180 -970 38190 -900
rect 38180 -990 38230 -970
rect 38180 -1060 38190 -990
rect 38180 -1080 38230 -1060
rect 38180 -1150 38190 -1080
rect 38470 -1100 38500 -860
rect 38260 -1150 38280 -1100
rect 38350 -1150 38370 -1100
rect 38440 -1150 38500 -1100
rect 38180 -1170 38500 -1150
rect 38180 -1240 38190 -1170
rect 38260 -1190 38280 -1170
rect 38350 -1190 38370 -1170
rect 38440 -1190 38500 -1170
rect 38180 -1260 38230 -1240
rect 38180 -1330 38190 -1260
rect 38180 -1350 38230 -1330
rect 38180 -1420 38190 -1350
rect 38180 -1430 38230 -1420
rect 38470 -1430 38500 -1190
rect 38180 -1440 38500 -1430
rect 38180 -1510 38190 -1440
rect 38260 -1510 38280 -1440
rect 38350 -1510 38370 -1440
rect 38440 -1510 38500 -1440
rect 38180 -1520 38500 -1510
rect 38180 -1530 38230 -1520
rect 38180 -1600 38190 -1530
rect 38180 -1620 38230 -1600
rect 38180 -1690 38190 -1620
rect 38180 -1710 38230 -1690
rect 38180 -1780 38190 -1710
rect 38470 -1760 38500 -1520
rect 38260 -1780 38280 -1760
rect 38350 -1780 38370 -1760
rect 38440 -1780 38500 -1760
rect 38180 -1800 38500 -1780
rect 38180 -1870 38190 -1800
rect 38260 -1850 38280 -1800
rect 38350 -1850 38370 -1800
rect 38440 -1850 38500 -1800
rect 38180 -1890 38230 -1870
rect 38180 -1960 38190 -1890
rect 38180 -1980 38230 -1960
rect 38180 -2050 38190 -1980
rect 38180 -2070 38230 -2050
rect 38180 -2140 38190 -2070
rect 38470 -2090 38500 -1850
rect 38260 -2140 38280 -2090
rect 38350 -2140 38370 -2090
rect 38440 -2140 38500 -2090
rect 38180 -2160 38500 -2140
rect 38180 -2230 38190 -2160
rect 38260 -2180 38280 -2160
rect 38350 -2180 38370 -2160
rect 38440 -2180 38500 -2160
rect 38180 -2250 38230 -2230
rect 38180 -2320 38190 -2250
rect 38180 -2340 38230 -2320
rect 38180 -2410 38190 -2340
rect 38180 -2420 38230 -2410
rect 38470 -2420 38500 -2180
rect 38180 -2430 38500 -2420
rect 38180 -2500 38190 -2430
rect 38260 -2500 38280 -2430
rect 38350 -2500 38370 -2430
rect 38440 -2500 38500 -2430
rect 38180 -2510 38500 -2500
rect 38180 -2520 38230 -2510
rect 38180 -2590 38190 -2520
rect 38180 -2610 38230 -2590
rect 38180 -2680 38190 -2610
rect 38180 -2700 38230 -2680
rect 38180 -2770 38190 -2700
rect 38470 -2750 38500 -2510
rect 38260 -2770 38280 -2750
rect 38350 -2770 38370 -2750
rect 38440 -2770 38500 -2750
rect 38180 -2790 38500 -2770
rect 38180 -2860 38190 -2790
rect 38260 -2840 38280 -2790
rect 38350 -2840 38370 -2790
rect 38440 -2840 38500 -2790
rect 38180 -2880 38230 -2860
rect 38180 -2950 38190 -2880
rect 38180 -2970 38230 -2950
rect 38180 -3040 38190 -2970
rect 38180 -3060 38230 -3040
rect 38180 -3130 38190 -3060
rect 38470 -3080 38500 -2840
rect 38260 -3130 38280 -3080
rect 38350 -3130 38370 -3080
rect 38440 -3130 38500 -3080
rect 38180 -3150 38500 -3130
rect 38180 -3220 38190 -3150
rect 38260 -3170 38280 -3150
rect 38350 -3170 38370 -3150
rect 38440 -3170 38500 -3150
rect 38180 -3240 38230 -3220
rect 38180 -3310 38190 -3240
rect 38180 -3330 38230 -3310
rect 38180 -3400 38190 -3330
rect 38180 -3410 38230 -3400
rect 38470 -3410 38500 -3170
rect 38180 -3460 38500 -3410
rect 38180 -3530 38190 -3460
rect 38260 -3530 38280 -3460
rect 38350 -3530 38370 -3460
rect 38440 -3530 38500 -3460
rect 38180 -3540 38500 -3530
rect 38180 -3550 38230 -3540
rect 38180 -3620 38190 -3550
rect 38180 -3640 38230 -3620
rect 38180 -3710 38190 -3640
rect 38180 -3730 38230 -3710
rect 38180 -3800 38190 -3730
rect 38470 -3780 38500 -3540
rect 38260 -3800 38280 -3780
rect 38350 -3800 38370 -3780
rect 38440 -3800 38500 -3780
rect 38180 -3820 38500 -3800
rect 38180 -3890 38190 -3820
rect 38260 -3870 38280 -3820
rect 38350 -3870 38370 -3820
rect 38440 -3870 38500 -3820
rect 38180 -3910 38230 -3890
rect 38180 -3980 38190 -3910
rect 38180 -4000 38230 -3980
rect 38180 -4070 38190 -4000
rect 38180 -4090 38230 -4070
rect 38180 -4160 38190 -4090
rect 38470 -4110 38500 -3870
rect 38260 -4160 38280 -4110
rect 38350 -4160 38370 -4110
rect 38440 -4160 38500 -4110
rect 38180 -4180 38500 -4160
rect 38180 -4250 38190 -4180
rect 38260 -4200 38280 -4180
rect 38350 -4200 38370 -4180
rect 38440 -4200 38500 -4180
rect 38180 -4270 38230 -4250
rect 38180 -4340 38190 -4270
rect 38180 -4360 38230 -4340
rect 38180 -4430 38190 -4360
rect 38180 -4440 38230 -4430
rect 38470 -4440 38500 -4200
rect 38180 -4450 38500 -4440
rect 38180 -4520 38190 -4450
rect 38260 -4520 38280 -4450
rect 38350 -4520 38370 -4450
rect 38440 -4520 38500 -4450
rect 38180 -4530 38500 -4520
rect 38180 -4540 38230 -4530
rect 38180 -4610 38190 -4540
rect 38180 -4630 38230 -4610
rect 38180 -4700 38190 -4630
rect 38180 -4720 38230 -4700
rect 38180 -4790 38190 -4720
rect 38470 -4770 38500 -4530
rect 38260 -4790 38280 -4770
rect 38350 -4790 38370 -4770
rect 38440 -4790 38500 -4770
rect 38180 -4810 38500 -4790
rect 38180 -4880 38190 -4810
rect 38260 -4860 38280 -4810
rect 38350 -4860 38370 -4810
rect 38440 -4860 38500 -4810
rect 38180 -4900 38230 -4880
rect 38180 -4970 38190 -4900
rect 38180 -4990 38230 -4970
rect 38180 -5060 38190 -4990
rect 38180 -5080 38230 -5060
rect 38180 -5150 38190 -5080
rect 38470 -5100 38500 -4860
rect 38260 -5150 38280 -5100
rect 38350 -5150 38370 -5100
rect 38440 -5150 38500 -5100
rect 38180 -5170 38500 -5150
rect 38180 -5240 38190 -5170
rect 38260 -5190 38280 -5170
rect 38350 -5190 38370 -5170
rect 38440 -5190 38500 -5170
rect 38180 -5260 38230 -5240
rect 38180 -5330 38190 -5260
rect 38180 -5350 38230 -5330
rect 38180 -5420 38190 -5350
rect 38180 -5430 38230 -5420
rect 38470 -5430 38500 -5190
rect 38180 -5440 38500 -5430
rect 38180 -5510 38190 -5440
rect 38260 -5510 38280 -5440
rect 38350 -5510 38370 -5440
rect 38440 -5510 38500 -5440
rect 38180 -5520 38500 -5510
rect 38180 -5530 38230 -5520
rect 38180 -5600 38190 -5530
rect 38180 -5620 38230 -5600
rect 38180 -5690 38190 -5620
rect 38180 -5710 38230 -5690
rect 38180 -5780 38190 -5710
rect 38470 -5760 38500 -5520
rect 38260 -5780 38280 -5760
rect 38350 -5780 38370 -5760
rect 38440 -5780 38500 -5760
rect 38180 -5800 38500 -5780
rect 38180 -5870 38190 -5800
rect 38260 -5850 38280 -5800
rect 38350 -5850 38370 -5800
rect 38440 -5850 38500 -5800
rect 38180 -5890 38230 -5870
rect 38180 -5960 38190 -5890
rect 38180 -5980 38230 -5960
rect 38180 -6050 38190 -5980
rect 38180 -6070 38230 -6050
rect 38180 -6140 38190 -6070
rect 38470 -6090 38500 -5850
rect 38260 -6140 38280 -6090
rect 38350 -6140 38370 -6090
rect 38440 -6140 38500 -6090
rect 38180 -6160 38500 -6140
rect 38180 -6230 38190 -6160
rect 38260 -6180 38280 -6160
rect 38350 -6180 38370 -6160
rect 38440 -6180 38500 -6160
rect 38180 -6250 38230 -6230
rect 38180 -6320 38190 -6250
rect 38180 -6340 38230 -6320
rect 38180 -6410 38190 -6340
rect 38180 -6420 38230 -6410
rect 38470 -6420 38500 -6180
rect 38180 -6450 38500 -6420
rect 30680 -10520 31010 -10510
rect 30680 -10590 30700 -10520
rect 30770 -10590 31010 -10520
rect 30680 -10630 31010 -10590
rect 30680 -10700 30700 -10630
rect 30770 -10700 31010 -10630
rect 30680 -10740 31010 -10700
rect 30680 -10810 30700 -10740
rect 30770 -10810 31010 -10740
rect 30680 -10830 31010 -10810
rect 27015 -11105 30477 -10995
rect 27015 -11600 27125 -11105
rect 26680 -11710 27160 -11600
rect 1510 -12240 3110 -12220
rect 1510 -12300 1690 -12240
rect 1930 -12300 2020 -12240
rect 2260 -12300 2360 -12240
rect 2600 -12300 2690 -12240
rect 2930 -12300 3110 -12240
rect 1510 -12370 1540 -12300
rect 1610 -12370 1650 -12300
rect 1940 -12370 1980 -12300
rect 2270 -12370 2310 -12300
rect 2600 -12370 2640 -12300
rect 2930 -12370 2970 -12300
rect 3040 -12370 3110 -12300
rect 1510 -12410 1690 -12370
rect 1930 -12410 2020 -12370
rect 2260 -12410 2360 -12370
rect 2600 -12410 2690 -12370
rect 2930 -12410 3110 -12370
rect 1510 -12480 1540 -12410
rect 1610 -12480 1650 -12410
rect 1940 -12480 1980 -12410
rect 2270 -12480 2310 -12410
rect 2600 -12480 2640 -12410
rect 2930 -12480 2970 -12410
rect 3040 -12480 3110 -12410
rect 1510 -12510 3110 -12480
rect 11790 -12240 13390 -12220
rect 11790 -12300 11970 -12240
rect 12210 -12300 12300 -12240
rect 12540 -12300 12640 -12240
rect 12880 -12300 12970 -12240
rect 13210 -12300 13390 -12240
rect 11790 -12370 11820 -12300
rect 11890 -12370 11930 -12300
rect 12220 -12370 12260 -12300
rect 12550 -12370 12590 -12300
rect 12880 -12370 12920 -12300
rect 13210 -12370 13250 -12300
rect 13320 -12370 13390 -12300
rect 11790 -12410 11970 -12370
rect 12210 -12410 12300 -12370
rect 12540 -12410 12640 -12370
rect 12880 -12410 12970 -12370
rect 13210 -12410 13390 -12370
rect 11790 -12480 11820 -12410
rect 11890 -12480 11930 -12410
rect 12220 -12480 12260 -12410
rect 12550 -12480 12590 -12410
rect 12880 -12480 12920 -12410
rect 13210 -12480 13250 -12410
rect 13320 -12480 13390 -12410
rect 11790 -12510 13390 -12480
rect 21610 -14020 21930 -13990
rect 21610 -14090 21630 -14020
rect 21700 -14030 21730 -14020
rect 21800 -14030 21830 -14020
rect 21900 -14090 21930 -14020
rect 21610 -14120 21650 -14090
rect 21890 -14120 21930 -14090
rect 21610 -14190 21630 -14120
rect 21900 -14190 21930 -14120
rect 21610 -14220 21650 -14190
rect 21890 -14220 21930 -14190
rect 21610 -14290 21630 -14220
rect 21700 -14290 21730 -14270
rect 21800 -14290 21830 -14270
rect 21900 -14290 21930 -14220
rect 21610 -14310 21930 -14290
rect 22900 -14870 23220 -14840
rect 22900 -14940 22920 -14870
rect 22990 -14940 23020 -14870
rect 23090 -14940 23120 -14870
rect 23190 -14940 23220 -14870
rect 22900 -14970 23220 -14940
rect 22900 -15040 22920 -14970
rect 22990 -15040 23020 -14970
rect 23090 -15040 23120 -14970
rect 23190 -15040 23220 -14970
rect 22900 -15070 23220 -15040
rect 22900 -15140 22920 -15070
rect 22990 -15140 23020 -15070
rect 23090 -15140 23120 -15070
rect 23190 -15140 23220 -15070
rect 22900 -16370 23220 -15140
rect 22900 -16690 30930 -16370
rect 26480 -17620 26960 -17500
rect 26480 -17730 26600 -17620
rect -2710 -17750 26600 -17730
rect -2710 -17820 6460 -17750
rect 6530 -17820 6560 -17750
rect 6630 -17820 6660 -17750
rect 6730 -17820 8170 -17750
rect 8240 -17820 8270 -17750
rect 8340 -17820 8370 -17750
rect 8440 -17820 26600 -17750
rect -2710 -17850 26600 -17820
rect 6440 -17860 6750 -17850
rect 6440 -17930 6460 -17860
rect 6530 -17930 6560 -17860
rect 6630 -17930 6660 -17860
rect 6730 -17930 6750 -17860
rect 6440 -17970 6750 -17930
rect 6440 -18040 6460 -17970
rect 6530 -18040 6560 -17970
rect 6630 -18040 6660 -17970
rect 6730 -18040 6750 -17970
rect 6440 -18080 6750 -18040
rect 6440 -18150 6460 -18080
rect 6530 -18150 6560 -18080
rect 6630 -18150 6660 -18080
rect 6730 -18150 6750 -18080
rect 6440 -18170 6750 -18150
rect 8150 -17860 8460 -17850
rect 8150 -17930 8170 -17860
rect 8240 -17930 8270 -17860
rect 8340 -17930 8370 -17860
rect 8440 -17930 8460 -17860
rect 8150 -17970 8460 -17930
rect 8150 -18040 8170 -17970
rect 8240 -18040 8270 -17970
rect 8340 -18040 8370 -17970
rect 8440 -18040 8460 -17970
rect 8150 -18080 8460 -18040
rect 8150 -18150 8170 -18080
rect 8240 -18150 8270 -18080
rect 8340 -18150 8370 -18080
rect 8440 -18150 8460 -18080
rect 8150 -18170 8460 -18150
rect 21610 -20100 21930 -20070
rect 21610 -20170 21630 -20100
rect 21700 -20110 21730 -20100
rect 21800 -20110 21830 -20100
rect 21900 -20170 21930 -20100
rect 21610 -20200 21650 -20170
rect 21890 -20200 21930 -20170
rect 21610 -20270 21630 -20200
rect 21900 -20270 21930 -20200
rect 21610 -20300 21650 -20270
rect 21890 -20300 21930 -20270
rect 21610 -20370 21630 -20300
rect 21700 -20370 21730 -20350
rect 21800 -20370 21830 -20350
rect 21900 -20370 21930 -20300
rect 21610 -20390 21930 -20370
rect 22680 -20730 23000 -20700
rect 22680 -20800 22700 -20730
rect 22770 -20800 22800 -20730
rect 22870 -20800 22900 -20730
rect 22970 -20800 23000 -20730
rect 22680 -20830 23000 -20800
rect 22680 -20900 22700 -20830
rect 22770 -20900 22800 -20830
rect 22870 -20900 22900 -20830
rect 22970 -20900 23000 -20830
rect 22680 -20930 23000 -20900
rect 22680 -21000 22700 -20930
rect 22770 -21000 22800 -20930
rect 22870 -21000 22900 -20930
rect 22970 -21000 23000 -20930
rect 22680 -22230 23000 -21000
rect 22680 -22550 30710 -22230
rect 1550 -22660 3150 -22630
rect 1550 -22730 1620 -22660
rect 1690 -22730 1730 -22660
rect 2020 -22730 2060 -22660
rect 2350 -22730 2390 -22660
rect 2680 -22730 2720 -22660
rect 3010 -22730 3050 -22660
rect 3120 -22730 3150 -22660
rect 1550 -22770 1730 -22730
rect 1970 -22770 2060 -22730
rect 2300 -22770 2400 -22730
rect 2640 -22770 2730 -22730
rect 2970 -22770 3150 -22730
rect 1550 -22840 1620 -22770
rect 1690 -22840 1730 -22770
rect 2020 -22840 2060 -22770
rect 2350 -22840 2390 -22770
rect 2680 -22840 2720 -22770
rect 3010 -22840 3050 -22770
rect 3120 -22840 3150 -22770
rect 1550 -22900 1730 -22840
rect 1970 -22900 2060 -22840
rect 2300 -22900 2400 -22840
rect 2640 -22900 2730 -22840
rect 2970 -22900 3150 -22840
rect 1550 -22910 3150 -22900
rect 11750 -22660 13350 -22630
rect 11750 -22730 11820 -22660
rect 11890 -22730 11930 -22660
rect 12220 -22730 12260 -22660
rect 12550 -22730 12590 -22660
rect 12880 -22730 12920 -22660
rect 13210 -22730 13250 -22660
rect 13320 -22730 13350 -22660
rect 11750 -22770 11930 -22730
rect 12170 -22770 12260 -22730
rect 12500 -22770 12600 -22730
rect 12840 -22770 12930 -22730
rect 13170 -22770 13350 -22730
rect 11750 -22840 11820 -22770
rect 11890 -22840 11930 -22770
rect 12220 -22840 12260 -22770
rect 12550 -22840 12590 -22770
rect 12880 -22840 12920 -22770
rect 13210 -22840 13250 -22770
rect 13320 -22840 13350 -22770
rect 11750 -22900 11930 -22840
rect 12170 -22900 12260 -22840
rect 12500 -22900 12600 -22840
rect 12840 -22900 12930 -22840
rect 13170 -22900 13350 -22840
rect 11750 -22910 13350 -22900
<< via4 >>
rect -5180 21580 -4940 21610
rect -4850 21580 -4610 21610
rect -4520 21580 -4280 21610
rect -4190 21580 -3950 21610
rect -3860 21580 -3620 21610
rect -3530 21580 -3290 21610
rect -3200 21580 -2960 21610
rect -2870 21580 -2630 21610
rect -2540 21580 -2300 21610
rect -2170 21580 -1930 21610
rect -1840 21580 -1600 21610
rect -1510 21580 -1270 21610
rect -1180 21580 -940 21610
rect -850 21580 -610 21610
rect -520 21580 -280 21610
rect -190 21580 50 21610
rect 140 21580 380 21610
rect 470 21580 710 21610
rect 840 21580 1080 21610
rect 1170 21580 1410 21610
rect 1500 21580 1740 21610
rect 1830 21580 2070 21610
rect 2160 21580 2400 21610
rect 2490 21580 2730 21610
rect 2820 21580 3060 21610
rect 3150 21580 3390 21610
rect 3480 21580 3720 21610
rect 3850 21580 4090 21610
rect 4180 21580 4420 21610
rect 4510 21580 4750 21610
rect 4840 21580 5080 21610
rect 5170 21580 5410 21610
rect 5500 21580 5740 21610
rect 5830 21580 6070 21610
rect 6160 21580 6400 21610
rect 6490 21580 6730 21610
rect -5180 21510 -5170 21580
rect -5170 21510 -5100 21580
rect -5100 21510 -5080 21580
rect -5080 21510 -5010 21580
rect -5010 21510 -4990 21580
rect -4990 21510 -4940 21580
rect -4850 21510 -4830 21580
rect -4830 21510 -4810 21580
rect -4810 21510 -4740 21580
rect -4740 21510 -4720 21580
rect -4720 21510 -4650 21580
rect -4650 21510 -4630 21580
rect -4630 21510 -4610 21580
rect -4520 21510 -4470 21580
rect -4470 21510 -4450 21580
rect -4450 21510 -4380 21580
rect -4380 21510 -4360 21580
rect -4360 21510 -4290 21580
rect -4290 21510 -4280 21580
rect -4190 21510 -4180 21580
rect -4180 21510 -4110 21580
rect -4110 21510 -4090 21580
rect -4090 21510 -4020 21580
rect -4020 21510 -4000 21580
rect -4000 21510 -3950 21580
rect -3860 21510 -3840 21580
rect -3840 21510 -3820 21580
rect -3820 21510 -3750 21580
rect -3750 21510 -3730 21580
rect -3730 21510 -3660 21580
rect -3660 21510 -3640 21580
rect -3640 21510 -3620 21580
rect -3530 21510 -3480 21580
rect -3480 21510 -3460 21580
rect -3460 21510 -3390 21580
rect -3390 21510 -3370 21580
rect -3370 21510 -3300 21580
rect -3300 21510 -3290 21580
rect -3200 21510 -3190 21580
rect -3190 21510 -3120 21580
rect -3120 21510 -3100 21580
rect -3100 21510 -3030 21580
rect -3030 21510 -3010 21580
rect -3010 21510 -2960 21580
rect -2870 21510 -2850 21580
rect -2850 21510 -2830 21580
rect -2830 21510 -2760 21580
rect -2760 21510 -2740 21580
rect -2740 21510 -2670 21580
rect -2670 21510 -2650 21580
rect -2650 21510 -2630 21580
rect -2540 21510 -2490 21580
rect -2490 21510 -2470 21580
rect -2470 21510 -2400 21580
rect -2400 21510 -2380 21580
rect -2380 21510 -2310 21580
rect -2310 21510 -2300 21580
rect -2170 21510 -2160 21580
rect -2160 21510 -2090 21580
rect -2090 21510 -2070 21580
rect -2070 21510 -2000 21580
rect -2000 21510 -1980 21580
rect -1980 21510 -1930 21580
rect -1840 21510 -1820 21580
rect -1820 21510 -1800 21580
rect -1800 21510 -1730 21580
rect -1730 21510 -1710 21580
rect -1710 21510 -1640 21580
rect -1640 21510 -1620 21580
rect -1620 21510 -1600 21580
rect -1510 21510 -1460 21580
rect -1460 21510 -1440 21580
rect -1440 21510 -1370 21580
rect -1370 21510 -1350 21580
rect -1350 21510 -1280 21580
rect -1280 21510 -1270 21580
rect -1180 21510 -1170 21580
rect -1170 21510 -1100 21580
rect -1100 21510 -1080 21580
rect -1080 21510 -1010 21580
rect -1010 21510 -990 21580
rect -990 21510 -940 21580
rect -850 21510 -830 21580
rect -830 21510 -810 21580
rect -810 21510 -740 21580
rect -740 21510 -720 21580
rect -720 21510 -650 21580
rect -650 21510 -630 21580
rect -630 21510 -610 21580
rect -520 21510 -470 21580
rect -470 21510 -450 21580
rect -450 21510 -380 21580
rect -380 21510 -360 21580
rect -360 21510 -290 21580
rect -290 21510 -280 21580
rect -190 21510 -180 21580
rect -180 21510 -110 21580
rect -110 21510 -90 21580
rect -90 21510 -20 21580
rect -20 21510 0 21580
rect 0 21510 50 21580
rect 140 21510 160 21580
rect 160 21510 180 21580
rect 180 21510 250 21580
rect 250 21510 270 21580
rect 270 21510 340 21580
rect 340 21510 360 21580
rect 360 21510 380 21580
rect 470 21510 520 21580
rect 520 21510 540 21580
rect 540 21510 610 21580
rect 610 21510 630 21580
rect 630 21510 700 21580
rect 700 21510 710 21580
rect 840 21510 850 21580
rect 850 21510 920 21580
rect 920 21510 940 21580
rect 940 21510 1010 21580
rect 1010 21510 1030 21580
rect 1030 21510 1080 21580
rect 1170 21510 1190 21580
rect 1190 21510 1210 21580
rect 1210 21510 1280 21580
rect 1280 21510 1300 21580
rect 1300 21510 1370 21580
rect 1370 21510 1390 21580
rect 1390 21510 1410 21580
rect 1500 21510 1550 21580
rect 1550 21510 1570 21580
rect 1570 21510 1640 21580
rect 1640 21510 1660 21580
rect 1660 21510 1730 21580
rect 1730 21510 1740 21580
rect 1830 21510 1840 21580
rect 1840 21510 1910 21580
rect 1910 21510 1930 21580
rect 1930 21510 2000 21580
rect 2000 21510 2020 21580
rect 2020 21510 2070 21580
rect 2160 21510 2180 21580
rect 2180 21510 2200 21580
rect 2200 21510 2270 21580
rect 2270 21510 2290 21580
rect 2290 21510 2360 21580
rect 2360 21510 2380 21580
rect 2380 21510 2400 21580
rect 2490 21510 2540 21580
rect 2540 21510 2560 21580
rect 2560 21510 2630 21580
rect 2630 21510 2650 21580
rect 2650 21510 2720 21580
rect 2720 21510 2730 21580
rect 2820 21510 2830 21580
rect 2830 21510 2900 21580
rect 2900 21510 2920 21580
rect 2920 21510 2990 21580
rect 2990 21510 3010 21580
rect 3010 21510 3060 21580
rect 3150 21510 3170 21580
rect 3170 21510 3190 21580
rect 3190 21510 3260 21580
rect 3260 21510 3280 21580
rect 3280 21510 3350 21580
rect 3350 21510 3370 21580
rect 3370 21510 3390 21580
rect 3480 21510 3530 21580
rect 3530 21510 3550 21580
rect 3550 21510 3620 21580
rect 3620 21510 3640 21580
rect 3640 21510 3710 21580
rect 3710 21510 3720 21580
rect 3850 21510 3860 21580
rect 3860 21510 3930 21580
rect 3930 21510 3950 21580
rect 3950 21510 4020 21580
rect 4020 21510 4040 21580
rect 4040 21510 4090 21580
rect 4180 21510 4200 21580
rect 4200 21510 4220 21580
rect 4220 21510 4290 21580
rect 4290 21510 4310 21580
rect 4310 21510 4380 21580
rect 4380 21510 4400 21580
rect 4400 21510 4420 21580
rect 4510 21510 4560 21580
rect 4560 21510 4580 21580
rect 4580 21510 4650 21580
rect 4650 21510 4670 21580
rect 4670 21510 4740 21580
rect 4740 21510 4750 21580
rect 4840 21510 4850 21580
rect 4850 21510 4920 21580
rect 4920 21510 4940 21580
rect 4940 21510 5010 21580
rect 5010 21510 5030 21580
rect 5030 21510 5080 21580
rect 5170 21510 5190 21580
rect 5190 21510 5210 21580
rect 5210 21510 5280 21580
rect 5280 21510 5300 21580
rect 5300 21510 5370 21580
rect 5370 21510 5390 21580
rect 5390 21510 5410 21580
rect 5500 21510 5550 21580
rect 5550 21510 5570 21580
rect 5570 21510 5640 21580
rect 5640 21510 5660 21580
rect 5660 21510 5730 21580
rect 5730 21510 5740 21580
rect 5830 21510 5840 21580
rect 5840 21510 5910 21580
rect 5910 21510 5930 21580
rect 5930 21510 6000 21580
rect 6000 21510 6020 21580
rect 6020 21510 6070 21580
rect 6160 21510 6180 21580
rect 6180 21510 6200 21580
rect 6200 21510 6270 21580
rect 6270 21510 6290 21580
rect 6290 21510 6360 21580
rect 6360 21510 6380 21580
rect 6380 21510 6400 21580
rect 6490 21510 6540 21580
rect 6540 21510 6560 21580
rect 6560 21510 6630 21580
rect 6630 21510 6650 21580
rect 6650 21510 6720 21580
rect 6720 21510 6730 21580
rect -5180 21490 -4940 21510
rect -4850 21490 -4610 21510
rect -4520 21490 -4280 21510
rect -4190 21490 -3950 21510
rect -3860 21490 -3620 21510
rect -3530 21490 -3290 21510
rect -3200 21490 -2960 21510
rect -2870 21490 -2630 21510
rect -2540 21490 -2300 21510
rect -2170 21490 -1930 21510
rect -1840 21490 -1600 21510
rect -1510 21490 -1270 21510
rect -1180 21490 -940 21510
rect -850 21490 -610 21510
rect -520 21490 -280 21510
rect -190 21490 50 21510
rect 140 21490 380 21510
rect 470 21490 710 21510
rect 840 21490 1080 21510
rect 1170 21490 1410 21510
rect 1500 21490 1740 21510
rect 1830 21490 2070 21510
rect 2160 21490 2400 21510
rect 2490 21490 2730 21510
rect 2820 21490 3060 21510
rect 3150 21490 3390 21510
rect 3480 21490 3720 21510
rect 3850 21490 4090 21510
rect 4180 21490 4420 21510
rect 4510 21490 4750 21510
rect 4840 21490 5080 21510
rect 5170 21490 5410 21510
rect 5500 21490 5740 21510
rect 5830 21490 6070 21510
rect 6160 21490 6400 21510
rect 6490 21490 6730 21510
rect -5180 21420 -5170 21490
rect -5170 21420 -5100 21490
rect -5100 21420 -5080 21490
rect -5080 21420 -5010 21490
rect -5010 21420 -4990 21490
rect -4990 21420 -4940 21490
rect -4850 21420 -4830 21490
rect -4830 21420 -4810 21490
rect -4810 21420 -4740 21490
rect -4740 21420 -4720 21490
rect -4720 21420 -4650 21490
rect -4650 21420 -4630 21490
rect -4630 21420 -4610 21490
rect -4520 21420 -4470 21490
rect -4470 21420 -4450 21490
rect -4450 21420 -4380 21490
rect -4380 21420 -4360 21490
rect -4360 21420 -4290 21490
rect -4290 21420 -4280 21490
rect -4190 21420 -4180 21490
rect -4180 21420 -4110 21490
rect -4110 21420 -4090 21490
rect -4090 21420 -4020 21490
rect -4020 21420 -4000 21490
rect -4000 21420 -3950 21490
rect -3860 21420 -3840 21490
rect -3840 21420 -3820 21490
rect -3820 21420 -3750 21490
rect -3750 21420 -3730 21490
rect -3730 21420 -3660 21490
rect -3660 21420 -3640 21490
rect -3640 21420 -3620 21490
rect -3530 21420 -3480 21490
rect -3480 21420 -3460 21490
rect -3460 21420 -3390 21490
rect -3390 21420 -3370 21490
rect -3370 21420 -3300 21490
rect -3300 21420 -3290 21490
rect -3200 21420 -3190 21490
rect -3190 21420 -3120 21490
rect -3120 21420 -3100 21490
rect -3100 21420 -3030 21490
rect -3030 21420 -3010 21490
rect -3010 21420 -2960 21490
rect -2870 21420 -2850 21490
rect -2850 21420 -2830 21490
rect -2830 21420 -2760 21490
rect -2760 21420 -2740 21490
rect -2740 21420 -2670 21490
rect -2670 21420 -2650 21490
rect -2650 21420 -2630 21490
rect -2540 21420 -2490 21490
rect -2490 21420 -2470 21490
rect -2470 21420 -2400 21490
rect -2400 21420 -2380 21490
rect -2380 21420 -2310 21490
rect -2310 21420 -2300 21490
rect -2170 21420 -2160 21490
rect -2160 21420 -2090 21490
rect -2090 21420 -2070 21490
rect -2070 21420 -2000 21490
rect -2000 21420 -1980 21490
rect -1980 21420 -1930 21490
rect -1840 21420 -1820 21490
rect -1820 21420 -1800 21490
rect -1800 21420 -1730 21490
rect -1730 21420 -1710 21490
rect -1710 21420 -1640 21490
rect -1640 21420 -1620 21490
rect -1620 21420 -1600 21490
rect -1510 21420 -1460 21490
rect -1460 21420 -1440 21490
rect -1440 21420 -1370 21490
rect -1370 21420 -1350 21490
rect -1350 21420 -1280 21490
rect -1280 21420 -1270 21490
rect -1180 21420 -1170 21490
rect -1170 21420 -1100 21490
rect -1100 21420 -1080 21490
rect -1080 21420 -1010 21490
rect -1010 21420 -990 21490
rect -990 21420 -940 21490
rect -850 21420 -830 21490
rect -830 21420 -810 21490
rect -810 21420 -740 21490
rect -740 21420 -720 21490
rect -720 21420 -650 21490
rect -650 21420 -630 21490
rect -630 21420 -610 21490
rect -520 21420 -470 21490
rect -470 21420 -450 21490
rect -450 21420 -380 21490
rect -380 21420 -360 21490
rect -360 21420 -290 21490
rect -290 21420 -280 21490
rect -190 21420 -180 21490
rect -180 21420 -110 21490
rect -110 21420 -90 21490
rect -90 21420 -20 21490
rect -20 21420 0 21490
rect 0 21420 50 21490
rect 140 21420 160 21490
rect 160 21420 180 21490
rect 180 21420 250 21490
rect 250 21420 270 21490
rect 270 21420 340 21490
rect 340 21420 360 21490
rect 360 21420 380 21490
rect 470 21420 520 21490
rect 520 21420 540 21490
rect 540 21420 610 21490
rect 610 21420 630 21490
rect 630 21420 700 21490
rect 700 21420 710 21490
rect 840 21420 850 21490
rect 850 21420 920 21490
rect 920 21420 940 21490
rect 940 21420 1010 21490
rect 1010 21420 1030 21490
rect 1030 21420 1080 21490
rect 1170 21420 1190 21490
rect 1190 21420 1210 21490
rect 1210 21420 1280 21490
rect 1280 21420 1300 21490
rect 1300 21420 1370 21490
rect 1370 21420 1390 21490
rect 1390 21420 1410 21490
rect 1500 21420 1550 21490
rect 1550 21420 1570 21490
rect 1570 21420 1640 21490
rect 1640 21420 1660 21490
rect 1660 21420 1730 21490
rect 1730 21420 1740 21490
rect 1830 21420 1840 21490
rect 1840 21420 1910 21490
rect 1910 21420 1930 21490
rect 1930 21420 2000 21490
rect 2000 21420 2020 21490
rect 2020 21420 2070 21490
rect 2160 21420 2180 21490
rect 2180 21420 2200 21490
rect 2200 21420 2270 21490
rect 2270 21420 2290 21490
rect 2290 21420 2360 21490
rect 2360 21420 2380 21490
rect 2380 21420 2400 21490
rect 2490 21420 2540 21490
rect 2540 21420 2560 21490
rect 2560 21420 2630 21490
rect 2630 21420 2650 21490
rect 2650 21420 2720 21490
rect 2720 21420 2730 21490
rect 2820 21420 2830 21490
rect 2830 21420 2900 21490
rect 2900 21420 2920 21490
rect 2920 21420 2990 21490
rect 2990 21420 3010 21490
rect 3010 21420 3060 21490
rect 3150 21420 3170 21490
rect 3170 21420 3190 21490
rect 3190 21420 3260 21490
rect 3260 21420 3280 21490
rect 3280 21420 3350 21490
rect 3350 21420 3370 21490
rect 3370 21420 3390 21490
rect 3480 21420 3530 21490
rect 3530 21420 3550 21490
rect 3550 21420 3620 21490
rect 3620 21420 3640 21490
rect 3640 21420 3710 21490
rect 3710 21420 3720 21490
rect 3850 21420 3860 21490
rect 3860 21420 3930 21490
rect 3930 21420 3950 21490
rect 3950 21420 4020 21490
rect 4020 21420 4040 21490
rect 4040 21420 4090 21490
rect 4180 21420 4200 21490
rect 4200 21420 4220 21490
rect 4220 21420 4290 21490
rect 4290 21420 4310 21490
rect 4310 21420 4380 21490
rect 4380 21420 4400 21490
rect 4400 21420 4420 21490
rect 4510 21420 4560 21490
rect 4560 21420 4580 21490
rect 4580 21420 4650 21490
rect 4650 21420 4670 21490
rect 4670 21420 4740 21490
rect 4740 21420 4750 21490
rect 4840 21420 4850 21490
rect 4850 21420 4920 21490
rect 4920 21420 4940 21490
rect 4940 21420 5010 21490
rect 5010 21420 5030 21490
rect 5030 21420 5080 21490
rect 5170 21420 5190 21490
rect 5190 21420 5210 21490
rect 5210 21420 5280 21490
rect 5280 21420 5300 21490
rect 5300 21420 5370 21490
rect 5370 21420 5390 21490
rect 5390 21420 5410 21490
rect 5500 21420 5550 21490
rect 5550 21420 5570 21490
rect 5570 21420 5640 21490
rect 5640 21420 5660 21490
rect 5660 21420 5730 21490
rect 5730 21420 5740 21490
rect 5830 21420 5840 21490
rect 5840 21420 5910 21490
rect 5910 21420 5930 21490
rect 5930 21420 6000 21490
rect 6000 21420 6020 21490
rect 6020 21420 6070 21490
rect 6160 21420 6180 21490
rect 6180 21420 6200 21490
rect 6200 21420 6270 21490
rect 6270 21420 6290 21490
rect 6290 21420 6360 21490
rect 6360 21420 6380 21490
rect 6380 21420 6400 21490
rect 6490 21420 6540 21490
rect 6540 21420 6560 21490
rect 6560 21420 6630 21490
rect 6630 21420 6650 21490
rect 6650 21420 6720 21490
rect 6720 21420 6730 21490
rect -5180 21400 -4940 21420
rect -4850 21400 -4610 21420
rect -4520 21400 -4280 21420
rect -4190 21400 -3950 21420
rect -3860 21400 -3620 21420
rect -3530 21400 -3290 21420
rect -3200 21400 -2960 21420
rect -2870 21400 -2630 21420
rect -2540 21400 -2300 21420
rect -2170 21400 -1930 21420
rect -1840 21400 -1600 21420
rect -1510 21400 -1270 21420
rect -1180 21400 -940 21420
rect -850 21400 -610 21420
rect -520 21400 -280 21420
rect -190 21400 50 21420
rect 140 21400 380 21420
rect 470 21400 710 21420
rect 840 21400 1080 21420
rect 1170 21400 1410 21420
rect 1500 21400 1740 21420
rect 1830 21400 2070 21420
rect 2160 21400 2400 21420
rect 2490 21400 2730 21420
rect 2820 21400 3060 21420
rect 3150 21400 3390 21420
rect 3480 21400 3720 21420
rect 3850 21400 4090 21420
rect 4180 21400 4420 21420
rect 4510 21400 4750 21420
rect 4840 21400 5080 21420
rect 5170 21400 5410 21420
rect 5500 21400 5740 21420
rect 5830 21400 6070 21420
rect 6160 21400 6400 21420
rect 6490 21400 6730 21420
rect -5180 21370 -5170 21400
rect -5170 21370 -5100 21400
rect -5100 21370 -5080 21400
rect -5080 21370 -5010 21400
rect -5010 21370 -4990 21400
rect -4990 21370 -4940 21400
rect -4850 21370 -4830 21400
rect -4830 21370 -4810 21400
rect -4810 21370 -4740 21400
rect -4740 21370 -4720 21400
rect -4720 21370 -4650 21400
rect -4650 21370 -4630 21400
rect -4630 21370 -4610 21400
rect -4520 21370 -4470 21400
rect -4470 21370 -4450 21400
rect -4450 21370 -4380 21400
rect -4380 21370 -4360 21400
rect -4360 21370 -4290 21400
rect -4290 21370 -4280 21400
rect -4190 21370 -4180 21400
rect -4180 21370 -4110 21400
rect -4110 21370 -4090 21400
rect -4090 21370 -4020 21400
rect -4020 21370 -4000 21400
rect -4000 21370 -3950 21400
rect -3860 21370 -3840 21400
rect -3840 21370 -3820 21400
rect -3820 21370 -3750 21400
rect -3750 21370 -3730 21400
rect -3730 21370 -3660 21400
rect -3660 21370 -3640 21400
rect -3640 21370 -3620 21400
rect -3530 21370 -3480 21400
rect -3480 21370 -3460 21400
rect -3460 21370 -3390 21400
rect -3390 21370 -3370 21400
rect -3370 21370 -3300 21400
rect -3300 21370 -3290 21400
rect -3200 21370 -3190 21400
rect -3190 21370 -3120 21400
rect -3120 21370 -3100 21400
rect -3100 21370 -3030 21400
rect -3030 21370 -3010 21400
rect -3010 21370 -2960 21400
rect -2870 21370 -2850 21400
rect -2850 21370 -2830 21400
rect -2830 21370 -2760 21400
rect -2760 21370 -2740 21400
rect -2740 21370 -2670 21400
rect -2670 21370 -2650 21400
rect -2650 21370 -2630 21400
rect -2540 21370 -2490 21400
rect -2490 21370 -2470 21400
rect -2470 21370 -2400 21400
rect -2400 21370 -2380 21400
rect -2380 21370 -2310 21400
rect -2310 21370 -2300 21400
rect -2170 21370 -2160 21400
rect -2160 21370 -2090 21400
rect -2090 21370 -2070 21400
rect -2070 21370 -2000 21400
rect -2000 21370 -1980 21400
rect -1980 21370 -1930 21400
rect -1840 21370 -1820 21400
rect -1820 21370 -1800 21400
rect -1800 21370 -1730 21400
rect -1730 21370 -1710 21400
rect -1710 21370 -1640 21400
rect -1640 21370 -1620 21400
rect -1620 21370 -1600 21400
rect -1510 21370 -1460 21400
rect -1460 21370 -1440 21400
rect -1440 21370 -1370 21400
rect -1370 21370 -1350 21400
rect -1350 21370 -1280 21400
rect -1280 21370 -1270 21400
rect -1180 21370 -1170 21400
rect -1170 21370 -1100 21400
rect -1100 21370 -1080 21400
rect -1080 21370 -1010 21400
rect -1010 21370 -990 21400
rect -990 21370 -940 21400
rect -850 21370 -830 21400
rect -830 21370 -810 21400
rect -810 21370 -740 21400
rect -740 21370 -720 21400
rect -720 21370 -650 21400
rect -650 21370 -630 21400
rect -630 21370 -610 21400
rect -520 21370 -470 21400
rect -470 21370 -450 21400
rect -450 21370 -380 21400
rect -380 21370 -360 21400
rect -360 21370 -290 21400
rect -290 21370 -280 21400
rect -190 21370 -180 21400
rect -180 21370 -110 21400
rect -110 21370 -90 21400
rect -90 21370 -20 21400
rect -20 21370 0 21400
rect 0 21370 50 21400
rect 140 21370 160 21400
rect 160 21370 180 21400
rect 180 21370 250 21400
rect 250 21370 270 21400
rect 270 21370 340 21400
rect 340 21370 360 21400
rect 360 21370 380 21400
rect 470 21370 520 21400
rect 520 21370 540 21400
rect 540 21370 610 21400
rect 610 21370 630 21400
rect 630 21370 700 21400
rect 700 21370 710 21400
rect 840 21370 850 21400
rect 850 21370 920 21400
rect 920 21370 940 21400
rect 940 21370 1010 21400
rect 1010 21370 1030 21400
rect 1030 21370 1080 21400
rect 1170 21370 1190 21400
rect 1190 21370 1210 21400
rect 1210 21370 1280 21400
rect 1280 21370 1300 21400
rect 1300 21370 1370 21400
rect 1370 21370 1390 21400
rect 1390 21370 1410 21400
rect 1500 21370 1550 21400
rect 1550 21370 1570 21400
rect 1570 21370 1640 21400
rect 1640 21370 1660 21400
rect 1660 21370 1730 21400
rect 1730 21370 1740 21400
rect 1830 21370 1840 21400
rect 1840 21370 1910 21400
rect 1910 21370 1930 21400
rect 1930 21370 2000 21400
rect 2000 21370 2020 21400
rect 2020 21370 2070 21400
rect 2160 21370 2180 21400
rect 2180 21370 2200 21400
rect 2200 21370 2270 21400
rect 2270 21370 2290 21400
rect 2290 21370 2360 21400
rect 2360 21370 2380 21400
rect 2380 21370 2400 21400
rect 2490 21370 2540 21400
rect 2540 21370 2560 21400
rect 2560 21370 2630 21400
rect 2630 21370 2650 21400
rect 2650 21370 2720 21400
rect 2720 21370 2730 21400
rect 2820 21370 2830 21400
rect 2830 21370 2900 21400
rect 2900 21370 2920 21400
rect 2920 21370 2990 21400
rect 2990 21370 3010 21400
rect 3010 21370 3060 21400
rect 3150 21370 3170 21400
rect 3170 21370 3190 21400
rect 3190 21370 3260 21400
rect 3260 21370 3280 21400
rect 3280 21370 3350 21400
rect 3350 21370 3370 21400
rect 3370 21370 3390 21400
rect 3480 21370 3530 21400
rect 3530 21370 3550 21400
rect 3550 21370 3620 21400
rect 3620 21370 3640 21400
rect 3640 21370 3710 21400
rect 3710 21370 3720 21400
rect 3850 21370 3860 21400
rect 3860 21370 3930 21400
rect 3930 21370 3950 21400
rect 3950 21370 4020 21400
rect 4020 21370 4040 21400
rect 4040 21370 4090 21400
rect 4180 21370 4200 21400
rect 4200 21370 4220 21400
rect 4220 21370 4290 21400
rect 4290 21370 4310 21400
rect 4310 21370 4380 21400
rect 4380 21370 4400 21400
rect 4400 21370 4420 21400
rect 4510 21370 4560 21400
rect 4560 21370 4580 21400
rect 4580 21370 4650 21400
rect 4650 21370 4670 21400
rect 4670 21370 4740 21400
rect 4740 21370 4750 21400
rect 4840 21370 4850 21400
rect 4850 21370 4920 21400
rect 4920 21370 4940 21400
rect 4940 21370 5010 21400
rect 5010 21370 5030 21400
rect 5030 21370 5080 21400
rect 5170 21370 5190 21400
rect 5190 21370 5210 21400
rect 5210 21370 5280 21400
rect 5280 21370 5300 21400
rect 5300 21370 5370 21400
rect 5370 21370 5390 21400
rect 5390 21370 5410 21400
rect 5500 21370 5550 21400
rect 5550 21370 5570 21400
rect 5570 21370 5640 21400
rect 5640 21370 5660 21400
rect 5660 21370 5730 21400
rect 5730 21370 5740 21400
rect 5830 21370 5840 21400
rect 5840 21370 5910 21400
rect 5910 21370 5930 21400
rect 5930 21370 6000 21400
rect 6000 21370 6020 21400
rect 6020 21370 6070 21400
rect 6160 21370 6180 21400
rect 6180 21370 6200 21400
rect 6200 21370 6270 21400
rect 6270 21370 6290 21400
rect 6290 21370 6360 21400
rect 6360 21370 6380 21400
rect 6380 21370 6400 21400
rect 6490 21370 6540 21400
rect 6540 21370 6560 21400
rect 6560 21370 6630 21400
rect 6630 21370 6650 21400
rect 6650 21370 6720 21400
rect 6720 21370 6730 21400
rect 8170 21580 8410 21610
rect 8500 21580 8740 21610
rect 8830 21580 9070 21610
rect 9160 21580 9400 21610
rect 9490 21580 9730 21610
rect 9820 21580 10060 21610
rect 10150 21580 10390 21610
rect 10480 21580 10720 21610
rect 10810 21580 11050 21610
rect 11180 21580 11420 21610
rect 11510 21580 11750 21610
rect 11840 21580 12080 21610
rect 12170 21580 12410 21610
rect 12500 21580 12740 21610
rect 12830 21580 13070 21610
rect 13160 21580 13400 21610
rect 13490 21580 13730 21610
rect 13820 21580 14060 21610
rect 14190 21580 14430 21610
rect 14520 21580 14760 21610
rect 14850 21580 15090 21610
rect 15180 21580 15420 21610
rect 15510 21580 15750 21610
rect 15840 21580 16080 21610
rect 16170 21580 16410 21610
rect 16500 21580 16740 21610
rect 16830 21580 17070 21610
rect 17200 21580 17440 21610
rect 17530 21580 17770 21610
rect 17860 21580 18100 21610
rect 18190 21580 18430 21610
rect 18520 21580 18760 21610
rect 18850 21580 19090 21610
rect 19180 21580 19420 21610
rect 19510 21580 19750 21610
rect 19840 21580 20080 21610
rect 8170 21510 8180 21580
rect 8180 21510 8250 21580
rect 8250 21510 8270 21580
rect 8270 21510 8340 21580
rect 8340 21510 8360 21580
rect 8360 21510 8410 21580
rect 8500 21510 8520 21580
rect 8520 21510 8540 21580
rect 8540 21510 8610 21580
rect 8610 21510 8630 21580
rect 8630 21510 8700 21580
rect 8700 21510 8720 21580
rect 8720 21510 8740 21580
rect 8830 21510 8880 21580
rect 8880 21510 8900 21580
rect 8900 21510 8970 21580
rect 8970 21510 8990 21580
rect 8990 21510 9060 21580
rect 9060 21510 9070 21580
rect 9160 21510 9170 21580
rect 9170 21510 9240 21580
rect 9240 21510 9260 21580
rect 9260 21510 9330 21580
rect 9330 21510 9350 21580
rect 9350 21510 9400 21580
rect 9490 21510 9510 21580
rect 9510 21510 9530 21580
rect 9530 21510 9600 21580
rect 9600 21510 9620 21580
rect 9620 21510 9690 21580
rect 9690 21510 9710 21580
rect 9710 21510 9730 21580
rect 9820 21510 9870 21580
rect 9870 21510 9890 21580
rect 9890 21510 9960 21580
rect 9960 21510 9980 21580
rect 9980 21510 10050 21580
rect 10050 21510 10060 21580
rect 10150 21510 10160 21580
rect 10160 21510 10230 21580
rect 10230 21510 10250 21580
rect 10250 21510 10320 21580
rect 10320 21510 10340 21580
rect 10340 21510 10390 21580
rect 10480 21510 10500 21580
rect 10500 21510 10520 21580
rect 10520 21510 10590 21580
rect 10590 21510 10610 21580
rect 10610 21510 10680 21580
rect 10680 21510 10700 21580
rect 10700 21510 10720 21580
rect 10810 21510 10860 21580
rect 10860 21510 10880 21580
rect 10880 21510 10950 21580
rect 10950 21510 10970 21580
rect 10970 21510 11040 21580
rect 11040 21510 11050 21580
rect 11180 21510 11190 21580
rect 11190 21510 11260 21580
rect 11260 21510 11280 21580
rect 11280 21510 11350 21580
rect 11350 21510 11370 21580
rect 11370 21510 11420 21580
rect 11510 21510 11530 21580
rect 11530 21510 11550 21580
rect 11550 21510 11620 21580
rect 11620 21510 11640 21580
rect 11640 21510 11710 21580
rect 11710 21510 11730 21580
rect 11730 21510 11750 21580
rect 11840 21510 11890 21580
rect 11890 21510 11910 21580
rect 11910 21510 11980 21580
rect 11980 21510 12000 21580
rect 12000 21510 12070 21580
rect 12070 21510 12080 21580
rect 12170 21510 12180 21580
rect 12180 21510 12250 21580
rect 12250 21510 12270 21580
rect 12270 21510 12340 21580
rect 12340 21510 12360 21580
rect 12360 21510 12410 21580
rect 12500 21510 12520 21580
rect 12520 21510 12540 21580
rect 12540 21510 12610 21580
rect 12610 21510 12630 21580
rect 12630 21510 12700 21580
rect 12700 21510 12720 21580
rect 12720 21510 12740 21580
rect 12830 21510 12880 21580
rect 12880 21510 12900 21580
rect 12900 21510 12970 21580
rect 12970 21510 12990 21580
rect 12990 21510 13060 21580
rect 13060 21510 13070 21580
rect 13160 21510 13170 21580
rect 13170 21510 13240 21580
rect 13240 21510 13260 21580
rect 13260 21510 13330 21580
rect 13330 21510 13350 21580
rect 13350 21510 13400 21580
rect 13490 21510 13510 21580
rect 13510 21510 13530 21580
rect 13530 21510 13600 21580
rect 13600 21510 13620 21580
rect 13620 21510 13690 21580
rect 13690 21510 13710 21580
rect 13710 21510 13730 21580
rect 13820 21510 13870 21580
rect 13870 21510 13890 21580
rect 13890 21510 13960 21580
rect 13960 21510 13980 21580
rect 13980 21510 14050 21580
rect 14050 21510 14060 21580
rect 14190 21510 14200 21580
rect 14200 21510 14270 21580
rect 14270 21510 14290 21580
rect 14290 21510 14360 21580
rect 14360 21510 14380 21580
rect 14380 21510 14430 21580
rect 14520 21510 14540 21580
rect 14540 21510 14560 21580
rect 14560 21510 14630 21580
rect 14630 21510 14650 21580
rect 14650 21510 14720 21580
rect 14720 21510 14740 21580
rect 14740 21510 14760 21580
rect 14850 21510 14900 21580
rect 14900 21510 14920 21580
rect 14920 21510 14990 21580
rect 14990 21510 15010 21580
rect 15010 21510 15080 21580
rect 15080 21510 15090 21580
rect 15180 21510 15190 21580
rect 15190 21510 15260 21580
rect 15260 21510 15280 21580
rect 15280 21510 15350 21580
rect 15350 21510 15370 21580
rect 15370 21510 15420 21580
rect 15510 21510 15530 21580
rect 15530 21510 15550 21580
rect 15550 21510 15620 21580
rect 15620 21510 15640 21580
rect 15640 21510 15710 21580
rect 15710 21510 15730 21580
rect 15730 21510 15750 21580
rect 15840 21510 15890 21580
rect 15890 21510 15910 21580
rect 15910 21510 15980 21580
rect 15980 21510 16000 21580
rect 16000 21510 16070 21580
rect 16070 21510 16080 21580
rect 16170 21510 16180 21580
rect 16180 21510 16250 21580
rect 16250 21510 16270 21580
rect 16270 21510 16340 21580
rect 16340 21510 16360 21580
rect 16360 21510 16410 21580
rect 16500 21510 16520 21580
rect 16520 21510 16540 21580
rect 16540 21510 16610 21580
rect 16610 21510 16630 21580
rect 16630 21510 16700 21580
rect 16700 21510 16720 21580
rect 16720 21510 16740 21580
rect 16830 21510 16880 21580
rect 16880 21510 16900 21580
rect 16900 21510 16970 21580
rect 16970 21510 16990 21580
rect 16990 21510 17060 21580
rect 17060 21510 17070 21580
rect 17200 21510 17210 21580
rect 17210 21510 17280 21580
rect 17280 21510 17300 21580
rect 17300 21510 17370 21580
rect 17370 21510 17390 21580
rect 17390 21510 17440 21580
rect 17530 21510 17550 21580
rect 17550 21510 17570 21580
rect 17570 21510 17640 21580
rect 17640 21510 17660 21580
rect 17660 21510 17730 21580
rect 17730 21510 17750 21580
rect 17750 21510 17770 21580
rect 17860 21510 17910 21580
rect 17910 21510 17930 21580
rect 17930 21510 18000 21580
rect 18000 21510 18020 21580
rect 18020 21510 18090 21580
rect 18090 21510 18100 21580
rect 18190 21510 18200 21580
rect 18200 21510 18270 21580
rect 18270 21510 18290 21580
rect 18290 21510 18360 21580
rect 18360 21510 18380 21580
rect 18380 21510 18430 21580
rect 18520 21510 18540 21580
rect 18540 21510 18560 21580
rect 18560 21510 18630 21580
rect 18630 21510 18650 21580
rect 18650 21510 18720 21580
rect 18720 21510 18740 21580
rect 18740 21510 18760 21580
rect 18850 21510 18900 21580
rect 18900 21510 18920 21580
rect 18920 21510 18990 21580
rect 18990 21510 19010 21580
rect 19010 21510 19080 21580
rect 19080 21510 19090 21580
rect 19180 21510 19190 21580
rect 19190 21510 19260 21580
rect 19260 21510 19280 21580
rect 19280 21510 19350 21580
rect 19350 21510 19370 21580
rect 19370 21510 19420 21580
rect 19510 21510 19530 21580
rect 19530 21510 19550 21580
rect 19550 21510 19620 21580
rect 19620 21510 19640 21580
rect 19640 21510 19710 21580
rect 19710 21510 19730 21580
rect 19730 21510 19750 21580
rect 19840 21510 19890 21580
rect 19890 21510 19910 21580
rect 19910 21510 19980 21580
rect 19980 21510 20000 21580
rect 20000 21510 20070 21580
rect 20070 21510 20080 21580
rect 8170 21490 8410 21510
rect 8500 21490 8740 21510
rect 8830 21490 9070 21510
rect 9160 21490 9400 21510
rect 9490 21490 9730 21510
rect 9820 21490 10060 21510
rect 10150 21490 10390 21510
rect 10480 21490 10720 21510
rect 10810 21490 11050 21510
rect 11180 21490 11420 21510
rect 11510 21490 11750 21510
rect 11840 21490 12080 21510
rect 12170 21490 12410 21510
rect 12500 21490 12740 21510
rect 12830 21490 13070 21510
rect 13160 21490 13400 21510
rect 13490 21490 13730 21510
rect 13820 21490 14060 21510
rect 14190 21490 14430 21510
rect 14520 21490 14760 21510
rect 14850 21490 15090 21510
rect 15180 21490 15420 21510
rect 15510 21490 15750 21510
rect 15840 21490 16080 21510
rect 16170 21490 16410 21510
rect 16500 21490 16740 21510
rect 16830 21490 17070 21510
rect 17200 21490 17440 21510
rect 17530 21490 17770 21510
rect 17860 21490 18100 21510
rect 18190 21490 18430 21510
rect 18520 21490 18760 21510
rect 18850 21490 19090 21510
rect 19180 21490 19420 21510
rect 19510 21490 19750 21510
rect 19840 21490 20080 21510
rect 8170 21420 8180 21490
rect 8180 21420 8250 21490
rect 8250 21420 8270 21490
rect 8270 21420 8340 21490
rect 8340 21420 8360 21490
rect 8360 21420 8410 21490
rect 8500 21420 8520 21490
rect 8520 21420 8540 21490
rect 8540 21420 8610 21490
rect 8610 21420 8630 21490
rect 8630 21420 8700 21490
rect 8700 21420 8720 21490
rect 8720 21420 8740 21490
rect 8830 21420 8880 21490
rect 8880 21420 8900 21490
rect 8900 21420 8970 21490
rect 8970 21420 8990 21490
rect 8990 21420 9060 21490
rect 9060 21420 9070 21490
rect 9160 21420 9170 21490
rect 9170 21420 9240 21490
rect 9240 21420 9260 21490
rect 9260 21420 9330 21490
rect 9330 21420 9350 21490
rect 9350 21420 9400 21490
rect 9490 21420 9510 21490
rect 9510 21420 9530 21490
rect 9530 21420 9600 21490
rect 9600 21420 9620 21490
rect 9620 21420 9690 21490
rect 9690 21420 9710 21490
rect 9710 21420 9730 21490
rect 9820 21420 9870 21490
rect 9870 21420 9890 21490
rect 9890 21420 9960 21490
rect 9960 21420 9980 21490
rect 9980 21420 10050 21490
rect 10050 21420 10060 21490
rect 10150 21420 10160 21490
rect 10160 21420 10230 21490
rect 10230 21420 10250 21490
rect 10250 21420 10320 21490
rect 10320 21420 10340 21490
rect 10340 21420 10390 21490
rect 10480 21420 10500 21490
rect 10500 21420 10520 21490
rect 10520 21420 10590 21490
rect 10590 21420 10610 21490
rect 10610 21420 10680 21490
rect 10680 21420 10700 21490
rect 10700 21420 10720 21490
rect 10810 21420 10860 21490
rect 10860 21420 10880 21490
rect 10880 21420 10950 21490
rect 10950 21420 10970 21490
rect 10970 21420 11040 21490
rect 11040 21420 11050 21490
rect 11180 21420 11190 21490
rect 11190 21420 11260 21490
rect 11260 21420 11280 21490
rect 11280 21420 11350 21490
rect 11350 21420 11370 21490
rect 11370 21420 11420 21490
rect 11510 21420 11530 21490
rect 11530 21420 11550 21490
rect 11550 21420 11620 21490
rect 11620 21420 11640 21490
rect 11640 21420 11710 21490
rect 11710 21420 11730 21490
rect 11730 21420 11750 21490
rect 11840 21420 11890 21490
rect 11890 21420 11910 21490
rect 11910 21420 11980 21490
rect 11980 21420 12000 21490
rect 12000 21420 12070 21490
rect 12070 21420 12080 21490
rect 12170 21420 12180 21490
rect 12180 21420 12250 21490
rect 12250 21420 12270 21490
rect 12270 21420 12340 21490
rect 12340 21420 12360 21490
rect 12360 21420 12410 21490
rect 12500 21420 12520 21490
rect 12520 21420 12540 21490
rect 12540 21420 12610 21490
rect 12610 21420 12630 21490
rect 12630 21420 12700 21490
rect 12700 21420 12720 21490
rect 12720 21420 12740 21490
rect 12830 21420 12880 21490
rect 12880 21420 12900 21490
rect 12900 21420 12970 21490
rect 12970 21420 12990 21490
rect 12990 21420 13060 21490
rect 13060 21420 13070 21490
rect 13160 21420 13170 21490
rect 13170 21420 13240 21490
rect 13240 21420 13260 21490
rect 13260 21420 13330 21490
rect 13330 21420 13350 21490
rect 13350 21420 13400 21490
rect 13490 21420 13510 21490
rect 13510 21420 13530 21490
rect 13530 21420 13600 21490
rect 13600 21420 13620 21490
rect 13620 21420 13690 21490
rect 13690 21420 13710 21490
rect 13710 21420 13730 21490
rect 13820 21420 13870 21490
rect 13870 21420 13890 21490
rect 13890 21420 13960 21490
rect 13960 21420 13980 21490
rect 13980 21420 14050 21490
rect 14050 21420 14060 21490
rect 14190 21420 14200 21490
rect 14200 21420 14270 21490
rect 14270 21420 14290 21490
rect 14290 21420 14360 21490
rect 14360 21420 14380 21490
rect 14380 21420 14430 21490
rect 14520 21420 14540 21490
rect 14540 21420 14560 21490
rect 14560 21420 14630 21490
rect 14630 21420 14650 21490
rect 14650 21420 14720 21490
rect 14720 21420 14740 21490
rect 14740 21420 14760 21490
rect 14850 21420 14900 21490
rect 14900 21420 14920 21490
rect 14920 21420 14990 21490
rect 14990 21420 15010 21490
rect 15010 21420 15080 21490
rect 15080 21420 15090 21490
rect 15180 21420 15190 21490
rect 15190 21420 15260 21490
rect 15260 21420 15280 21490
rect 15280 21420 15350 21490
rect 15350 21420 15370 21490
rect 15370 21420 15420 21490
rect 15510 21420 15530 21490
rect 15530 21420 15550 21490
rect 15550 21420 15620 21490
rect 15620 21420 15640 21490
rect 15640 21420 15710 21490
rect 15710 21420 15730 21490
rect 15730 21420 15750 21490
rect 15840 21420 15890 21490
rect 15890 21420 15910 21490
rect 15910 21420 15980 21490
rect 15980 21420 16000 21490
rect 16000 21420 16070 21490
rect 16070 21420 16080 21490
rect 16170 21420 16180 21490
rect 16180 21420 16250 21490
rect 16250 21420 16270 21490
rect 16270 21420 16340 21490
rect 16340 21420 16360 21490
rect 16360 21420 16410 21490
rect 16500 21420 16520 21490
rect 16520 21420 16540 21490
rect 16540 21420 16610 21490
rect 16610 21420 16630 21490
rect 16630 21420 16700 21490
rect 16700 21420 16720 21490
rect 16720 21420 16740 21490
rect 16830 21420 16880 21490
rect 16880 21420 16900 21490
rect 16900 21420 16970 21490
rect 16970 21420 16990 21490
rect 16990 21420 17060 21490
rect 17060 21420 17070 21490
rect 17200 21420 17210 21490
rect 17210 21420 17280 21490
rect 17280 21420 17300 21490
rect 17300 21420 17370 21490
rect 17370 21420 17390 21490
rect 17390 21420 17440 21490
rect 17530 21420 17550 21490
rect 17550 21420 17570 21490
rect 17570 21420 17640 21490
rect 17640 21420 17660 21490
rect 17660 21420 17730 21490
rect 17730 21420 17750 21490
rect 17750 21420 17770 21490
rect 17860 21420 17910 21490
rect 17910 21420 17930 21490
rect 17930 21420 18000 21490
rect 18000 21420 18020 21490
rect 18020 21420 18090 21490
rect 18090 21420 18100 21490
rect 18190 21420 18200 21490
rect 18200 21420 18270 21490
rect 18270 21420 18290 21490
rect 18290 21420 18360 21490
rect 18360 21420 18380 21490
rect 18380 21420 18430 21490
rect 18520 21420 18540 21490
rect 18540 21420 18560 21490
rect 18560 21420 18630 21490
rect 18630 21420 18650 21490
rect 18650 21420 18720 21490
rect 18720 21420 18740 21490
rect 18740 21420 18760 21490
rect 18850 21420 18900 21490
rect 18900 21420 18920 21490
rect 18920 21420 18990 21490
rect 18990 21420 19010 21490
rect 19010 21420 19080 21490
rect 19080 21420 19090 21490
rect 19180 21420 19190 21490
rect 19190 21420 19260 21490
rect 19260 21420 19280 21490
rect 19280 21420 19350 21490
rect 19350 21420 19370 21490
rect 19370 21420 19420 21490
rect 19510 21420 19530 21490
rect 19530 21420 19550 21490
rect 19550 21420 19620 21490
rect 19620 21420 19640 21490
rect 19640 21420 19710 21490
rect 19710 21420 19730 21490
rect 19730 21420 19750 21490
rect 19840 21420 19890 21490
rect 19890 21420 19910 21490
rect 19910 21420 19980 21490
rect 19980 21420 20000 21490
rect 20000 21420 20070 21490
rect 20070 21420 20080 21490
rect 8170 21400 8410 21420
rect 8500 21400 8740 21420
rect 8830 21400 9070 21420
rect 9160 21400 9400 21420
rect 9490 21400 9730 21420
rect 9820 21400 10060 21420
rect 10150 21400 10390 21420
rect 10480 21400 10720 21420
rect 10810 21400 11050 21420
rect 11180 21400 11420 21420
rect 11510 21400 11750 21420
rect 11840 21400 12080 21420
rect 12170 21400 12410 21420
rect 12500 21400 12740 21420
rect 12830 21400 13070 21420
rect 13160 21400 13400 21420
rect 13490 21400 13730 21420
rect 13820 21400 14060 21420
rect 14190 21400 14430 21420
rect 14520 21400 14760 21420
rect 14850 21400 15090 21420
rect 15180 21400 15420 21420
rect 15510 21400 15750 21420
rect 15840 21400 16080 21420
rect 16170 21400 16410 21420
rect 16500 21400 16740 21420
rect 16830 21400 17070 21420
rect 17200 21400 17440 21420
rect 17530 21400 17770 21420
rect 17860 21400 18100 21420
rect 18190 21400 18430 21420
rect 18520 21400 18760 21420
rect 18850 21400 19090 21420
rect 19180 21400 19420 21420
rect 19510 21400 19750 21420
rect 19840 21400 20080 21420
rect 8170 21370 8180 21400
rect 8180 21370 8250 21400
rect 8250 21370 8270 21400
rect 8270 21370 8340 21400
rect 8340 21370 8360 21400
rect 8360 21370 8410 21400
rect 8500 21370 8520 21400
rect 8520 21370 8540 21400
rect 8540 21370 8610 21400
rect 8610 21370 8630 21400
rect 8630 21370 8700 21400
rect 8700 21370 8720 21400
rect 8720 21370 8740 21400
rect 8830 21370 8880 21400
rect 8880 21370 8900 21400
rect 8900 21370 8970 21400
rect 8970 21370 8990 21400
rect 8990 21370 9060 21400
rect 9060 21370 9070 21400
rect 9160 21370 9170 21400
rect 9170 21370 9240 21400
rect 9240 21370 9260 21400
rect 9260 21370 9330 21400
rect 9330 21370 9350 21400
rect 9350 21370 9400 21400
rect 9490 21370 9510 21400
rect 9510 21370 9530 21400
rect 9530 21370 9600 21400
rect 9600 21370 9620 21400
rect 9620 21370 9690 21400
rect 9690 21370 9710 21400
rect 9710 21370 9730 21400
rect 9820 21370 9870 21400
rect 9870 21370 9890 21400
rect 9890 21370 9960 21400
rect 9960 21370 9980 21400
rect 9980 21370 10050 21400
rect 10050 21370 10060 21400
rect 10150 21370 10160 21400
rect 10160 21370 10230 21400
rect 10230 21370 10250 21400
rect 10250 21370 10320 21400
rect 10320 21370 10340 21400
rect 10340 21370 10390 21400
rect 10480 21370 10500 21400
rect 10500 21370 10520 21400
rect 10520 21370 10590 21400
rect 10590 21370 10610 21400
rect 10610 21370 10680 21400
rect 10680 21370 10700 21400
rect 10700 21370 10720 21400
rect 10810 21370 10860 21400
rect 10860 21370 10880 21400
rect 10880 21370 10950 21400
rect 10950 21370 10970 21400
rect 10970 21370 11040 21400
rect 11040 21370 11050 21400
rect 11180 21370 11190 21400
rect 11190 21370 11260 21400
rect 11260 21370 11280 21400
rect 11280 21370 11350 21400
rect 11350 21370 11370 21400
rect 11370 21370 11420 21400
rect 11510 21370 11530 21400
rect 11530 21370 11550 21400
rect 11550 21370 11620 21400
rect 11620 21370 11640 21400
rect 11640 21370 11710 21400
rect 11710 21370 11730 21400
rect 11730 21370 11750 21400
rect 11840 21370 11890 21400
rect 11890 21370 11910 21400
rect 11910 21370 11980 21400
rect 11980 21370 12000 21400
rect 12000 21370 12070 21400
rect 12070 21370 12080 21400
rect 12170 21370 12180 21400
rect 12180 21370 12250 21400
rect 12250 21370 12270 21400
rect 12270 21370 12340 21400
rect 12340 21370 12360 21400
rect 12360 21370 12410 21400
rect 12500 21370 12520 21400
rect 12520 21370 12540 21400
rect 12540 21370 12610 21400
rect 12610 21370 12630 21400
rect 12630 21370 12700 21400
rect 12700 21370 12720 21400
rect 12720 21370 12740 21400
rect 12830 21370 12880 21400
rect 12880 21370 12900 21400
rect 12900 21370 12970 21400
rect 12970 21370 12990 21400
rect 12990 21370 13060 21400
rect 13060 21370 13070 21400
rect 13160 21370 13170 21400
rect 13170 21370 13240 21400
rect 13240 21370 13260 21400
rect 13260 21370 13330 21400
rect 13330 21370 13350 21400
rect 13350 21370 13400 21400
rect 13490 21370 13510 21400
rect 13510 21370 13530 21400
rect 13530 21370 13600 21400
rect 13600 21370 13620 21400
rect 13620 21370 13690 21400
rect 13690 21370 13710 21400
rect 13710 21370 13730 21400
rect 13820 21370 13870 21400
rect 13870 21370 13890 21400
rect 13890 21370 13960 21400
rect 13960 21370 13980 21400
rect 13980 21370 14050 21400
rect 14050 21370 14060 21400
rect 14190 21370 14200 21400
rect 14200 21370 14270 21400
rect 14270 21370 14290 21400
rect 14290 21370 14360 21400
rect 14360 21370 14380 21400
rect 14380 21370 14430 21400
rect 14520 21370 14540 21400
rect 14540 21370 14560 21400
rect 14560 21370 14630 21400
rect 14630 21370 14650 21400
rect 14650 21370 14720 21400
rect 14720 21370 14740 21400
rect 14740 21370 14760 21400
rect 14850 21370 14900 21400
rect 14900 21370 14920 21400
rect 14920 21370 14990 21400
rect 14990 21370 15010 21400
rect 15010 21370 15080 21400
rect 15080 21370 15090 21400
rect 15180 21370 15190 21400
rect 15190 21370 15260 21400
rect 15260 21370 15280 21400
rect 15280 21370 15350 21400
rect 15350 21370 15370 21400
rect 15370 21370 15420 21400
rect 15510 21370 15530 21400
rect 15530 21370 15550 21400
rect 15550 21370 15620 21400
rect 15620 21370 15640 21400
rect 15640 21370 15710 21400
rect 15710 21370 15730 21400
rect 15730 21370 15750 21400
rect 15840 21370 15890 21400
rect 15890 21370 15910 21400
rect 15910 21370 15980 21400
rect 15980 21370 16000 21400
rect 16000 21370 16070 21400
rect 16070 21370 16080 21400
rect 16170 21370 16180 21400
rect 16180 21370 16250 21400
rect 16250 21370 16270 21400
rect 16270 21370 16340 21400
rect 16340 21370 16360 21400
rect 16360 21370 16410 21400
rect 16500 21370 16520 21400
rect 16520 21370 16540 21400
rect 16540 21370 16610 21400
rect 16610 21370 16630 21400
rect 16630 21370 16700 21400
rect 16700 21370 16720 21400
rect 16720 21370 16740 21400
rect 16830 21370 16880 21400
rect 16880 21370 16900 21400
rect 16900 21370 16970 21400
rect 16970 21370 16990 21400
rect 16990 21370 17060 21400
rect 17060 21370 17070 21400
rect 17200 21370 17210 21400
rect 17210 21370 17280 21400
rect 17280 21370 17300 21400
rect 17300 21370 17370 21400
rect 17370 21370 17390 21400
rect 17390 21370 17440 21400
rect 17530 21370 17550 21400
rect 17550 21370 17570 21400
rect 17570 21370 17640 21400
rect 17640 21370 17660 21400
rect 17660 21370 17730 21400
rect 17730 21370 17750 21400
rect 17750 21370 17770 21400
rect 17860 21370 17910 21400
rect 17910 21370 17930 21400
rect 17930 21370 18000 21400
rect 18000 21370 18020 21400
rect 18020 21370 18090 21400
rect 18090 21370 18100 21400
rect 18190 21370 18200 21400
rect 18200 21370 18270 21400
rect 18270 21370 18290 21400
rect 18290 21370 18360 21400
rect 18360 21370 18380 21400
rect 18380 21370 18430 21400
rect 18520 21370 18540 21400
rect 18540 21370 18560 21400
rect 18560 21370 18630 21400
rect 18630 21370 18650 21400
rect 18650 21370 18720 21400
rect 18720 21370 18740 21400
rect 18740 21370 18760 21400
rect 18850 21370 18900 21400
rect 18900 21370 18920 21400
rect 18920 21370 18990 21400
rect 18990 21370 19010 21400
rect 19010 21370 19080 21400
rect 19080 21370 19090 21400
rect 19180 21370 19190 21400
rect 19190 21370 19260 21400
rect 19260 21370 19280 21400
rect 19280 21370 19350 21400
rect 19350 21370 19370 21400
rect 19370 21370 19420 21400
rect 19510 21370 19530 21400
rect 19530 21370 19550 21400
rect 19550 21370 19620 21400
rect 19620 21370 19640 21400
rect 19640 21370 19710 21400
rect 19710 21370 19730 21400
rect 19730 21370 19750 21400
rect 19840 21370 19890 21400
rect 19890 21370 19910 21400
rect 19910 21370 19980 21400
rect 19980 21370 20000 21400
rect 20000 21370 20070 21400
rect 20070 21370 20080 21400
rect 1720 6850 1960 6910
rect 2050 6850 2290 6910
rect 2390 6850 2630 6910
rect 2720 6850 2960 6910
rect 1720 6780 1750 6850
rect 1750 6780 1790 6850
rect 1790 6780 1860 6850
rect 1860 6780 1900 6850
rect 1900 6780 1960 6850
rect 2050 6780 2080 6850
rect 2080 6780 2120 6850
rect 2120 6780 2190 6850
rect 2190 6780 2230 6850
rect 2230 6780 2290 6850
rect 2390 6780 2410 6850
rect 2410 6780 2450 6850
rect 2450 6780 2520 6850
rect 2520 6780 2560 6850
rect 2560 6780 2630 6850
rect 2720 6780 2740 6850
rect 2740 6780 2780 6850
rect 2780 6780 2850 6850
rect 2850 6780 2890 6850
rect 2890 6780 2960 6850
rect 1720 6740 1960 6780
rect 2050 6740 2290 6780
rect 2390 6740 2630 6780
rect 2720 6740 2960 6780
rect 1720 6670 1750 6740
rect 1750 6670 1790 6740
rect 1790 6670 1860 6740
rect 1860 6670 1900 6740
rect 1900 6670 1960 6740
rect 2050 6670 2080 6740
rect 2080 6670 2120 6740
rect 2120 6670 2190 6740
rect 2190 6670 2230 6740
rect 2230 6670 2290 6740
rect 2390 6670 2410 6740
rect 2410 6670 2450 6740
rect 2450 6670 2520 6740
rect 2520 6670 2560 6740
rect 2560 6670 2630 6740
rect 2720 6670 2740 6740
rect 2740 6670 2780 6740
rect 2780 6670 2850 6740
rect 2850 6670 2890 6740
rect 2890 6670 2960 6740
rect 11940 6880 12180 6940
rect 12270 6880 12510 6940
rect 12610 6880 12850 6940
rect 12940 6880 13180 6940
rect 11940 6810 11970 6880
rect 11970 6810 12010 6880
rect 12010 6810 12080 6880
rect 12080 6810 12120 6880
rect 12120 6810 12180 6880
rect 12270 6810 12300 6880
rect 12300 6810 12340 6880
rect 12340 6810 12410 6880
rect 12410 6810 12450 6880
rect 12450 6810 12510 6880
rect 12610 6810 12630 6880
rect 12630 6810 12670 6880
rect 12670 6810 12740 6880
rect 12740 6810 12780 6880
rect 12780 6810 12850 6880
rect 12940 6810 12960 6880
rect 12960 6810 13000 6880
rect 13000 6810 13070 6880
rect 13070 6810 13110 6880
rect 13110 6810 13180 6880
rect 11940 6770 12180 6810
rect 12270 6770 12510 6810
rect 12610 6770 12850 6810
rect 12940 6770 13180 6810
rect 11940 6700 11970 6770
rect 11970 6700 12010 6770
rect 12010 6700 12080 6770
rect 12080 6700 12120 6770
rect 12120 6700 12180 6770
rect 12270 6700 12300 6770
rect 12300 6700 12340 6770
rect 12340 6700 12410 6770
rect 12410 6700 12450 6770
rect 12450 6700 12510 6770
rect 12610 6700 12630 6770
rect 12630 6700 12670 6770
rect 12670 6700 12740 6770
rect 12740 6700 12780 6770
rect 12780 6700 12850 6770
rect 12940 6700 12960 6770
rect 12960 6700 13000 6770
rect 13000 6700 13070 6770
rect 13070 6700 13110 6770
rect 13110 6700 13180 6770
rect 23510 7210 23880 7270
rect 23510 7140 23560 7210
rect 23560 7140 23600 7210
rect 23600 7140 23670 7210
rect 23670 7140 23710 7210
rect 23710 7140 23780 7210
rect 23780 7140 23820 7210
rect 23820 7140 23880 7210
rect 23510 7100 23880 7140
rect 23510 7030 23560 7100
rect 23560 7030 23600 7100
rect 23600 7030 23670 7100
rect 23670 7030 23710 7100
rect 23710 7030 23780 7100
rect 23780 7030 23820 7100
rect 23820 7030 23880 7100
rect 25910 7210 26280 7270
rect 25910 7140 25960 7210
rect 25960 7140 26000 7210
rect 26000 7140 26070 7210
rect 26070 7140 26110 7210
rect 26110 7140 26180 7210
rect 26180 7140 26220 7210
rect 26220 7140 26280 7210
rect 25910 7100 26280 7140
rect 25910 7030 25960 7100
rect 25960 7030 26000 7100
rect 26000 7030 26070 7100
rect 26070 7030 26110 7100
rect 26110 7030 26180 7100
rect 26180 7030 26220 7100
rect 26220 7030 26280 7100
rect 1260 -860 1330 -790
rect 1330 -860 1370 -790
rect 1370 -860 1440 -790
rect 1440 -860 1480 -790
rect 1480 -860 1500 -790
rect 1590 -860 1660 -790
rect 1660 -860 1700 -790
rect 1700 -860 1770 -790
rect 1770 -860 1810 -790
rect 1810 -860 1830 -790
rect 1930 -860 1990 -790
rect 1990 -860 2030 -790
rect 2030 -860 2100 -790
rect 2100 -860 2140 -790
rect 2140 -860 2170 -790
rect 2260 -860 2320 -790
rect 2320 -860 2360 -790
rect 2360 -860 2430 -790
rect 2430 -860 2470 -790
rect 2470 -860 2500 -790
rect 1260 -900 1500 -860
rect 1590 -900 1830 -860
rect 1930 -900 2170 -860
rect 2260 -900 2500 -860
rect 1260 -970 1330 -900
rect 1330 -970 1370 -900
rect 1370 -970 1440 -900
rect 1440 -970 1480 -900
rect 1480 -970 1500 -900
rect 1590 -970 1660 -900
rect 1660 -970 1700 -900
rect 1700 -970 1770 -900
rect 1770 -970 1810 -900
rect 1810 -970 1830 -900
rect 1930 -970 1990 -900
rect 1990 -970 2030 -900
rect 2030 -970 2100 -900
rect 2100 -970 2140 -900
rect 2140 -970 2170 -900
rect 2260 -970 2320 -900
rect 2320 -970 2360 -900
rect 2360 -970 2430 -900
rect 2430 -970 2470 -900
rect 2470 -970 2500 -900
rect 1260 -1030 1500 -970
rect 1590 -1030 1830 -970
rect 1930 -1030 2170 -970
rect 2260 -1030 2500 -970
rect 12400 -860 12430 -790
rect 12430 -860 12470 -790
rect 12470 -860 12540 -790
rect 12540 -860 12580 -790
rect 12580 -860 12640 -790
rect 12730 -860 12760 -790
rect 12760 -860 12800 -790
rect 12800 -860 12870 -790
rect 12870 -860 12910 -790
rect 12910 -860 12970 -790
rect 13070 -860 13090 -790
rect 13090 -860 13130 -790
rect 13130 -860 13200 -790
rect 13200 -860 13240 -790
rect 13240 -860 13310 -790
rect 13400 -860 13420 -790
rect 13420 -860 13460 -790
rect 13460 -860 13530 -790
rect 13530 -860 13570 -790
rect 13570 -860 13640 -790
rect 12400 -900 12640 -860
rect 12730 -900 12970 -860
rect 13070 -900 13310 -860
rect 13400 -900 13640 -860
rect 12400 -970 12430 -900
rect 12430 -970 12470 -900
rect 12470 -970 12540 -900
rect 12540 -970 12580 -900
rect 12580 -970 12640 -900
rect 12730 -970 12760 -900
rect 12760 -970 12800 -900
rect 12800 -970 12870 -900
rect 12870 -970 12910 -900
rect 12910 -970 12970 -900
rect 13070 -970 13090 -900
rect 13090 -970 13130 -900
rect 13130 -970 13200 -900
rect 13200 -970 13240 -900
rect 13240 -970 13310 -900
rect 13400 -970 13420 -900
rect 13420 -970 13460 -900
rect 13460 -970 13530 -900
rect 13530 -970 13570 -900
rect 13570 -970 13640 -900
rect 12400 -1030 12640 -970
rect 12730 -1030 12970 -970
rect 13070 -1030 13310 -970
rect 13400 -1030 13640 -970
rect 1720 -2780 1960 -2720
rect 2050 -2780 2290 -2720
rect 2390 -2780 2630 -2720
rect 2720 -2780 2960 -2720
rect 1720 -2850 1750 -2780
rect 1750 -2850 1790 -2780
rect 1790 -2850 1860 -2780
rect 1860 -2850 1900 -2780
rect 1900 -2850 1960 -2780
rect 2050 -2850 2080 -2780
rect 2080 -2850 2120 -2780
rect 2120 -2850 2190 -2780
rect 2190 -2850 2230 -2780
rect 2230 -2850 2290 -2780
rect 2390 -2850 2410 -2780
rect 2410 -2850 2450 -2780
rect 2450 -2850 2520 -2780
rect 2520 -2850 2560 -2780
rect 2560 -2850 2630 -2780
rect 2720 -2850 2740 -2780
rect 2740 -2850 2780 -2780
rect 2780 -2850 2850 -2780
rect 2850 -2850 2890 -2780
rect 2890 -2850 2960 -2780
rect 1720 -2890 1960 -2850
rect 2050 -2890 2290 -2850
rect 2390 -2890 2630 -2850
rect 2720 -2890 2960 -2850
rect 1720 -2960 1750 -2890
rect 1750 -2960 1790 -2890
rect 1790 -2960 1860 -2890
rect 1860 -2960 1900 -2890
rect 1900 -2960 1960 -2890
rect 2050 -2960 2080 -2890
rect 2080 -2960 2120 -2890
rect 2120 -2960 2190 -2890
rect 2190 -2960 2230 -2890
rect 2230 -2960 2290 -2890
rect 2390 -2960 2410 -2890
rect 2410 -2960 2450 -2890
rect 2450 -2960 2520 -2890
rect 2520 -2960 2560 -2890
rect 2560 -2960 2630 -2890
rect 2720 -2960 2740 -2890
rect 2740 -2960 2780 -2890
rect 2780 -2960 2850 -2890
rect 2850 -2960 2890 -2890
rect 2890 -2960 2960 -2890
rect 11940 -2780 12180 -2720
rect 12270 -2780 12510 -2720
rect 12610 -2780 12850 -2720
rect 12940 -2780 13180 -2720
rect 11940 -2850 11970 -2780
rect 11970 -2850 12010 -2780
rect 12010 -2850 12080 -2780
rect 12080 -2850 12120 -2780
rect 12120 -2850 12180 -2780
rect 12270 -2850 12300 -2780
rect 12300 -2850 12340 -2780
rect 12340 -2850 12410 -2780
rect 12410 -2850 12450 -2780
rect 12450 -2850 12510 -2780
rect 12610 -2850 12630 -2780
rect 12630 -2850 12670 -2780
rect 12670 -2850 12740 -2780
rect 12740 -2850 12780 -2780
rect 12780 -2850 12850 -2780
rect 12940 -2850 12960 -2780
rect 12960 -2850 13000 -2780
rect 13000 -2850 13070 -2780
rect 13070 -2850 13110 -2780
rect 13110 -2850 13180 -2780
rect 11940 -2890 12180 -2850
rect 12270 -2890 12510 -2850
rect 12610 -2890 12850 -2850
rect 12940 -2890 13180 -2850
rect 11940 -2960 11970 -2890
rect 11970 -2960 12010 -2890
rect 12010 -2960 12080 -2890
rect 12080 -2960 12120 -2890
rect 12120 -2960 12180 -2890
rect 12270 -2960 12300 -2890
rect 12300 -2960 12340 -2890
rect 12340 -2960 12410 -2890
rect 12410 -2960 12450 -2890
rect 12450 -2960 12510 -2890
rect 12610 -2960 12630 -2890
rect 12630 -2960 12670 -2890
rect 12670 -2960 12740 -2890
rect 12740 -2960 12780 -2890
rect 12780 -2960 12850 -2890
rect 12940 -2960 12960 -2890
rect 12960 -2960 13000 -2890
rect 13000 -2960 13070 -2890
rect 13070 -2960 13110 -2890
rect 13110 -2960 13180 -2890
rect 22480 2530 22540 2600
rect 22540 2530 22580 2600
rect 22580 2530 22650 2600
rect 22650 2530 22690 2600
rect 22690 2530 22760 2600
rect 22760 2530 22800 2600
rect 22800 2530 22850 2600
rect 22480 2490 22850 2530
rect 22480 2420 22540 2490
rect 22540 2420 22580 2490
rect 22580 2420 22650 2490
rect 22650 2420 22690 2490
rect 22690 2420 22760 2490
rect 22760 2420 22800 2490
rect 22800 2420 22850 2490
rect 22480 2360 22850 2420
rect 26960 2530 27020 2600
rect 27020 2530 27060 2600
rect 27060 2530 27130 2600
rect 27130 2530 27170 2600
rect 27170 2530 27240 2600
rect 27240 2530 27280 2600
rect 27280 2530 27330 2600
rect 26960 2490 27330 2530
rect 26960 2420 27020 2490
rect 27020 2420 27060 2490
rect 27060 2420 27130 2490
rect 27130 2420 27170 2490
rect 27170 2420 27240 2490
rect 27240 2420 27280 2490
rect 27280 2420 27330 2490
rect 26960 2360 27330 2420
rect 23510 920 23880 980
rect 23510 850 23560 920
rect 23560 850 23600 920
rect 23600 850 23670 920
rect 23670 850 23710 920
rect 23710 850 23780 920
rect 23780 850 23820 920
rect 23820 850 23880 920
rect 23510 810 23880 850
rect 23510 740 23560 810
rect 23560 740 23600 810
rect 23600 740 23670 810
rect 23670 740 23710 810
rect 23710 740 23780 810
rect 23780 740 23820 810
rect 23820 740 23880 810
rect 25910 920 26280 980
rect 25910 850 25960 920
rect 25960 850 26000 920
rect 26000 850 26070 920
rect 26070 850 26110 920
rect 26110 850 26180 920
rect 26180 850 26220 920
rect 26220 850 26280 920
rect 25910 810 26280 850
rect 25910 740 25960 810
rect 25960 740 26000 810
rect 26000 740 26070 810
rect 26070 740 26110 810
rect 26110 740 26180 810
rect 26180 740 26220 810
rect 26220 740 26280 810
rect 38230 7750 38260 7770
rect 38260 7750 38280 7770
rect 38280 7750 38350 7770
rect 38350 7750 38370 7770
rect 38370 7750 38440 7770
rect 38440 7750 38470 7770
rect 38230 7730 38470 7750
rect 38230 7660 38260 7730
rect 38260 7660 38280 7730
rect 38280 7660 38350 7730
rect 38350 7660 38370 7730
rect 38370 7660 38440 7730
rect 38440 7660 38470 7730
rect 38230 7640 38470 7660
rect 38230 7570 38260 7640
rect 38260 7570 38280 7640
rect 38280 7570 38350 7640
rect 38350 7570 38370 7640
rect 38370 7570 38440 7640
rect 38440 7570 38470 7640
rect 38230 7550 38470 7570
rect 38230 7530 38260 7550
rect 38260 7530 38280 7550
rect 38280 7530 38350 7550
rect 38350 7530 38370 7550
rect 38370 7530 38440 7550
rect 38440 7530 38470 7550
rect 38230 7390 38260 7440
rect 38260 7390 38280 7440
rect 38280 7390 38350 7440
rect 38350 7390 38370 7440
rect 38370 7390 38440 7440
rect 38440 7390 38470 7440
rect 38230 7370 38470 7390
rect 38230 7300 38260 7370
rect 38260 7300 38280 7370
rect 38280 7300 38350 7370
rect 38350 7300 38370 7370
rect 38370 7300 38440 7370
rect 38440 7300 38470 7370
rect 38230 7280 38470 7300
rect 38230 7210 38260 7280
rect 38260 7210 38280 7280
rect 38280 7210 38350 7280
rect 38350 7210 38370 7280
rect 38370 7210 38440 7280
rect 38440 7210 38470 7280
rect 38230 7200 38470 7210
rect 38230 7060 38470 7070
rect 38230 6990 38260 7060
rect 38260 6990 38280 7060
rect 38280 6990 38350 7060
rect 38350 6990 38370 7060
rect 38370 6990 38440 7060
rect 38440 6990 38470 7060
rect 38230 6970 38470 6990
rect 38230 6900 38260 6970
rect 38260 6900 38280 6970
rect 38280 6900 38350 6970
rect 38350 6900 38370 6970
rect 38370 6900 38440 6970
rect 38440 6900 38470 6970
rect 38230 6880 38470 6900
rect 38230 6830 38260 6880
rect 38260 6830 38280 6880
rect 38280 6830 38350 6880
rect 38350 6830 38370 6880
rect 38370 6830 38440 6880
rect 38440 6830 38470 6880
rect 38230 6720 38260 6740
rect 38260 6720 38280 6740
rect 38280 6720 38350 6740
rect 38350 6720 38370 6740
rect 38370 6720 38440 6740
rect 38440 6720 38470 6740
rect 38230 6700 38470 6720
rect 38230 6630 38260 6700
rect 38260 6630 38280 6700
rect 38280 6630 38350 6700
rect 38350 6630 38370 6700
rect 38370 6630 38440 6700
rect 38440 6630 38470 6700
rect 38230 6610 38470 6630
rect 38230 6540 38260 6610
rect 38260 6540 38280 6610
rect 38280 6540 38350 6610
rect 38350 6540 38370 6610
rect 38370 6540 38440 6610
rect 38440 6540 38470 6610
rect 38230 6520 38470 6540
rect 38230 6500 38260 6520
rect 38260 6500 38280 6520
rect 38280 6500 38350 6520
rect 38350 6500 38370 6520
rect 38370 6500 38440 6520
rect 38440 6500 38470 6520
rect 38230 6360 38260 6410
rect 38260 6360 38280 6410
rect 38280 6360 38350 6410
rect 38350 6360 38370 6410
rect 38370 6360 38440 6410
rect 38440 6360 38470 6410
rect 38230 6340 38470 6360
rect 38230 6270 38260 6340
rect 38260 6270 38280 6340
rect 38280 6270 38350 6340
rect 38350 6270 38370 6340
rect 38370 6270 38440 6340
rect 38440 6270 38470 6340
rect 38230 6250 38470 6270
rect 38230 6180 38260 6250
rect 38260 6180 38280 6250
rect 38280 6180 38350 6250
rect 38350 6180 38370 6250
rect 38370 6180 38440 6250
rect 38440 6180 38470 6250
rect 38230 6170 38470 6180
rect 38230 6070 38470 6080
rect 38230 6000 38260 6070
rect 38260 6000 38280 6070
rect 38280 6000 38350 6070
rect 38350 6000 38370 6070
rect 38370 6000 38440 6070
rect 38440 6000 38470 6070
rect 38230 5980 38470 6000
rect 38230 5910 38260 5980
rect 38260 5910 38280 5980
rect 38280 5910 38350 5980
rect 38350 5910 38370 5980
rect 38370 5910 38440 5980
rect 38440 5910 38470 5980
rect 38230 5890 38470 5910
rect 38230 5840 38260 5890
rect 38260 5840 38280 5890
rect 38280 5840 38350 5890
rect 38350 5840 38370 5890
rect 38370 5840 38440 5890
rect 38440 5840 38470 5890
rect 38230 5730 38260 5750
rect 38260 5730 38280 5750
rect 38280 5730 38350 5750
rect 38350 5730 38370 5750
rect 38370 5730 38440 5750
rect 38440 5730 38470 5750
rect 38230 5710 38470 5730
rect 38230 5640 38260 5710
rect 38260 5640 38280 5710
rect 38280 5640 38350 5710
rect 38350 5640 38370 5710
rect 38370 5640 38440 5710
rect 38440 5640 38470 5710
rect 38230 5620 38470 5640
rect 38230 5550 38260 5620
rect 38260 5550 38280 5620
rect 38280 5550 38350 5620
rect 38350 5550 38370 5620
rect 38370 5550 38440 5620
rect 38440 5550 38470 5620
rect 38230 5530 38470 5550
rect 38230 5510 38260 5530
rect 38260 5510 38280 5530
rect 38280 5510 38350 5530
rect 38350 5510 38370 5530
rect 38370 5510 38440 5530
rect 38440 5510 38470 5530
rect 38230 5370 38260 5420
rect 38260 5370 38280 5420
rect 38280 5370 38350 5420
rect 38350 5370 38370 5420
rect 38370 5370 38440 5420
rect 38440 5370 38470 5420
rect 38230 5350 38470 5370
rect 38230 5280 38260 5350
rect 38260 5280 38280 5350
rect 38280 5280 38350 5350
rect 38350 5280 38370 5350
rect 38370 5280 38440 5350
rect 38440 5280 38470 5350
rect 38230 5260 38470 5280
rect 38230 5190 38260 5260
rect 38260 5190 38280 5260
rect 38280 5190 38350 5260
rect 38350 5190 38370 5260
rect 38370 5190 38440 5260
rect 38440 5190 38470 5260
rect 38230 5180 38470 5190
rect 38230 5080 38470 5090
rect 38230 5010 38260 5080
rect 38260 5010 38280 5080
rect 38280 5010 38350 5080
rect 38350 5010 38370 5080
rect 38370 5010 38440 5080
rect 38440 5010 38470 5080
rect 38230 4990 38470 5010
rect 38230 4920 38260 4990
rect 38260 4920 38280 4990
rect 38280 4920 38350 4990
rect 38350 4920 38370 4990
rect 38370 4920 38440 4990
rect 38440 4920 38470 4990
rect 38230 4900 38470 4920
rect 38230 4850 38260 4900
rect 38260 4850 38280 4900
rect 38280 4850 38350 4900
rect 38350 4850 38370 4900
rect 38370 4850 38440 4900
rect 38440 4850 38470 4900
rect 38230 4740 38260 4760
rect 38260 4740 38280 4760
rect 38280 4740 38350 4760
rect 38350 4740 38370 4760
rect 38370 4740 38440 4760
rect 38440 4740 38470 4760
rect 38230 4720 38470 4740
rect 38230 4650 38260 4720
rect 38260 4650 38280 4720
rect 38280 4650 38350 4720
rect 38350 4650 38370 4720
rect 38370 4650 38440 4720
rect 38440 4650 38470 4720
rect 38230 4630 38470 4650
rect 38230 4560 38260 4630
rect 38260 4560 38280 4630
rect 38280 4560 38350 4630
rect 38350 4560 38370 4630
rect 38370 4560 38440 4630
rect 38440 4560 38470 4630
rect 38230 4540 38470 4560
rect 38230 4520 38260 4540
rect 38260 4520 38280 4540
rect 38280 4520 38350 4540
rect 38350 4520 38370 4540
rect 38370 4520 38440 4540
rect 38440 4520 38470 4540
rect 38230 4380 38260 4430
rect 38260 4380 38280 4430
rect 38280 4380 38350 4430
rect 38350 4380 38370 4430
rect 38370 4380 38440 4430
rect 38440 4380 38470 4430
rect 38230 4360 38470 4380
rect 38230 4290 38260 4360
rect 38260 4290 38280 4360
rect 38280 4290 38350 4360
rect 38350 4290 38370 4360
rect 38370 4290 38440 4360
rect 38440 4290 38470 4360
rect 38230 4270 38470 4290
rect 38230 4200 38260 4270
rect 38260 4200 38280 4270
rect 38280 4200 38350 4270
rect 38350 4200 38370 4270
rect 38370 4200 38440 4270
rect 38440 4200 38470 4270
rect 38230 4190 38470 4200
rect 38230 4050 38470 4060
rect 38230 3980 38260 4050
rect 38260 3980 38280 4050
rect 38280 3980 38350 4050
rect 38350 3980 38370 4050
rect 38370 3980 38440 4050
rect 38440 3980 38470 4050
rect 38230 3960 38470 3980
rect 38230 3890 38260 3960
rect 38260 3890 38280 3960
rect 38280 3890 38350 3960
rect 38350 3890 38370 3960
rect 38370 3890 38440 3960
rect 38440 3890 38470 3960
rect 38230 3870 38470 3890
rect 38230 3820 38260 3870
rect 38260 3820 38280 3870
rect 38280 3820 38350 3870
rect 38350 3820 38370 3870
rect 38370 3820 38440 3870
rect 38440 3820 38470 3870
rect 38230 3710 38260 3730
rect 38260 3710 38280 3730
rect 38280 3710 38350 3730
rect 38350 3710 38370 3730
rect 38370 3710 38440 3730
rect 38440 3710 38470 3730
rect 38230 3690 38470 3710
rect 38230 3620 38260 3690
rect 38260 3620 38280 3690
rect 38280 3620 38350 3690
rect 38350 3620 38370 3690
rect 38370 3620 38440 3690
rect 38440 3620 38470 3690
rect 38230 3600 38470 3620
rect 38230 3530 38260 3600
rect 38260 3530 38280 3600
rect 38280 3530 38350 3600
rect 38350 3530 38370 3600
rect 38370 3530 38440 3600
rect 38440 3530 38470 3600
rect 38230 3510 38470 3530
rect 38230 3490 38260 3510
rect 38260 3490 38280 3510
rect 38280 3490 38350 3510
rect 38350 3490 38370 3510
rect 38370 3490 38440 3510
rect 38440 3490 38470 3510
rect 38230 3350 38260 3400
rect 38260 3350 38280 3400
rect 38280 3350 38350 3400
rect 38350 3350 38370 3400
rect 38370 3350 38440 3400
rect 38440 3350 38470 3400
rect 38230 3330 38470 3350
rect 38230 3260 38260 3330
rect 38260 3260 38280 3330
rect 38280 3260 38350 3330
rect 38350 3260 38370 3330
rect 38370 3260 38440 3330
rect 38440 3260 38470 3330
rect 38230 3240 38470 3260
rect 38230 3170 38260 3240
rect 38260 3170 38280 3240
rect 38280 3170 38350 3240
rect 38350 3170 38370 3240
rect 38370 3170 38440 3240
rect 38440 3170 38470 3240
rect 38230 3160 38470 3170
rect 38230 3060 38470 3070
rect 38230 2990 38260 3060
rect 38260 2990 38280 3060
rect 38280 2990 38350 3060
rect 38350 2990 38370 3060
rect 38370 2990 38440 3060
rect 38440 2990 38470 3060
rect 38230 2970 38470 2990
rect 38230 2900 38260 2970
rect 38260 2900 38280 2970
rect 38280 2900 38350 2970
rect 38350 2900 38370 2970
rect 38370 2900 38440 2970
rect 38440 2900 38470 2970
rect 38230 2880 38470 2900
rect 38230 2830 38260 2880
rect 38260 2830 38280 2880
rect 38280 2830 38350 2880
rect 38350 2830 38370 2880
rect 38370 2830 38440 2880
rect 38440 2830 38470 2880
rect 38230 2720 38260 2740
rect 38260 2720 38280 2740
rect 38280 2720 38350 2740
rect 38350 2720 38370 2740
rect 38370 2720 38440 2740
rect 38440 2720 38470 2740
rect 38230 2700 38470 2720
rect 38230 2630 38260 2700
rect 38260 2630 38280 2700
rect 38280 2630 38350 2700
rect 38350 2630 38370 2700
rect 38370 2630 38440 2700
rect 38440 2630 38470 2700
rect 38230 2610 38470 2630
rect 38230 2540 38260 2610
rect 38260 2540 38280 2610
rect 38280 2540 38350 2610
rect 38350 2540 38370 2610
rect 38370 2540 38440 2610
rect 38440 2540 38470 2610
rect 38230 2520 38470 2540
rect 38230 2500 38260 2520
rect 38260 2500 38280 2520
rect 38280 2500 38350 2520
rect 38350 2500 38370 2520
rect 38370 2500 38440 2520
rect 38440 2500 38470 2520
rect 38230 2360 38260 2410
rect 38260 2360 38280 2410
rect 38280 2360 38350 2410
rect 38350 2360 38370 2410
rect 38370 2360 38440 2410
rect 38440 2360 38470 2410
rect 38230 2340 38470 2360
rect 38230 2270 38260 2340
rect 38260 2270 38280 2340
rect 38280 2270 38350 2340
rect 38350 2270 38370 2340
rect 38370 2270 38440 2340
rect 38440 2270 38470 2340
rect 38230 2250 38470 2270
rect 38230 2180 38260 2250
rect 38260 2180 38280 2250
rect 38280 2180 38350 2250
rect 38350 2180 38370 2250
rect 38370 2180 38440 2250
rect 38440 2180 38470 2250
rect 38230 2170 38470 2180
rect 38230 2070 38470 2080
rect 38230 2000 38260 2070
rect 38260 2000 38280 2070
rect 38280 2000 38350 2070
rect 38350 2000 38370 2070
rect 38370 2000 38440 2070
rect 38440 2000 38470 2070
rect 38230 1980 38470 2000
rect 38230 1910 38260 1980
rect 38260 1910 38280 1980
rect 38280 1910 38350 1980
rect 38350 1910 38370 1980
rect 38370 1910 38440 1980
rect 38440 1910 38470 1980
rect 38230 1890 38470 1910
rect 38230 1840 38260 1890
rect 38260 1840 38280 1890
rect 38280 1840 38350 1890
rect 38350 1840 38370 1890
rect 38370 1840 38440 1890
rect 38440 1840 38470 1890
rect 38230 1730 38260 1750
rect 38260 1730 38280 1750
rect 38280 1730 38350 1750
rect 38350 1730 38370 1750
rect 38370 1730 38440 1750
rect 38440 1730 38470 1750
rect 38230 1710 38470 1730
rect 38230 1640 38260 1710
rect 38260 1640 38280 1710
rect 38280 1640 38350 1710
rect 38350 1640 38370 1710
rect 38370 1640 38440 1710
rect 38440 1640 38470 1710
rect 38230 1620 38470 1640
rect 38230 1550 38260 1620
rect 38260 1550 38280 1620
rect 38280 1550 38350 1620
rect 38350 1550 38370 1620
rect 38370 1550 38440 1620
rect 38440 1550 38470 1620
rect 38230 1530 38470 1550
rect 38230 1510 38260 1530
rect 38260 1510 38280 1530
rect 38280 1510 38350 1530
rect 38350 1510 38370 1530
rect 38370 1510 38440 1530
rect 38440 1510 38470 1530
rect 38230 1370 38260 1420
rect 38260 1370 38280 1420
rect 38280 1370 38350 1420
rect 38350 1370 38370 1420
rect 38370 1370 38440 1420
rect 38440 1370 38470 1420
rect 38230 1350 38470 1370
rect 38230 1280 38260 1350
rect 38260 1280 38280 1350
rect 38280 1280 38350 1350
rect 38350 1280 38370 1350
rect 38370 1280 38440 1350
rect 38440 1280 38470 1350
rect 38230 1260 38470 1280
rect 38230 1190 38260 1260
rect 38260 1190 38280 1260
rect 38280 1190 38350 1260
rect 38350 1190 38370 1260
rect 38370 1190 38440 1260
rect 38440 1190 38470 1260
rect 38230 1180 38470 1190
rect 22480 -3760 22540 -3690
rect 22540 -3760 22580 -3690
rect 22580 -3760 22650 -3690
rect 22650 -3760 22690 -3690
rect 22690 -3760 22760 -3690
rect 22760 -3760 22800 -3690
rect 22800 -3760 22850 -3690
rect 22480 -3800 22850 -3760
rect 22480 -3870 22540 -3800
rect 22540 -3870 22580 -3800
rect 22580 -3870 22650 -3800
rect 22650 -3870 22690 -3800
rect 22690 -3870 22760 -3800
rect 22760 -3870 22800 -3800
rect 22800 -3870 22850 -3800
rect 22480 -3930 22850 -3870
rect 26960 -3760 27020 -3690
rect 27020 -3760 27060 -3690
rect 27060 -3760 27130 -3690
rect 27130 -3760 27170 -3690
rect 27170 -3760 27240 -3690
rect 27240 -3760 27280 -3690
rect 27280 -3760 27330 -3690
rect 26960 -3800 27330 -3760
rect 26960 -3870 27020 -3800
rect 27020 -3870 27060 -3800
rect 27060 -3870 27130 -3800
rect 27130 -3870 27170 -3800
rect 27170 -3870 27240 -3800
rect 27240 -3870 27280 -3800
rect 27280 -3870 27330 -3800
rect 26960 -3930 27330 -3870
rect -1170 -6400 -1160 -6370
rect -1160 -6400 -1090 -6370
rect -1090 -6400 -1070 -6370
rect -1070 -6400 -1000 -6370
rect -1000 -6400 -980 -6370
rect -980 -6400 -930 -6370
rect -840 -6400 -820 -6370
rect -820 -6400 -800 -6370
rect -800 -6400 -730 -6370
rect -730 -6400 -710 -6370
rect -710 -6400 -640 -6370
rect -640 -6400 -620 -6370
rect -620 -6400 -600 -6370
rect -510 -6400 -460 -6370
rect -460 -6400 -440 -6370
rect -440 -6400 -370 -6370
rect -370 -6400 -350 -6370
rect -350 -6400 -280 -6370
rect -280 -6400 -270 -6370
rect -180 -6400 -170 -6370
rect -170 -6400 -100 -6370
rect -100 -6400 -80 -6370
rect -80 -6400 -10 -6370
rect -10 -6400 10 -6370
rect 10 -6400 60 -6370
rect -1170 -6420 -930 -6400
rect -840 -6420 -600 -6400
rect -510 -6420 -270 -6400
rect -180 -6420 60 -6400
rect -1170 -6490 -1160 -6420
rect -1160 -6490 -1090 -6420
rect -1090 -6490 -1070 -6420
rect -1070 -6490 -1000 -6420
rect -1000 -6490 -980 -6420
rect -980 -6490 -930 -6420
rect -840 -6490 -820 -6420
rect -820 -6490 -800 -6420
rect -800 -6490 -730 -6420
rect -730 -6490 -710 -6420
rect -710 -6490 -640 -6420
rect -640 -6490 -620 -6420
rect -620 -6490 -600 -6420
rect -510 -6490 -460 -6420
rect -460 -6490 -440 -6420
rect -440 -6490 -370 -6420
rect -370 -6490 -350 -6420
rect -350 -6490 -280 -6420
rect -280 -6490 -270 -6420
rect -180 -6490 -170 -6420
rect -170 -6490 -100 -6420
rect -100 -6490 -80 -6420
rect -80 -6490 -10 -6420
rect -10 -6490 10 -6420
rect 10 -6490 60 -6420
rect -1170 -6510 -930 -6490
rect -840 -6510 -600 -6490
rect -510 -6510 -270 -6490
rect -180 -6510 60 -6490
rect -1170 -6580 -1160 -6510
rect -1160 -6580 -1090 -6510
rect -1090 -6580 -1070 -6510
rect -1070 -6580 -1000 -6510
rect -1000 -6580 -980 -6510
rect -980 -6580 -930 -6510
rect -840 -6580 -820 -6510
rect -820 -6580 -800 -6510
rect -800 -6580 -730 -6510
rect -730 -6580 -710 -6510
rect -710 -6580 -640 -6510
rect -640 -6580 -620 -6510
rect -620 -6580 -600 -6510
rect -510 -6580 -460 -6510
rect -460 -6580 -440 -6510
rect -440 -6580 -370 -6510
rect -370 -6580 -350 -6510
rect -350 -6580 -280 -6510
rect -280 -6580 -270 -6510
rect -180 -6580 -170 -6510
rect -170 -6580 -100 -6510
rect -100 -6580 -80 -6510
rect -80 -6580 -10 -6510
rect -10 -6580 10 -6510
rect 10 -6580 60 -6510
rect -1170 -6610 -930 -6580
rect -840 -6610 -600 -6580
rect -510 -6610 -270 -6580
rect -180 -6610 60 -6580
rect 14720 -6400 14770 -6370
rect 14770 -6400 14790 -6370
rect 14790 -6400 14860 -6370
rect 14860 -6400 14880 -6370
rect 14880 -6400 14950 -6370
rect 14950 -6400 14960 -6370
rect 15050 -6400 15060 -6370
rect 15060 -6400 15130 -6370
rect 15130 -6400 15150 -6370
rect 15150 -6400 15220 -6370
rect 15220 -6400 15240 -6370
rect 15240 -6400 15290 -6370
rect 15380 -6400 15400 -6370
rect 15400 -6400 15420 -6370
rect 15420 -6400 15490 -6370
rect 15490 -6400 15510 -6370
rect 15510 -6400 15580 -6370
rect 15580 -6400 15600 -6370
rect 15600 -6400 15620 -6370
rect 15710 -6400 15760 -6370
rect 15760 -6400 15780 -6370
rect 15780 -6400 15850 -6370
rect 15850 -6400 15870 -6370
rect 15870 -6400 15940 -6370
rect 15940 -6400 15950 -6370
rect 14720 -6420 14960 -6400
rect 15050 -6420 15290 -6400
rect 15380 -6420 15620 -6400
rect 15710 -6420 15950 -6400
rect 14720 -6490 14770 -6420
rect 14770 -6490 14790 -6420
rect 14790 -6490 14860 -6420
rect 14860 -6490 14880 -6420
rect 14880 -6490 14950 -6420
rect 14950 -6490 14960 -6420
rect 15050 -6490 15060 -6420
rect 15060 -6490 15130 -6420
rect 15130 -6490 15150 -6420
rect 15150 -6490 15220 -6420
rect 15220 -6490 15240 -6420
rect 15240 -6490 15290 -6420
rect 15380 -6490 15400 -6420
rect 15400 -6490 15420 -6420
rect 15420 -6490 15490 -6420
rect 15490 -6490 15510 -6420
rect 15510 -6490 15580 -6420
rect 15580 -6490 15600 -6420
rect 15600 -6490 15620 -6420
rect 15710 -6490 15760 -6420
rect 15760 -6490 15780 -6420
rect 15780 -6490 15850 -6420
rect 15850 -6490 15870 -6420
rect 15870 -6490 15940 -6420
rect 15940 -6490 15950 -6420
rect 14720 -6510 14960 -6490
rect 15050 -6510 15290 -6490
rect 15380 -6510 15620 -6490
rect 15710 -6510 15950 -6490
rect 14720 -6580 14770 -6510
rect 14770 -6580 14790 -6510
rect 14790 -6580 14860 -6510
rect 14860 -6580 14880 -6510
rect 14880 -6580 14950 -6510
rect 14950 -6580 14960 -6510
rect 15050 -6580 15060 -6510
rect 15060 -6580 15130 -6510
rect 15130 -6580 15150 -6510
rect 15150 -6580 15220 -6510
rect 15220 -6580 15240 -6510
rect 15240 -6580 15290 -6510
rect 15380 -6580 15400 -6510
rect 15400 -6580 15420 -6510
rect 15420 -6580 15490 -6510
rect 15490 -6580 15510 -6510
rect 15510 -6580 15580 -6510
rect 15580 -6580 15600 -6510
rect 15600 -6580 15620 -6510
rect 15710 -6580 15760 -6510
rect 15760 -6580 15780 -6510
rect 15780 -6580 15850 -6510
rect 15850 -6580 15870 -6510
rect 15870 -6580 15940 -6510
rect 15940 -6580 15950 -6510
rect 14720 -6610 14960 -6580
rect 15050 -6610 15290 -6580
rect 15380 -6610 15620 -6580
rect 15710 -6610 15950 -6580
rect 21650 -8430 21700 -8370
rect 21700 -8430 21730 -8370
rect 21730 -8430 21800 -8370
rect 21800 -8430 21830 -8370
rect 21830 -8430 21890 -8370
rect 21650 -8460 21890 -8430
rect 21650 -8530 21700 -8460
rect 21700 -8530 21730 -8460
rect 21730 -8530 21800 -8460
rect 21800 -8530 21830 -8460
rect 21830 -8530 21890 -8460
rect 21650 -8560 21890 -8530
rect 21650 -8610 21700 -8560
rect 21700 -8610 21730 -8560
rect 21730 -8610 21800 -8560
rect 21800 -8610 21830 -8560
rect 21830 -8610 21890 -8560
rect 1260 -10410 1330 -10340
rect 1330 -10410 1370 -10340
rect 1370 -10410 1440 -10340
rect 1440 -10410 1480 -10340
rect 1480 -10410 1500 -10340
rect 1590 -10410 1660 -10340
rect 1660 -10410 1700 -10340
rect 1700 -10410 1770 -10340
rect 1770 -10410 1810 -10340
rect 1810 -10410 1830 -10340
rect 1930 -10410 1990 -10340
rect 1990 -10410 2030 -10340
rect 2030 -10410 2100 -10340
rect 2100 -10410 2140 -10340
rect 2140 -10410 2170 -10340
rect 2260 -10410 2320 -10340
rect 2320 -10410 2360 -10340
rect 2360 -10410 2430 -10340
rect 2430 -10410 2470 -10340
rect 2470 -10410 2500 -10340
rect 1260 -10450 1500 -10410
rect 1590 -10450 1830 -10410
rect 1930 -10450 2170 -10410
rect 2260 -10450 2500 -10410
rect 1260 -10520 1330 -10450
rect 1330 -10520 1370 -10450
rect 1370 -10520 1440 -10450
rect 1440 -10520 1480 -10450
rect 1480 -10520 1500 -10450
rect 1590 -10520 1660 -10450
rect 1660 -10520 1700 -10450
rect 1700 -10520 1770 -10450
rect 1770 -10520 1810 -10450
rect 1810 -10520 1830 -10450
rect 1930 -10520 1990 -10450
rect 1990 -10520 2030 -10450
rect 2030 -10520 2100 -10450
rect 2100 -10520 2140 -10450
rect 2140 -10520 2170 -10450
rect 2260 -10520 2320 -10450
rect 2320 -10520 2360 -10450
rect 2360 -10520 2430 -10450
rect 2430 -10520 2470 -10450
rect 2470 -10520 2500 -10450
rect 1260 -10580 1500 -10520
rect 1590 -10580 1830 -10520
rect 1930 -10580 2170 -10520
rect 2260 -10580 2500 -10520
rect 12400 -10440 12470 -10370
rect 12470 -10440 12510 -10370
rect 12510 -10440 12580 -10370
rect 12580 -10440 12620 -10370
rect 12620 -10440 12640 -10370
rect 12730 -10440 12800 -10370
rect 12800 -10440 12840 -10370
rect 12840 -10440 12910 -10370
rect 12910 -10440 12950 -10370
rect 12950 -10440 12970 -10370
rect 13070 -10440 13130 -10370
rect 13130 -10440 13170 -10370
rect 13170 -10440 13240 -10370
rect 13240 -10440 13280 -10370
rect 13280 -10440 13310 -10370
rect 13400 -10440 13460 -10370
rect 13460 -10440 13500 -10370
rect 13500 -10440 13570 -10370
rect 13570 -10440 13610 -10370
rect 13610 -10440 13640 -10370
rect 12400 -10480 12640 -10440
rect 12730 -10480 12970 -10440
rect 13070 -10480 13310 -10440
rect 13400 -10480 13640 -10440
rect 12400 -10550 12470 -10480
rect 12470 -10550 12510 -10480
rect 12510 -10550 12580 -10480
rect 12580 -10550 12620 -10480
rect 12620 -10550 12640 -10480
rect 12730 -10550 12800 -10480
rect 12800 -10550 12840 -10480
rect 12840 -10550 12910 -10480
rect 12910 -10550 12950 -10480
rect 12950 -10550 12970 -10480
rect 13070 -10550 13130 -10480
rect 13130 -10550 13170 -10480
rect 13170 -10550 13240 -10480
rect 13240 -10550 13280 -10480
rect 13280 -10550 13310 -10480
rect 13400 -10550 13460 -10480
rect 13460 -10550 13500 -10480
rect 13500 -10550 13570 -10480
rect 13570 -10550 13610 -10480
rect 13610 -10550 13640 -10480
rect 12400 -10610 12640 -10550
rect 12730 -10610 12970 -10550
rect 13070 -10610 13310 -10550
rect 13400 -10610 13640 -10550
rect 38230 150 38260 170
rect 38260 150 38280 170
rect 38280 150 38350 170
rect 38350 150 38370 170
rect 38370 150 38440 170
rect 38440 150 38470 170
rect 38230 130 38470 150
rect 38230 60 38260 130
rect 38260 60 38280 130
rect 38280 60 38350 130
rect 38350 60 38370 130
rect 38370 60 38440 130
rect 38440 60 38470 130
rect 38230 40 38470 60
rect 38230 -30 38260 40
rect 38260 -30 38280 40
rect 38280 -30 38350 40
rect 38350 -30 38370 40
rect 38370 -30 38440 40
rect 38440 -30 38470 40
rect 38230 -50 38470 -30
rect 38230 -70 38260 -50
rect 38260 -70 38280 -50
rect 38280 -70 38350 -50
rect 38350 -70 38370 -50
rect 38370 -70 38440 -50
rect 38440 -70 38470 -50
rect 38230 -210 38260 -160
rect 38260 -210 38280 -160
rect 38280 -210 38350 -160
rect 38350 -210 38370 -160
rect 38370 -210 38440 -160
rect 38440 -210 38470 -160
rect 38230 -230 38470 -210
rect 38230 -300 38260 -230
rect 38260 -300 38280 -230
rect 38280 -300 38350 -230
rect 38350 -300 38370 -230
rect 38370 -300 38440 -230
rect 38440 -300 38470 -230
rect 38230 -320 38470 -300
rect 38230 -390 38260 -320
rect 38260 -390 38280 -320
rect 38280 -390 38350 -320
rect 38350 -390 38370 -320
rect 38370 -390 38440 -320
rect 38440 -390 38470 -320
rect 38230 -400 38470 -390
rect 38230 -540 38470 -530
rect 38230 -610 38260 -540
rect 38260 -610 38280 -540
rect 38280 -610 38350 -540
rect 38350 -610 38370 -540
rect 38370 -610 38440 -540
rect 38440 -610 38470 -540
rect 38230 -630 38470 -610
rect 38230 -700 38260 -630
rect 38260 -700 38280 -630
rect 38280 -700 38350 -630
rect 38350 -700 38370 -630
rect 38370 -700 38440 -630
rect 38440 -700 38470 -630
rect 38230 -720 38470 -700
rect 38230 -770 38260 -720
rect 38260 -770 38280 -720
rect 38280 -770 38350 -720
rect 38350 -770 38370 -720
rect 38370 -770 38440 -720
rect 38440 -770 38470 -720
rect 38230 -880 38260 -860
rect 38260 -880 38280 -860
rect 38280 -880 38350 -860
rect 38350 -880 38370 -860
rect 38370 -880 38440 -860
rect 38440 -880 38470 -860
rect 38230 -900 38470 -880
rect 38230 -970 38260 -900
rect 38260 -970 38280 -900
rect 38280 -970 38350 -900
rect 38350 -970 38370 -900
rect 38370 -970 38440 -900
rect 38440 -970 38470 -900
rect 38230 -990 38470 -970
rect 38230 -1060 38260 -990
rect 38260 -1060 38280 -990
rect 38280 -1060 38350 -990
rect 38350 -1060 38370 -990
rect 38370 -1060 38440 -990
rect 38440 -1060 38470 -990
rect 38230 -1080 38470 -1060
rect 38230 -1100 38260 -1080
rect 38260 -1100 38280 -1080
rect 38280 -1100 38350 -1080
rect 38350 -1100 38370 -1080
rect 38370 -1100 38440 -1080
rect 38440 -1100 38470 -1080
rect 38230 -1240 38260 -1190
rect 38260 -1240 38280 -1190
rect 38280 -1240 38350 -1190
rect 38350 -1240 38370 -1190
rect 38370 -1240 38440 -1190
rect 38440 -1240 38470 -1190
rect 38230 -1260 38470 -1240
rect 38230 -1330 38260 -1260
rect 38260 -1330 38280 -1260
rect 38280 -1330 38350 -1260
rect 38350 -1330 38370 -1260
rect 38370 -1330 38440 -1260
rect 38440 -1330 38470 -1260
rect 38230 -1350 38470 -1330
rect 38230 -1420 38260 -1350
rect 38260 -1420 38280 -1350
rect 38280 -1420 38350 -1350
rect 38350 -1420 38370 -1350
rect 38370 -1420 38440 -1350
rect 38440 -1420 38470 -1350
rect 38230 -1430 38470 -1420
rect 38230 -1530 38470 -1520
rect 38230 -1600 38260 -1530
rect 38260 -1600 38280 -1530
rect 38280 -1600 38350 -1530
rect 38350 -1600 38370 -1530
rect 38370 -1600 38440 -1530
rect 38440 -1600 38470 -1530
rect 38230 -1620 38470 -1600
rect 38230 -1690 38260 -1620
rect 38260 -1690 38280 -1620
rect 38280 -1690 38350 -1620
rect 38350 -1690 38370 -1620
rect 38370 -1690 38440 -1620
rect 38440 -1690 38470 -1620
rect 38230 -1710 38470 -1690
rect 38230 -1760 38260 -1710
rect 38260 -1760 38280 -1710
rect 38280 -1760 38350 -1710
rect 38350 -1760 38370 -1710
rect 38370 -1760 38440 -1710
rect 38440 -1760 38470 -1710
rect 38230 -1870 38260 -1850
rect 38260 -1870 38280 -1850
rect 38280 -1870 38350 -1850
rect 38350 -1870 38370 -1850
rect 38370 -1870 38440 -1850
rect 38440 -1870 38470 -1850
rect 38230 -1890 38470 -1870
rect 38230 -1960 38260 -1890
rect 38260 -1960 38280 -1890
rect 38280 -1960 38350 -1890
rect 38350 -1960 38370 -1890
rect 38370 -1960 38440 -1890
rect 38440 -1960 38470 -1890
rect 38230 -1980 38470 -1960
rect 38230 -2050 38260 -1980
rect 38260 -2050 38280 -1980
rect 38280 -2050 38350 -1980
rect 38350 -2050 38370 -1980
rect 38370 -2050 38440 -1980
rect 38440 -2050 38470 -1980
rect 38230 -2070 38470 -2050
rect 38230 -2090 38260 -2070
rect 38260 -2090 38280 -2070
rect 38280 -2090 38350 -2070
rect 38350 -2090 38370 -2070
rect 38370 -2090 38440 -2070
rect 38440 -2090 38470 -2070
rect 38230 -2230 38260 -2180
rect 38260 -2230 38280 -2180
rect 38280 -2230 38350 -2180
rect 38350 -2230 38370 -2180
rect 38370 -2230 38440 -2180
rect 38440 -2230 38470 -2180
rect 38230 -2250 38470 -2230
rect 38230 -2320 38260 -2250
rect 38260 -2320 38280 -2250
rect 38280 -2320 38350 -2250
rect 38350 -2320 38370 -2250
rect 38370 -2320 38440 -2250
rect 38440 -2320 38470 -2250
rect 38230 -2340 38470 -2320
rect 38230 -2410 38260 -2340
rect 38260 -2410 38280 -2340
rect 38280 -2410 38350 -2340
rect 38350 -2410 38370 -2340
rect 38370 -2410 38440 -2340
rect 38440 -2410 38470 -2340
rect 38230 -2420 38470 -2410
rect 38230 -2520 38470 -2510
rect 38230 -2590 38260 -2520
rect 38260 -2590 38280 -2520
rect 38280 -2590 38350 -2520
rect 38350 -2590 38370 -2520
rect 38370 -2590 38440 -2520
rect 38440 -2590 38470 -2520
rect 38230 -2610 38470 -2590
rect 38230 -2680 38260 -2610
rect 38260 -2680 38280 -2610
rect 38280 -2680 38350 -2610
rect 38350 -2680 38370 -2610
rect 38370 -2680 38440 -2610
rect 38440 -2680 38470 -2610
rect 38230 -2700 38470 -2680
rect 38230 -2750 38260 -2700
rect 38260 -2750 38280 -2700
rect 38280 -2750 38350 -2700
rect 38350 -2750 38370 -2700
rect 38370 -2750 38440 -2700
rect 38440 -2750 38470 -2700
rect 38230 -2860 38260 -2840
rect 38260 -2860 38280 -2840
rect 38280 -2860 38350 -2840
rect 38350 -2860 38370 -2840
rect 38370 -2860 38440 -2840
rect 38440 -2860 38470 -2840
rect 38230 -2880 38470 -2860
rect 38230 -2950 38260 -2880
rect 38260 -2950 38280 -2880
rect 38280 -2950 38350 -2880
rect 38350 -2950 38370 -2880
rect 38370 -2950 38440 -2880
rect 38440 -2950 38470 -2880
rect 38230 -2970 38470 -2950
rect 38230 -3040 38260 -2970
rect 38260 -3040 38280 -2970
rect 38280 -3040 38350 -2970
rect 38350 -3040 38370 -2970
rect 38370 -3040 38440 -2970
rect 38440 -3040 38470 -2970
rect 38230 -3060 38470 -3040
rect 38230 -3080 38260 -3060
rect 38260 -3080 38280 -3060
rect 38280 -3080 38350 -3060
rect 38350 -3080 38370 -3060
rect 38370 -3080 38440 -3060
rect 38440 -3080 38470 -3060
rect 38230 -3220 38260 -3170
rect 38260 -3220 38280 -3170
rect 38280 -3220 38350 -3170
rect 38350 -3220 38370 -3170
rect 38370 -3220 38440 -3170
rect 38440 -3220 38470 -3170
rect 38230 -3240 38470 -3220
rect 38230 -3310 38260 -3240
rect 38260 -3310 38280 -3240
rect 38280 -3310 38350 -3240
rect 38350 -3310 38370 -3240
rect 38370 -3310 38440 -3240
rect 38440 -3310 38470 -3240
rect 38230 -3330 38470 -3310
rect 38230 -3400 38260 -3330
rect 38260 -3400 38280 -3330
rect 38280 -3400 38350 -3330
rect 38350 -3400 38370 -3330
rect 38370 -3400 38440 -3330
rect 38440 -3400 38470 -3330
rect 38230 -3410 38470 -3400
rect 38230 -3550 38470 -3540
rect 38230 -3620 38260 -3550
rect 38260 -3620 38280 -3550
rect 38280 -3620 38350 -3550
rect 38350 -3620 38370 -3550
rect 38370 -3620 38440 -3550
rect 38440 -3620 38470 -3550
rect 38230 -3640 38470 -3620
rect 38230 -3710 38260 -3640
rect 38260 -3710 38280 -3640
rect 38280 -3710 38350 -3640
rect 38350 -3710 38370 -3640
rect 38370 -3710 38440 -3640
rect 38440 -3710 38470 -3640
rect 38230 -3730 38470 -3710
rect 38230 -3780 38260 -3730
rect 38260 -3780 38280 -3730
rect 38280 -3780 38350 -3730
rect 38350 -3780 38370 -3730
rect 38370 -3780 38440 -3730
rect 38440 -3780 38470 -3730
rect 38230 -3890 38260 -3870
rect 38260 -3890 38280 -3870
rect 38280 -3890 38350 -3870
rect 38350 -3890 38370 -3870
rect 38370 -3890 38440 -3870
rect 38440 -3890 38470 -3870
rect 38230 -3910 38470 -3890
rect 38230 -3980 38260 -3910
rect 38260 -3980 38280 -3910
rect 38280 -3980 38350 -3910
rect 38350 -3980 38370 -3910
rect 38370 -3980 38440 -3910
rect 38440 -3980 38470 -3910
rect 38230 -4000 38470 -3980
rect 38230 -4070 38260 -4000
rect 38260 -4070 38280 -4000
rect 38280 -4070 38350 -4000
rect 38350 -4070 38370 -4000
rect 38370 -4070 38440 -4000
rect 38440 -4070 38470 -4000
rect 38230 -4090 38470 -4070
rect 38230 -4110 38260 -4090
rect 38260 -4110 38280 -4090
rect 38280 -4110 38350 -4090
rect 38350 -4110 38370 -4090
rect 38370 -4110 38440 -4090
rect 38440 -4110 38470 -4090
rect 38230 -4250 38260 -4200
rect 38260 -4250 38280 -4200
rect 38280 -4250 38350 -4200
rect 38350 -4250 38370 -4200
rect 38370 -4250 38440 -4200
rect 38440 -4250 38470 -4200
rect 38230 -4270 38470 -4250
rect 38230 -4340 38260 -4270
rect 38260 -4340 38280 -4270
rect 38280 -4340 38350 -4270
rect 38350 -4340 38370 -4270
rect 38370 -4340 38440 -4270
rect 38440 -4340 38470 -4270
rect 38230 -4360 38470 -4340
rect 38230 -4430 38260 -4360
rect 38260 -4430 38280 -4360
rect 38280 -4430 38350 -4360
rect 38350 -4430 38370 -4360
rect 38370 -4430 38440 -4360
rect 38440 -4430 38470 -4360
rect 38230 -4440 38470 -4430
rect 38230 -4540 38470 -4530
rect 38230 -4610 38260 -4540
rect 38260 -4610 38280 -4540
rect 38280 -4610 38350 -4540
rect 38350 -4610 38370 -4540
rect 38370 -4610 38440 -4540
rect 38440 -4610 38470 -4540
rect 38230 -4630 38470 -4610
rect 38230 -4700 38260 -4630
rect 38260 -4700 38280 -4630
rect 38280 -4700 38350 -4630
rect 38350 -4700 38370 -4630
rect 38370 -4700 38440 -4630
rect 38440 -4700 38470 -4630
rect 38230 -4720 38470 -4700
rect 38230 -4770 38260 -4720
rect 38260 -4770 38280 -4720
rect 38280 -4770 38350 -4720
rect 38350 -4770 38370 -4720
rect 38370 -4770 38440 -4720
rect 38440 -4770 38470 -4720
rect 38230 -4880 38260 -4860
rect 38260 -4880 38280 -4860
rect 38280 -4880 38350 -4860
rect 38350 -4880 38370 -4860
rect 38370 -4880 38440 -4860
rect 38440 -4880 38470 -4860
rect 38230 -4900 38470 -4880
rect 38230 -4970 38260 -4900
rect 38260 -4970 38280 -4900
rect 38280 -4970 38350 -4900
rect 38350 -4970 38370 -4900
rect 38370 -4970 38440 -4900
rect 38440 -4970 38470 -4900
rect 38230 -4990 38470 -4970
rect 38230 -5060 38260 -4990
rect 38260 -5060 38280 -4990
rect 38280 -5060 38350 -4990
rect 38350 -5060 38370 -4990
rect 38370 -5060 38440 -4990
rect 38440 -5060 38470 -4990
rect 38230 -5080 38470 -5060
rect 38230 -5100 38260 -5080
rect 38260 -5100 38280 -5080
rect 38280 -5100 38350 -5080
rect 38350 -5100 38370 -5080
rect 38370 -5100 38440 -5080
rect 38440 -5100 38470 -5080
rect 38230 -5240 38260 -5190
rect 38260 -5240 38280 -5190
rect 38280 -5240 38350 -5190
rect 38350 -5240 38370 -5190
rect 38370 -5240 38440 -5190
rect 38440 -5240 38470 -5190
rect 38230 -5260 38470 -5240
rect 38230 -5330 38260 -5260
rect 38260 -5330 38280 -5260
rect 38280 -5330 38350 -5260
rect 38350 -5330 38370 -5260
rect 38370 -5330 38440 -5260
rect 38440 -5330 38470 -5260
rect 38230 -5350 38470 -5330
rect 38230 -5420 38260 -5350
rect 38260 -5420 38280 -5350
rect 38280 -5420 38350 -5350
rect 38350 -5420 38370 -5350
rect 38370 -5420 38440 -5350
rect 38440 -5420 38470 -5350
rect 38230 -5430 38470 -5420
rect 38230 -5530 38470 -5520
rect 38230 -5600 38260 -5530
rect 38260 -5600 38280 -5530
rect 38280 -5600 38350 -5530
rect 38350 -5600 38370 -5530
rect 38370 -5600 38440 -5530
rect 38440 -5600 38470 -5530
rect 38230 -5620 38470 -5600
rect 38230 -5690 38260 -5620
rect 38260 -5690 38280 -5620
rect 38280 -5690 38350 -5620
rect 38350 -5690 38370 -5620
rect 38370 -5690 38440 -5620
rect 38440 -5690 38470 -5620
rect 38230 -5710 38470 -5690
rect 38230 -5760 38260 -5710
rect 38260 -5760 38280 -5710
rect 38280 -5760 38350 -5710
rect 38350 -5760 38370 -5710
rect 38370 -5760 38440 -5710
rect 38440 -5760 38470 -5710
rect 38230 -5870 38260 -5850
rect 38260 -5870 38280 -5850
rect 38280 -5870 38350 -5850
rect 38350 -5870 38370 -5850
rect 38370 -5870 38440 -5850
rect 38440 -5870 38470 -5850
rect 38230 -5890 38470 -5870
rect 38230 -5960 38260 -5890
rect 38260 -5960 38280 -5890
rect 38280 -5960 38350 -5890
rect 38350 -5960 38370 -5890
rect 38370 -5960 38440 -5890
rect 38440 -5960 38470 -5890
rect 38230 -5980 38470 -5960
rect 38230 -6050 38260 -5980
rect 38260 -6050 38280 -5980
rect 38280 -6050 38350 -5980
rect 38350 -6050 38370 -5980
rect 38370 -6050 38440 -5980
rect 38440 -6050 38470 -5980
rect 38230 -6070 38470 -6050
rect 38230 -6090 38260 -6070
rect 38260 -6090 38280 -6070
rect 38280 -6090 38350 -6070
rect 38350 -6090 38370 -6070
rect 38370 -6090 38440 -6070
rect 38440 -6090 38470 -6070
rect 38230 -6230 38260 -6180
rect 38260 -6230 38280 -6180
rect 38280 -6230 38350 -6180
rect 38350 -6230 38370 -6180
rect 38370 -6230 38440 -6180
rect 38440 -6230 38470 -6180
rect 38230 -6250 38470 -6230
rect 38230 -6320 38260 -6250
rect 38260 -6320 38280 -6250
rect 38280 -6320 38350 -6250
rect 38350 -6320 38370 -6250
rect 38370 -6320 38440 -6250
rect 38440 -6320 38470 -6250
rect 38230 -6340 38470 -6320
rect 38230 -6410 38260 -6340
rect 38260 -6410 38280 -6340
rect 38280 -6410 38350 -6340
rect 38350 -6410 38370 -6340
rect 38370 -6410 38440 -6340
rect 38440 -6410 38470 -6340
rect 38230 -6420 38470 -6410
rect 1690 -12300 1930 -12240
rect 2020 -12300 2260 -12240
rect 2360 -12300 2600 -12240
rect 2690 -12300 2930 -12240
rect 1690 -12370 1720 -12300
rect 1720 -12370 1760 -12300
rect 1760 -12370 1830 -12300
rect 1830 -12370 1870 -12300
rect 1870 -12370 1930 -12300
rect 2020 -12370 2050 -12300
rect 2050 -12370 2090 -12300
rect 2090 -12370 2160 -12300
rect 2160 -12370 2200 -12300
rect 2200 -12370 2260 -12300
rect 2360 -12370 2380 -12300
rect 2380 -12370 2420 -12300
rect 2420 -12370 2490 -12300
rect 2490 -12370 2530 -12300
rect 2530 -12370 2600 -12300
rect 2690 -12370 2710 -12300
rect 2710 -12370 2750 -12300
rect 2750 -12370 2820 -12300
rect 2820 -12370 2860 -12300
rect 2860 -12370 2930 -12300
rect 1690 -12410 1930 -12370
rect 2020 -12410 2260 -12370
rect 2360 -12410 2600 -12370
rect 2690 -12410 2930 -12370
rect 1690 -12480 1720 -12410
rect 1720 -12480 1760 -12410
rect 1760 -12480 1830 -12410
rect 1830 -12480 1870 -12410
rect 1870 -12480 1930 -12410
rect 2020 -12480 2050 -12410
rect 2050 -12480 2090 -12410
rect 2090 -12480 2160 -12410
rect 2160 -12480 2200 -12410
rect 2200 -12480 2260 -12410
rect 2360 -12480 2380 -12410
rect 2380 -12480 2420 -12410
rect 2420 -12480 2490 -12410
rect 2490 -12480 2530 -12410
rect 2530 -12480 2600 -12410
rect 2690 -12480 2710 -12410
rect 2710 -12480 2750 -12410
rect 2750 -12480 2820 -12410
rect 2820 -12480 2860 -12410
rect 2860 -12480 2930 -12410
rect 11970 -12300 12210 -12240
rect 12300 -12300 12540 -12240
rect 12640 -12300 12880 -12240
rect 12970 -12300 13210 -12240
rect 11970 -12370 12000 -12300
rect 12000 -12370 12040 -12300
rect 12040 -12370 12110 -12300
rect 12110 -12370 12150 -12300
rect 12150 -12370 12210 -12300
rect 12300 -12370 12330 -12300
rect 12330 -12370 12370 -12300
rect 12370 -12370 12440 -12300
rect 12440 -12370 12480 -12300
rect 12480 -12370 12540 -12300
rect 12640 -12370 12660 -12300
rect 12660 -12370 12700 -12300
rect 12700 -12370 12770 -12300
rect 12770 -12370 12810 -12300
rect 12810 -12370 12880 -12300
rect 12970 -12370 12990 -12300
rect 12990 -12370 13030 -12300
rect 13030 -12370 13100 -12300
rect 13100 -12370 13140 -12300
rect 13140 -12370 13210 -12300
rect 11970 -12410 12210 -12370
rect 12300 -12410 12540 -12370
rect 12640 -12410 12880 -12370
rect 12970 -12410 13210 -12370
rect 11970 -12480 12000 -12410
rect 12000 -12480 12040 -12410
rect 12040 -12480 12110 -12410
rect 12110 -12480 12150 -12410
rect 12150 -12480 12210 -12410
rect 12300 -12480 12330 -12410
rect 12330 -12480 12370 -12410
rect 12370 -12480 12440 -12410
rect 12440 -12480 12480 -12410
rect 12480 -12480 12540 -12410
rect 12640 -12480 12660 -12410
rect 12660 -12480 12700 -12410
rect 12700 -12480 12770 -12410
rect 12770 -12480 12810 -12410
rect 12810 -12480 12880 -12410
rect 12970 -12480 12990 -12410
rect 12990 -12480 13030 -12410
rect 13030 -12480 13100 -12410
rect 13100 -12480 13140 -12410
rect 13140 -12480 13210 -12410
rect 21650 -14090 21700 -14030
rect 21700 -14090 21730 -14030
rect 21730 -14090 21800 -14030
rect 21800 -14090 21830 -14030
rect 21830 -14090 21890 -14030
rect 21650 -14120 21890 -14090
rect 21650 -14190 21700 -14120
rect 21700 -14190 21730 -14120
rect 21730 -14190 21800 -14120
rect 21800 -14190 21830 -14120
rect 21830 -14190 21890 -14120
rect 21650 -14220 21890 -14190
rect 21650 -14270 21700 -14220
rect 21700 -14270 21730 -14220
rect 21730 -14270 21800 -14220
rect 21800 -14270 21830 -14220
rect 21830 -14270 21890 -14220
rect 21650 -20170 21700 -20110
rect 21700 -20170 21730 -20110
rect 21730 -20170 21800 -20110
rect 21800 -20170 21830 -20110
rect 21830 -20170 21890 -20110
rect 21650 -20200 21890 -20170
rect 21650 -20270 21700 -20200
rect 21700 -20270 21730 -20200
rect 21730 -20270 21800 -20200
rect 21800 -20270 21830 -20200
rect 21830 -20270 21890 -20200
rect 21650 -20300 21890 -20270
rect 21650 -20350 21700 -20300
rect 21700 -20350 21730 -20300
rect 21730 -20350 21800 -20300
rect 21800 -20350 21830 -20300
rect 21830 -20350 21890 -20300
rect 1730 -22730 1800 -22660
rect 1800 -22730 1840 -22660
rect 1840 -22730 1910 -22660
rect 1910 -22730 1950 -22660
rect 1950 -22730 1970 -22660
rect 2060 -22730 2130 -22660
rect 2130 -22730 2170 -22660
rect 2170 -22730 2240 -22660
rect 2240 -22730 2280 -22660
rect 2280 -22730 2300 -22660
rect 2400 -22730 2460 -22660
rect 2460 -22730 2500 -22660
rect 2500 -22730 2570 -22660
rect 2570 -22730 2610 -22660
rect 2610 -22730 2640 -22660
rect 2730 -22730 2790 -22660
rect 2790 -22730 2830 -22660
rect 2830 -22730 2900 -22660
rect 2900 -22730 2940 -22660
rect 2940 -22730 2970 -22660
rect 1730 -22770 1970 -22730
rect 2060 -22770 2300 -22730
rect 2400 -22770 2640 -22730
rect 2730 -22770 2970 -22730
rect 1730 -22840 1800 -22770
rect 1800 -22840 1840 -22770
rect 1840 -22840 1910 -22770
rect 1910 -22840 1950 -22770
rect 1950 -22840 1970 -22770
rect 2060 -22840 2130 -22770
rect 2130 -22840 2170 -22770
rect 2170 -22840 2240 -22770
rect 2240 -22840 2280 -22770
rect 2280 -22840 2300 -22770
rect 2400 -22840 2460 -22770
rect 2460 -22840 2500 -22770
rect 2500 -22840 2570 -22770
rect 2570 -22840 2610 -22770
rect 2610 -22840 2640 -22770
rect 2730 -22840 2790 -22770
rect 2790 -22840 2830 -22770
rect 2830 -22840 2900 -22770
rect 2900 -22840 2940 -22770
rect 2940 -22840 2970 -22770
rect 1730 -22900 1970 -22840
rect 2060 -22900 2300 -22840
rect 2400 -22900 2640 -22840
rect 2730 -22900 2970 -22840
rect 11930 -22730 12000 -22660
rect 12000 -22730 12040 -22660
rect 12040 -22730 12110 -22660
rect 12110 -22730 12150 -22660
rect 12150 -22730 12170 -22660
rect 12260 -22730 12330 -22660
rect 12330 -22730 12370 -22660
rect 12370 -22730 12440 -22660
rect 12440 -22730 12480 -22660
rect 12480 -22730 12500 -22660
rect 12600 -22730 12660 -22660
rect 12660 -22730 12700 -22660
rect 12700 -22730 12770 -22660
rect 12770 -22730 12810 -22660
rect 12810 -22730 12840 -22660
rect 12930 -22730 12990 -22660
rect 12990 -22730 13030 -22660
rect 13030 -22730 13100 -22660
rect 13100 -22730 13140 -22660
rect 13140 -22730 13170 -22660
rect 11930 -22770 12170 -22730
rect 12260 -22770 12500 -22730
rect 12600 -22770 12840 -22730
rect 12930 -22770 13170 -22730
rect 11930 -22840 12000 -22770
rect 12000 -22840 12040 -22770
rect 12040 -22840 12110 -22770
rect 12110 -22840 12150 -22770
rect 12150 -22840 12170 -22770
rect 12260 -22840 12330 -22770
rect 12330 -22840 12370 -22770
rect 12370 -22840 12440 -22770
rect 12440 -22840 12480 -22770
rect 12480 -22840 12500 -22770
rect 12600 -22840 12660 -22770
rect 12660 -22840 12700 -22770
rect 12700 -22840 12770 -22770
rect 12770 -22840 12810 -22770
rect 12810 -22840 12840 -22770
rect 12930 -22840 12990 -22770
rect 12990 -22840 13030 -22770
rect 13030 -22840 13100 -22770
rect 13100 -22840 13140 -22770
rect 13140 -22840 13170 -22770
rect 11930 -22900 12170 -22840
rect 12260 -22900 12500 -22840
rect 12600 -22900 12840 -22840
rect 12930 -22900 13170 -22840
<< mimcap2 >>
rect -5510 20830 6730 20960
rect -5510 20590 -5200 20830
rect -4960 20590 -4870 20830
rect -4630 20590 -4540 20830
rect -4300 20590 -4210 20830
rect -3970 20590 -3880 20830
rect -3640 20590 -3550 20830
rect -3310 20590 -3220 20830
rect -2980 20590 -2890 20830
rect -2650 20590 -2560 20830
rect -2320 20590 -2230 20830
rect -1990 20590 -1900 20830
rect -1660 20590 -1570 20830
rect -1330 20590 -1240 20830
rect -1000 20590 -910 20830
rect -670 20590 -580 20830
rect -340 20590 -250 20830
rect -10 20590 80 20830
rect 320 20590 410 20830
rect 650 20590 740 20830
rect 980 20590 1070 20830
rect 1310 20590 1400 20830
rect 1640 20590 1730 20830
rect 1970 20590 2060 20830
rect 2300 20590 2390 20830
rect 2630 20590 2720 20830
rect 2960 20590 3050 20830
rect 3290 20590 3380 20830
rect 3620 20590 3710 20830
rect 3950 20590 4040 20830
rect 4280 20590 4370 20830
rect 4610 20590 4700 20830
rect 4940 20590 5030 20830
rect 5270 20590 5360 20830
rect 5600 20590 5690 20830
rect 5930 20590 6020 20830
rect 6260 20590 6350 20830
rect 6590 20590 6730 20830
rect -5510 20500 6730 20590
rect -5510 20260 -5200 20500
rect -4960 20260 -4870 20500
rect -4630 20260 -4540 20500
rect -4300 20260 -4210 20500
rect -3970 20260 -3880 20500
rect -3640 20260 -3550 20500
rect -3310 20260 -3220 20500
rect -2980 20260 -2890 20500
rect -2650 20260 -2560 20500
rect -2320 20260 -2230 20500
rect -1990 20260 -1900 20500
rect -1660 20260 -1570 20500
rect -1330 20260 -1240 20500
rect -1000 20260 -910 20500
rect -670 20260 -580 20500
rect -340 20260 -250 20500
rect -10 20260 80 20500
rect 320 20260 410 20500
rect 650 20260 740 20500
rect 980 20260 1070 20500
rect 1310 20260 1400 20500
rect 1640 20260 1730 20500
rect 1970 20260 2060 20500
rect 2300 20260 2390 20500
rect 2630 20260 2720 20500
rect 2960 20260 3050 20500
rect 3290 20260 3380 20500
rect 3620 20260 3710 20500
rect 3950 20260 4040 20500
rect 4280 20260 4370 20500
rect 4610 20260 4700 20500
rect 4940 20260 5030 20500
rect 5270 20260 5360 20500
rect 5600 20260 5690 20500
rect 5930 20260 6020 20500
rect 6260 20260 6350 20500
rect 6590 20260 6730 20500
rect -5510 20170 6730 20260
rect -5510 19930 -5200 20170
rect -4960 19930 -4870 20170
rect -4630 19930 -4540 20170
rect -4300 19930 -4210 20170
rect -3970 19930 -3880 20170
rect -3640 19930 -3550 20170
rect -3310 19930 -3220 20170
rect -2980 19930 -2890 20170
rect -2650 19930 -2560 20170
rect -2320 19930 -2230 20170
rect -1990 19930 -1900 20170
rect -1660 19930 -1570 20170
rect -1330 19930 -1240 20170
rect -1000 19930 -910 20170
rect -670 19930 -580 20170
rect -340 19930 -250 20170
rect -10 19930 80 20170
rect 320 19930 410 20170
rect 650 19930 740 20170
rect 980 19930 1070 20170
rect 1310 19930 1400 20170
rect 1640 19930 1730 20170
rect 1970 19930 2060 20170
rect 2300 19930 2390 20170
rect 2630 19930 2720 20170
rect 2960 19930 3050 20170
rect 3290 19930 3380 20170
rect 3620 19930 3710 20170
rect 3950 19930 4040 20170
rect 4280 19930 4370 20170
rect 4610 19930 4700 20170
rect 4940 19930 5030 20170
rect 5270 19930 5360 20170
rect 5600 19930 5690 20170
rect 5930 19930 6020 20170
rect 6260 19930 6350 20170
rect 6590 19930 6730 20170
rect -5510 19840 6730 19930
rect -5510 19600 -5200 19840
rect -4960 19600 -4870 19840
rect -4630 19600 -4540 19840
rect -4300 19600 -4210 19840
rect -3970 19600 -3880 19840
rect -3640 19600 -3550 19840
rect -3310 19600 -3220 19840
rect -2980 19600 -2890 19840
rect -2650 19600 -2560 19840
rect -2320 19600 -2230 19840
rect -1990 19600 -1900 19840
rect -1660 19600 -1570 19840
rect -1330 19600 -1240 19840
rect -1000 19600 -910 19840
rect -670 19600 -580 19840
rect -340 19600 -250 19840
rect -10 19600 80 19840
rect 320 19600 410 19840
rect 650 19600 740 19840
rect 980 19600 1070 19840
rect 1310 19600 1400 19840
rect 1640 19600 1730 19840
rect 1970 19600 2060 19840
rect 2300 19600 2390 19840
rect 2630 19600 2720 19840
rect 2960 19600 3050 19840
rect 3290 19600 3380 19840
rect 3620 19600 3710 19840
rect 3950 19600 4040 19840
rect 4280 19600 4370 19840
rect 4610 19600 4700 19840
rect 4940 19600 5030 19840
rect 5270 19600 5360 19840
rect 5600 19600 5690 19840
rect 5930 19600 6020 19840
rect 6260 19600 6350 19840
rect 6590 19600 6730 19840
rect -5510 19510 6730 19600
rect -5510 19270 -5200 19510
rect -4960 19270 -4870 19510
rect -4630 19270 -4540 19510
rect -4300 19270 -4210 19510
rect -3970 19270 -3880 19510
rect -3640 19270 -3550 19510
rect -3310 19270 -3220 19510
rect -2980 19270 -2890 19510
rect -2650 19270 -2560 19510
rect -2320 19270 -2230 19510
rect -1990 19270 -1900 19510
rect -1660 19270 -1570 19510
rect -1330 19270 -1240 19510
rect -1000 19270 -910 19510
rect -670 19270 -580 19510
rect -340 19270 -250 19510
rect -10 19270 80 19510
rect 320 19270 410 19510
rect 650 19270 740 19510
rect 980 19270 1070 19510
rect 1310 19270 1400 19510
rect 1640 19270 1730 19510
rect 1970 19270 2060 19510
rect 2300 19270 2390 19510
rect 2630 19270 2720 19510
rect 2960 19270 3050 19510
rect 3290 19270 3380 19510
rect 3620 19270 3710 19510
rect 3950 19270 4040 19510
rect 4280 19270 4370 19510
rect 4610 19270 4700 19510
rect 4940 19270 5030 19510
rect 5270 19270 5360 19510
rect 5600 19270 5690 19510
rect 5930 19270 6020 19510
rect 6260 19270 6350 19510
rect 6590 19270 6730 19510
rect -5510 19180 6730 19270
rect -5510 18940 -5200 19180
rect -4960 18940 -4870 19180
rect -4630 18940 -4540 19180
rect -4300 18940 -4210 19180
rect -3970 18940 -3880 19180
rect -3640 18940 -3550 19180
rect -3310 18940 -3220 19180
rect -2980 18940 -2890 19180
rect -2650 18940 -2560 19180
rect -2320 18940 -2230 19180
rect -1990 18940 -1900 19180
rect -1660 18940 -1570 19180
rect -1330 18940 -1240 19180
rect -1000 18940 -910 19180
rect -670 18940 -580 19180
rect -340 18940 -250 19180
rect -10 18940 80 19180
rect 320 18940 410 19180
rect 650 18940 740 19180
rect 980 18940 1070 19180
rect 1310 18940 1400 19180
rect 1640 18940 1730 19180
rect 1970 18940 2060 19180
rect 2300 18940 2390 19180
rect 2630 18940 2720 19180
rect 2960 18940 3050 19180
rect 3290 18940 3380 19180
rect 3620 18940 3710 19180
rect 3950 18940 4040 19180
rect 4280 18940 4370 19180
rect 4610 18940 4700 19180
rect 4940 18940 5030 19180
rect 5270 18940 5360 19180
rect 5600 18940 5690 19180
rect 5930 18940 6020 19180
rect 6260 18940 6350 19180
rect 6590 18940 6730 19180
rect -5510 18850 6730 18940
rect -5510 18610 -5200 18850
rect -4960 18610 -4870 18850
rect -4630 18610 -4540 18850
rect -4300 18610 -4210 18850
rect -3970 18610 -3880 18850
rect -3640 18610 -3550 18850
rect -3310 18610 -3220 18850
rect -2980 18610 -2890 18850
rect -2650 18610 -2560 18850
rect -2320 18610 -2230 18850
rect -1990 18610 -1900 18850
rect -1660 18610 -1570 18850
rect -1330 18610 -1240 18850
rect -1000 18610 -910 18850
rect -670 18610 -580 18850
rect -340 18610 -250 18850
rect -10 18610 80 18850
rect 320 18610 410 18850
rect 650 18610 740 18850
rect 980 18610 1070 18850
rect 1310 18610 1400 18850
rect 1640 18610 1730 18850
rect 1970 18610 2060 18850
rect 2300 18610 2390 18850
rect 2630 18610 2720 18850
rect 2960 18610 3050 18850
rect 3290 18610 3380 18850
rect 3620 18610 3710 18850
rect 3950 18610 4040 18850
rect 4280 18610 4370 18850
rect 4610 18610 4700 18850
rect 4940 18610 5030 18850
rect 5270 18610 5360 18850
rect 5600 18610 5690 18850
rect 5930 18610 6020 18850
rect 6260 18610 6350 18850
rect 6590 18610 6730 18850
rect -5510 18520 6730 18610
rect -5510 18280 -5200 18520
rect -4960 18280 -4870 18520
rect -4630 18280 -4540 18520
rect -4300 18280 -4210 18520
rect -3970 18280 -3880 18520
rect -3640 18280 -3550 18520
rect -3310 18280 -3220 18520
rect -2980 18280 -2890 18520
rect -2650 18280 -2560 18520
rect -2320 18280 -2230 18520
rect -1990 18280 -1900 18520
rect -1660 18280 -1570 18520
rect -1330 18280 -1240 18520
rect -1000 18280 -910 18520
rect -670 18280 -580 18520
rect -340 18280 -250 18520
rect -10 18280 80 18520
rect 320 18280 410 18520
rect 650 18280 740 18520
rect 980 18280 1070 18520
rect 1310 18280 1400 18520
rect 1640 18280 1730 18520
rect 1970 18280 2060 18520
rect 2300 18280 2390 18520
rect 2630 18280 2720 18520
rect 2960 18280 3050 18520
rect 3290 18280 3380 18520
rect 3620 18280 3710 18520
rect 3950 18280 4040 18520
rect 4280 18280 4370 18520
rect 4610 18280 4700 18520
rect 4940 18280 5030 18520
rect 5270 18280 5360 18520
rect 5600 18280 5690 18520
rect 5930 18280 6020 18520
rect 6260 18280 6350 18520
rect 6590 18280 6730 18520
rect -5510 18190 6730 18280
rect -5510 17950 -5200 18190
rect -4960 17950 -4870 18190
rect -4630 17950 -4540 18190
rect -4300 17950 -4210 18190
rect -3970 17950 -3880 18190
rect -3640 17950 -3550 18190
rect -3310 17950 -3220 18190
rect -2980 17950 -2890 18190
rect -2650 17950 -2560 18190
rect -2320 17950 -2230 18190
rect -1990 17950 -1900 18190
rect -1660 17950 -1570 18190
rect -1330 17950 -1240 18190
rect -1000 17950 -910 18190
rect -670 17950 -580 18190
rect -340 17950 -250 18190
rect -10 17950 80 18190
rect 320 17950 410 18190
rect 650 17950 740 18190
rect 980 17950 1070 18190
rect 1310 17950 1400 18190
rect 1640 17950 1730 18190
rect 1970 17950 2060 18190
rect 2300 17950 2390 18190
rect 2630 17950 2720 18190
rect 2960 17950 3050 18190
rect 3290 17950 3380 18190
rect 3620 17950 3710 18190
rect 3950 17950 4040 18190
rect 4280 17950 4370 18190
rect 4610 17950 4700 18190
rect 4940 17950 5030 18190
rect 5270 17950 5360 18190
rect 5600 17950 5690 18190
rect 5930 17950 6020 18190
rect 6260 17950 6350 18190
rect 6590 17950 6730 18190
rect -5510 17860 6730 17950
rect -5510 17620 -5200 17860
rect -4960 17620 -4870 17860
rect -4630 17620 -4540 17860
rect -4300 17620 -4210 17860
rect -3970 17620 -3880 17860
rect -3640 17620 -3550 17860
rect -3310 17620 -3220 17860
rect -2980 17620 -2890 17860
rect -2650 17620 -2560 17860
rect -2320 17620 -2230 17860
rect -1990 17620 -1900 17860
rect -1660 17620 -1570 17860
rect -1330 17620 -1240 17860
rect -1000 17620 -910 17860
rect -670 17620 -580 17860
rect -340 17620 -250 17860
rect -10 17620 80 17860
rect 320 17620 410 17860
rect 650 17620 740 17860
rect 980 17620 1070 17860
rect 1310 17620 1400 17860
rect 1640 17620 1730 17860
rect 1970 17620 2060 17860
rect 2300 17620 2390 17860
rect 2630 17620 2720 17860
rect 2960 17620 3050 17860
rect 3290 17620 3380 17860
rect 3620 17620 3710 17860
rect 3950 17620 4040 17860
rect 4280 17620 4370 17860
rect 4610 17620 4700 17860
rect 4940 17620 5030 17860
rect 5270 17620 5360 17860
rect 5600 17620 5690 17860
rect 5930 17620 6020 17860
rect 6260 17620 6350 17860
rect 6590 17620 6730 17860
rect -5510 17530 6730 17620
rect -5510 17290 -5200 17530
rect -4960 17290 -4870 17530
rect -4630 17290 -4540 17530
rect -4300 17290 -4210 17530
rect -3970 17290 -3880 17530
rect -3640 17290 -3550 17530
rect -3310 17290 -3220 17530
rect -2980 17290 -2890 17530
rect -2650 17290 -2560 17530
rect -2320 17290 -2230 17530
rect -1990 17290 -1900 17530
rect -1660 17290 -1570 17530
rect -1330 17290 -1240 17530
rect -1000 17290 -910 17530
rect -670 17290 -580 17530
rect -340 17290 -250 17530
rect -10 17290 80 17530
rect 320 17290 410 17530
rect 650 17290 740 17530
rect 980 17290 1070 17530
rect 1310 17290 1400 17530
rect 1640 17290 1730 17530
rect 1970 17290 2060 17530
rect 2300 17290 2390 17530
rect 2630 17290 2720 17530
rect 2960 17290 3050 17530
rect 3290 17290 3380 17530
rect 3620 17290 3710 17530
rect 3950 17290 4040 17530
rect 4280 17290 4370 17530
rect 4610 17290 4700 17530
rect 4940 17290 5030 17530
rect 5270 17290 5360 17530
rect 5600 17290 5690 17530
rect 5930 17290 6020 17530
rect 6260 17290 6350 17530
rect 6590 17290 6730 17530
rect -5510 17200 6730 17290
rect -5510 16960 -5200 17200
rect -4960 16960 -4870 17200
rect -4630 16960 -4540 17200
rect -4300 16960 -4210 17200
rect -3970 16960 -3880 17200
rect -3640 16960 -3550 17200
rect -3310 16960 -3220 17200
rect -2980 16960 -2890 17200
rect -2650 16960 -2560 17200
rect -2320 16960 -2230 17200
rect -1990 16960 -1900 17200
rect -1660 16960 -1570 17200
rect -1330 16960 -1240 17200
rect -1000 16960 -910 17200
rect -670 16960 -580 17200
rect -340 16960 -250 17200
rect -10 16960 80 17200
rect 320 16960 410 17200
rect 650 16960 740 17200
rect 980 16960 1070 17200
rect 1310 16960 1400 17200
rect 1640 16960 1730 17200
rect 1970 16960 2060 17200
rect 2300 16960 2390 17200
rect 2630 16960 2720 17200
rect 2960 16960 3050 17200
rect 3290 16960 3380 17200
rect 3620 16960 3710 17200
rect 3950 16960 4040 17200
rect 4280 16960 4370 17200
rect 4610 16960 4700 17200
rect 4940 16960 5030 17200
rect 5270 16960 5360 17200
rect 5600 16960 5690 17200
rect 5930 16960 6020 17200
rect 6260 16960 6350 17200
rect 6590 16960 6730 17200
rect -5510 16870 6730 16960
rect -5510 16630 -5200 16870
rect -4960 16630 -4870 16870
rect -4630 16630 -4540 16870
rect -4300 16630 -4210 16870
rect -3970 16630 -3880 16870
rect -3640 16630 -3550 16870
rect -3310 16630 -3220 16870
rect -2980 16630 -2890 16870
rect -2650 16630 -2560 16870
rect -2320 16630 -2230 16870
rect -1990 16630 -1900 16870
rect -1660 16630 -1570 16870
rect -1330 16630 -1240 16870
rect -1000 16630 -910 16870
rect -670 16630 -580 16870
rect -340 16630 -250 16870
rect -10 16630 80 16870
rect 320 16630 410 16870
rect 650 16630 740 16870
rect 980 16630 1070 16870
rect 1310 16630 1400 16870
rect 1640 16630 1730 16870
rect 1970 16630 2060 16870
rect 2300 16630 2390 16870
rect 2630 16630 2720 16870
rect 2960 16630 3050 16870
rect 3290 16630 3380 16870
rect 3620 16630 3710 16870
rect 3950 16630 4040 16870
rect 4280 16630 4370 16870
rect 4610 16630 4700 16870
rect 4940 16630 5030 16870
rect 5270 16630 5360 16870
rect 5600 16630 5690 16870
rect 5930 16630 6020 16870
rect 6260 16630 6350 16870
rect 6590 16630 6730 16870
rect -5510 16540 6730 16630
rect -5510 16300 -5200 16540
rect -4960 16300 -4870 16540
rect -4630 16300 -4540 16540
rect -4300 16300 -4210 16540
rect -3970 16300 -3880 16540
rect -3640 16300 -3550 16540
rect -3310 16300 -3220 16540
rect -2980 16300 -2890 16540
rect -2650 16300 -2560 16540
rect -2320 16300 -2230 16540
rect -1990 16300 -1900 16540
rect -1660 16300 -1570 16540
rect -1330 16300 -1240 16540
rect -1000 16300 -910 16540
rect -670 16300 -580 16540
rect -340 16300 -250 16540
rect -10 16300 80 16540
rect 320 16300 410 16540
rect 650 16300 740 16540
rect 980 16300 1070 16540
rect 1310 16300 1400 16540
rect 1640 16300 1730 16540
rect 1970 16300 2060 16540
rect 2300 16300 2390 16540
rect 2630 16300 2720 16540
rect 2960 16300 3050 16540
rect 3290 16300 3380 16540
rect 3620 16300 3710 16540
rect 3950 16300 4040 16540
rect 4280 16300 4370 16540
rect 4610 16300 4700 16540
rect 4940 16300 5030 16540
rect 5270 16300 5360 16540
rect 5600 16300 5690 16540
rect 5930 16300 6020 16540
rect 6260 16300 6350 16540
rect 6590 16300 6730 16540
rect -5510 16210 6730 16300
rect -5510 15970 -5200 16210
rect -4960 15970 -4870 16210
rect -4630 15970 -4540 16210
rect -4300 15970 -4210 16210
rect -3970 15970 -3880 16210
rect -3640 15970 -3550 16210
rect -3310 15970 -3220 16210
rect -2980 15970 -2890 16210
rect -2650 15970 -2560 16210
rect -2320 15970 -2230 16210
rect -1990 15970 -1900 16210
rect -1660 15970 -1570 16210
rect -1330 15970 -1240 16210
rect -1000 15970 -910 16210
rect -670 15970 -580 16210
rect -340 15970 -250 16210
rect -10 15970 80 16210
rect 320 15970 410 16210
rect 650 15970 740 16210
rect 980 15970 1070 16210
rect 1310 15970 1400 16210
rect 1640 15970 1730 16210
rect 1970 15970 2060 16210
rect 2300 15970 2390 16210
rect 2630 15970 2720 16210
rect 2960 15970 3050 16210
rect 3290 15970 3380 16210
rect 3620 15970 3710 16210
rect 3950 15970 4040 16210
rect 4280 15970 4370 16210
rect 4610 15970 4700 16210
rect 4940 15970 5030 16210
rect 5270 15970 5360 16210
rect 5600 15970 5690 16210
rect 5930 15970 6020 16210
rect 6260 15970 6350 16210
rect 6590 15970 6730 16210
rect -5510 15880 6730 15970
rect -5510 15640 -5200 15880
rect -4960 15640 -4870 15880
rect -4630 15640 -4540 15880
rect -4300 15640 -4210 15880
rect -3970 15640 -3880 15880
rect -3640 15640 -3550 15880
rect -3310 15640 -3220 15880
rect -2980 15640 -2890 15880
rect -2650 15640 -2560 15880
rect -2320 15640 -2230 15880
rect -1990 15640 -1900 15880
rect -1660 15640 -1570 15880
rect -1330 15640 -1240 15880
rect -1000 15640 -910 15880
rect -670 15640 -580 15880
rect -340 15640 -250 15880
rect -10 15640 80 15880
rect 320 15640 410 15880
rect 650 15640 740 15880
rect 980 15640 1070 15880
rect 1310 15640 1400 15880
rect 1640 15640 1730 15880
rect 1970 15640 2060 15880
rect 2300 15640 2390 15880
rect 2630 15640 2720 15880
rect 2960 15640 3050 15880
rect 3290 15640 3380 15880
rect 3620 15640 3710 15880
rect 3950 15640 4040 15880
rect 4280 15640 4370 15880
rect 4610 15640 4700 15880
rect 4940 15640 5030 15880
rect 5270 15640 5360 15880
rect 5600 15640 5690 15880
rect 5930 15640 6020 15880
rect 6260 15640 6350 15880
rect 6590 15640 6730 15880
rect -5510 15550 6730 15640
rect -5510 15310 -5200 15550
rect -4960 15310 -4870 15550
rect -4630 15310 -4540 15550
rect -4300 15310 -4210 15550
rect -3970 15310 -3880 15550
rect -3640 15310 -3550 15550
rect -3310 15310 -3220 15550
rect -2980 15310 -2890 15550
rect -2650 15310 -2560 15550
rect -2320 15310 -2230 15550
rect -1990 15310 -1900 15550
rect -1660 15310 -1570 15550
rect -1330 15310 -1240 15550
rect -1000 15310 -910 15550
rect -670 15310 -580 15550
rect -340 15310 -250 15550
rect -10 15310 80 15550
rect 320 15310 410 15550
rect 650 15310 740 15550
rect 980 15310 1070 15550
rect 1310 15310 1400 15550
rect 1640 15310 1730 15550
rect 1970 15310 2060 15550
rect 2300 15310 2390 15550
rect 2630 15310 2720 15550
rect 2960 15310 3050 15550
rect 3290 15310 3380 15550
rect 3620 15310 3710 15550
rect 3950 15310 4040 15550
rect 4280 15310 4370 15550
rect 4610 15310 4700 15550
rect 4940 15310 5030 15550
rect 5270 15310 5360 15550
rect 5600 15310 5690 15550
rect 5930 15310 6020 15550
rect 6260 15310 6350 15550
rect 6590 15310 6730 15550
rect -5510 15220 6730 15310
rect -5510 14980 -5200 15220
rect -4960 14980 -4870 15220
rect -4630 14980 -4540 15220
rect -4300 14980 -4210 15220
rect -3970 14980 -3880 15220
rect -3640 14980 -3550 15220
rect -3310 14980 -3220 15220
rect -2980 14980 -2890 15220
rect -2650 14980 -2560 15220
rect -2320 14980 -2230 15220
rect -1990 14980 -1900 15220
rect -1660 14980 -1570 15220
rect -1330 14980 -1240 15220
rect -1000 14980 -910 15220
rect -670 14980 -580 15220
rect -340 14980 -250 15220
rect -10 14980 80 15220
rect 320 14980 410 15220
rect 650 14980 740 15220
rect 980 14980 1070 15220
rect 1310 14980 1400 15220
rect 1640 14980 1730 15220
rect 1970 14980 2060 15220
rect 2300 14980 2390 15220
rect 2630 14980 2720 15220
rect 2960 14980 3050 15220
rect 3290 14980 3380 15220
rect 3620 14980 3710 15220
rect 3950 14980 4040 15220
rect 4280 14980 4370 15220
rect 4610 14980 4700 15220
rect 4940 14980 5030 15220
rect 5270 14980 5360 15220
rect 5600 14980 5690 15220
rect 5930 14980 6020 15220
rect 6260 14980 6350 15220
rect 6590 14980 6730 15220
rect -5510 14890 6730 14980
rect -5510 14650 -5200 14890
rect -4960 14650 -4870 14890
rect -4630 14650 -4540 14890
rect -4300 14650 -4210 14890
rect -3970 14650 -3880 14890
rect -3640 14650 -3550 14890
rect -3310 14650 -3220 14890
rect -2980 14650 -2890 14890
rect -2650 14650 -2560 14890
rect -2320 14650 -2230 14890
rect -1990 14650 -1900 14890
rect -1660 14650 -1570 14890
rect -1330 14650 -1240 14890
rect -1000 14650 -910 14890
rect -670 14650 -580 14890
rect -340 14650 -250 14890
rect -10 14650 80 14890
rect 320 14650 410 14890
rect 650 14650 740 14890
rect 980 14650 1070 14890
rect 1310 14650 1400 14890
rect 1640 14650 1730 14890
rect 1970 14650 2060 14890
rect 2300 14650 2390 14890
rect 2630 14650 2720 14890
rect 2960 14650 3050 14890
rect 3290 14650 3380 14890
rect 3620 14650 3710 14890
rect 3950 14650 4040 14890
rect 4280 14650 4370 14890
rect 4610 14650 4700 14890
rect 4940 14650 5030 14890
rect 5270 14650 5360 14890
rect 5600 14650 5690 14890
rect 5930 14650 6020 14890
rect 6260 14650 6350 14890
rect 6590 14650 6730 14890
rect -5510 14560 6730 14650
rect -5510 14320 -5200 14560
rect -4960 14320 -4870 14560
rect -4630 14320 -4540 14560
rect -4300 14320 -4210 14560
rect -3970 14320 -3880 14560
rect -3640 14320 -3550 14560
rect -3310 14320 -3220 14560
rect -2980 14320 -2890 14560
rect -2650 14320 -2560 14560
rect -2320 14320 -2230 14560
rect -1990 14320 -1900 14560
rect -1660 14320 -1570 14560
rect -1330 14320 -1240 14560
rect -1000 14320 -910 14560
rect -670 14320 -580 14560
rect -340 14320 -250 14560
rect -10 14320 80 14560
rect 320 14320 410 14560
rect 650 14320 740 14560
rect 980 14320 1070 14560
rect 1310 14320 1400 14560
rect 1640 14320 1730 14560
rect 1970 14320 2060 14560
rect 2300 14320 2390 14560
rect 2630 14320 2720 14560
rect 2960 14320 3050 14560
rect 3290 14320 3380 14560
rect 3620 14320 3710 14560
rect 3950 14320 4040 14560
rect 4280 14320 4370 14560
rect 4610 14320 4700 14560
rect 4940 14320 5030 14560
rect 5270 14320 5360 14560
rect 5600 14320 5690 14560
rect 5930 14320 6020 14560
rect 6260 14320 6350 14560
rect 6590 14320 6730 14560
rect -5510 14230 6730 14320
rect -5510 13990 -5200 14230
rect -4960 13990 -4870 14230
rect -4630 13990 -4540 14230
rect -4300 13990 -4210 14230
rect -3970 13990 -3880 14230
rect -3640 13990 -3550 14230
rect -3310 13990 -3220 14230
rect -2980 13990 -2890 14230
rect -2650 13990 -2560 14230
rect -2320 13990 -2230 14230
rect -1990 13990 -1900 14230
rect -1660 13990 -1570 14230
rect -1330 13990 -1240 14230
rect -1000 13990 -910 14230
rect -670 13990 -580 14230
rect -340 13990 -250 14230
rect -10 13990 80 14230
rect 320 13990 410 14230
rect 650 13990 740 14230
rect 980 13990 1070 14230
rect 1310 13990 1400 14230
rect 1640 13990 1730 14230
rect 1970 13990 2060 14230
rect 2300 13990 2390 14230
rect 2630 13990 2720 14230
rect 2960 13990 3050 14230
rect 3290 13990 3380 14230
rect 3620 13990 3710 14230
rect 3950 13990 4040 14230
rect 4280 13990 4370 14230
rect 4610 13990 4700 14230
rect 4940 13990 5030 14230
rect 5270 13990 5360 14230
rect 5600 13990 5690 14230
rect 5930 13990 6020 14230
rect 6260 13990 6350 14230
rect 6590 13990 6730 14230
rect -5510 13900 6730 13990
rect -5510 13660 -5200 13900
rect -4960 13660 -4870 13900
rect -4630 13660 -4540 13900
rect -4300 13660 -4210 13900
rect -3970 13660 -3880 13900
rect -3640 13660 -3550 13900
rect -3310 13660 -3220 13900
rect -2980 13660 -2890 13900
rect -2650 13660 -2560 13900
rect -2320 13660 -2230 13900
rect -1990 13660 -1900 13900
rect -1660 13660 -1570 13900
rect -1330 13660 -1240 13900
rect -1000 13660 -910 13900
rect -670 13660 -580 13900
rect -340 13660 -250 13900
rect -10 13660 80 13900
rect 320 13660 410 13900
rect 650 13660 740 13900
rect 980 13660 1070 13900
rect 1310 13660 1400 13900
rect 1640 13660 1730 13900
rect 1970 13660 2060 13900
rect 2300 13660 2390 13900
rect 2630 13660 2720 13900
rect 2960 13660 3050 13900
rect 3290 13660 3380 13900
rect 3620 13660 3710 13900
rect 3950 13660 4040 13900
rect 4280 13660 4370 13900
rect 4610 13660 4700 13900
rect 4940 13660 5030 13900
rect 5270 13660 5360 13900
rect 5600 13660 5690 13900
rect 5930 13660 6020 13900
rect 6260 13660 6350 13900
rect 6590 13660 6730 13900
rect -5510 13570 6730 13660
rect -5510 13330 -5200 13570
rect -4960 13330 -4870 13570
rect -4630 13330 -4540 13570
rect -4300 13330 -4210 13570
rect -3970 13330 -3880 13570
rect -3640 13330 -3550 13570
rect -3310 13330 -3220 13570
rect -2980 13330 -2890 13570
rect -2650 13330 -2560 13570
rect -2320 13330 -2230 13570
rect -1990 13330 -1900 13570
rect -1660 13330 -1570 13570
rect -1330 13330 -1240 13570
rect -1000 13330 -910 13570
rect -670 13330 -580 13570
rect -340 13330 -250 13570
rect -10 13330 80 13570
rect 320 13330 410 13570
rect 650 13330 740 13570
rect 980 13330 1070 13570
rect 1310 13330 1400 13570
rect 1640 13330 1730 13570
rect 1970 13330 2060 13570
rect 2300 13330 2390 13570
rect 2630 13330 2720 13570
rect 2960 13330 3050 13570
rect 3290 13330 3380 13570
rect 3620 13330 3710 13570
rect 3950 13330 4040 13570
rect 4280 13330 4370 13570
rect 4610 13330 4700 13570
rect 4940 13330 5030 13570
rect 5270 13330 5360 13570
rect 5600 13330 5690 13570
rect 5930 13330 6020 13570
rect 6260 13330 6350 13570
rect 6590 13330 6730 13570
rect -5510 13240 6730 13330
rect -5510 13000 -5200 13240
rect -4960 13000 -4870 13240
rect -4630 13000 -4540 13240
rect -4300 13000 -4210 13240
rect -3970 13000 -3880 13240
rect -3640 13000 -3550 13240
rect -3310 13000 -3220 13240
rect -2980 13000 -2890 13240
rect -2650 13000 -2560 13240
rect -2320 13000 -2230 13240
rect -1990 13000 -1900 13240
rect -1660 13000 -1570 13240
rect -1330 13000 -1240 13240
rect -1000 13000 -910 13240
rect -670 13000 -580 13240
rect -340 13000 -250 13240
rect -10 13000 80 13240
rect 320 13000 410 13240
rect 650 13000 740 13240
rect 980 13000 1070 13240
rect 1310 13000 1400 13240
rect 1640 13000 1730 13240
rect 1970 13000 2060 13240
rect 2300 13000 2390 13240
rect 2630 13000 2720 13240
rect 2960 13000 3050 13240
rect 3290 13000 3380 13240
rect 3620 13000 3710 13240
rect 3950 13000 4040 13240
rect 4280 13000 4370 13240
rect 4610 13000 4700 13240
rect 4940 13000 5030 13240
rect 5270 13000 5360 13240
rect 5600 13000 5690 13240
rect 5930 13000 6020 13240
rect 6260 13000 6350 13240
rect 6590 13000 6730 13240
rect -5510 12910 6730 13000
rect -5510 12670 -5200 12910
rect -4960 12670 -4870 12910
rect -4630 12670 -4540 12910
rect -4300 12670 -4210 12910
rect -3970 12670 -3880 12910
rect -3640 12670 -3550 12910
rect -3310 12670 -3220 12910
rect -2980 12670 -2890 12910
rect -2650 12670 -2560 12910
rect -2320 12670 -2230 12910
rect -1990 12670 -1900 12910
rect -1660 12670 -1570 12910
rect -1330 12670 -1240 12910
rect -1000 12670 -910 12910
rect -670 12670 -580 12910
rect -340 12670 -250 12910
rect -10 12670 80 12910
rect 320 12670 410 12910
rect 650 12670 740 12910
rect 980 12670 1070 12910
rect 1310 12670 1400 12910
rect 1640 12670 1730 12910
rect 1970 12670 2060 12910
rect 2300 12670 2390 12910
rect 2630 12670 2720 12910
rect 2960 12670 3050 12910
rect 3290 12670 3380 12910
rect 3620 12670 3710 12910
rect 3950 12670 4040 12910
rect 4280 12670 4370 12910
rect 4610 12670 4700 12910
rect 4940 12670 5030 12910
rect 5270 12670 5360 12910
rect 5600 12670 5690 12910
rect 5930 12670 6020 12910
rect 6260 12670 6350 12910
rect 6590 12670 6730 12910
rect -5510 12580 6730 12670
rect -5510 12340 -5200 12580
rect -4960 12340 -4870 12580
rect -4630 12340 -4540 12580
rect -4300 12340 -4210 12580
rect -3970 12340 -3880 12580
rect -3640 12340 -3550 12580
rect -3310 12340 -3220 12580
rect -2980 12340 -2890 12580
rect -2650 12340 -2560 12580
rect -2320 12340 -2230 12580
rect -1990 12340 -1900 12580
rect -1660 12340 -1570 12580
rect -1330 12340 -1240 12580
rect -1000 12340 -910 12580
rect -670 12340 -580 12580
rect -340 12340 -250 12580
rect -10 12340 80 12580
rect 320 12340 410 12580
rect 650 12340 740 12580
rect 980 12340 1070 12580
rect 1310 12340 1400 12580
rect 1640 12340 1730 12580
rect 1970 12340 2060 12580
rect 2300 12340 2390 12580
rect 2630 12340 2720 12580
rect 2960 12340 3050 12580
rect 3290 12340 3380 12580
rect 3620 12340 3710 12580
rect 3950 12340 4040 12580
rect 4280 12340 4370 12580
rect 4610 12340 4700 12580
rect 4940 12340 5030 12580
rect 5270 12340 5360 12580
rect 5600 12340 5690 12580
rect 5930 12340 6020 12580
rect 6260 12340 6350 12580
rect 6590 12340 6730 12580
rect -5510 12250 6730 12340
rect -5510 12010 -5200 12250
rect -4960 12010 -4870 12250
rect -4630 12010 -4540 12250
rect -4300 12010 -4210 12250
rect -3970 12010 -3880 12250
rect -3640 12010 -3550 12250
rect -3310 12010 -3220 12250
rect -2980 12010 -2890 12250
rect -2650 12010 -2560 12250
rect -2320 12010 -2230 12250
rect -1990 12010 -1900 12250
rect -1660 12010 -1570 12250
rect -1330 12010 -1240 12250
rect -1000 12010 -910 12250
rect -670 12010 -580 12250
rect -340 12010 -250 12250
rect -10 12010 80 12250
rect 320 12010 410 12250
rect 650 12010 740 12250
rect 980 12010 1070 12250
rect 1310 12010 1400 12250
rect 1640 12010 1730 12250
rect 1970 12010 2060 12250
rect 2300 12010 2390 12250
rect 2630 12010 2720 12250
rect 2960 12010 3050 12250
rect 3290 12010 3380 12250
rect 3620 12010 3710 12250
rect 3950 12010 4040 12250
rect 4280 12010 4370 12250
rect 4610 12010 4700 12250
rect 4940 12010 5030 12250
rect 5270 12010 5360 12250
rect 5600 12010 5690 12250
rect 5930 12010 6020 12250
rect 6260 12010 6350 12250
rect 6590 12010 6730 12250
rect -5510 11920 6730 12010
rect -5510 11680 -5200 11920
rect -4960 11680 -4870 11920
rect -4630 11680 -4540 11920
rect -4300 11680 -4210 11920
rect -3970 11680 -3880 11920
rect -3640 11680 -3550 11920
rect -3310 11680 -3220 11920
rect -2980 11680 -2890 11920
rect -2650 11680 -2560 11920
rect -2320 11680 -2230 11920
rect -1990 11680 -1900 11920
rect -1660 11680 -1570 11920
rect -1330 11680 -1240 11920
rect -1000 11680 -910 11920
rect -670 11680 -580 11920
rect -340 11680 -250 11920
rect -10 11680 80 11920
rect 320 11680 410 11920
rect 650 11680 740 11920
rect 980 11680 1070 11920
rect 1310 11680 1400 11920
rect 1640 11680 1730 11920
rect 1970 11680 2060 11920
rect 2300 11680 2390 11920
rect 2630 11680 2720 11920
rect 2960 11680 3050 11920
rect 3290 11680 3380 11920
rect 3620 11680 3710 11920
rect 3950 11680 4040 11920
rect 4280 11680 4370 11920
rect 4610 11680 4700 11920
rect 4940 11680 5030 11920
rect 5270 11680 5360 11920
rect 5600 11680 5690 11920
rect 5930 11680 6020 11920
rect 6260 11680 6350 11920
rect 6590 11680 6730 11920
rect -5510 11590 6730 11680
rect -5510 11350 -5200 11590
rect -4960 11350 -4870 11590
rect -4630 11350 -4540 11590
rect -4300 11350 -4210 11590
rect -3970 11350 -3880 11590
rect -3640 11350 -3550 11590
rect -3310 11350 -3220 11590
rect -2980 11350 -2890 11590
rect -2650 11350 -2560 11590
rect -2320 11350 -2230 11590
rect -1990 11350 -1900 11590
rect -1660 11350 -1570 11590
rect -1330 11350 -1240 11590
rect -1000 11350 -910 11590
rect -670 11350 -580 11590
rect -340 11350 -250 11590
rect -10 11350 80 11590
rect 320 11350 410 11590
rect 650 11350 740 11590
rect 980 11350 1070 11590
rect 1310 11350 1400 11590
rect 1640 11350 1730 11590
rect 1970 11350 2060 11590
rect 2300 11350 2390 11590
rect 2630 11350 2720 11590
rect 2960 11350 3050 11590
rect 3290 11350 3380 11590
rect 3620 11350 3710 11590
rect 3950 11350 4040 11590
rect 4280 11350 4370 11590
rect 4610 11350 4700 11590
rect 4940 11350 5030 11590
rect 5270 11350 5360 11590
rect 5600 11350 5690 11590
rect 5930 11350 6020 11590
rect 6260 11350 6350 11590
rect 6590 11350 6730 11590
rect -5510 11260 6730 11350
rect -5510 11020 -5200 11260
rect -4960 11020 -4870 11260
rect -4630 11020 -4540 11260
rect -4300 11020 -4210 11260
rect -3970 11020 -3880 11260
rect -3640 11020 -3550 11260
rect -3310 11020 -3220 11260
rect -2980 11020 -2890 11260
rect -2650 11020 -2560 11260
rect -2320 11020 -2230 11260
rect -1990 11020 -1900 11260
rect -1660 11020 -1570 11260
rect -1330 11020 -1240 11260
rect -1000 11020 -910 11260
rect -670 11020 -580 11260
rect -340 11020 -250 11260
rect -10 11020 80 11260
rect 320 11020 410 11260
rect 650 11020 740 11260
rect 980 11020 1070 11260
rect 1310 11020 1400 11260
rect 1640 11020 1730 11260
rect 1970 11020 2060 11260
rect 2300 11020 2390 11260
rect 2630 11020 2720 11260
rect 2960 11020 3050 11260
rect 3290 11020 3380 11260
rect 3620 11020 3710 11260
rect 3950 11020 4040 11260
rect 4280 11020 4370 11260
rect 4610 11020 4700 11260
rect 4940 11020 5030 11260
rect 5270 11020 5360 11260
rect 5600 11020 5690 11260
rect 5930 11020 6020 11260
rect 6260 11020 6350 11260
rect 6590 11020 6730 11260
rect -5510 10930 6730 11020
rect -5510 10690 -5200 10930
rect -4960 10690 -4870 10930
rect -4630 10690 -4540 10930
rect -4300 10690 -4210 10930
rect -3970 10690 -3880 10930
rect -3640 10690 -3550 10930
rect -3310 10690 -3220 10930
rect -2980 10690 -2890 10930
rect -2650 10690 -2560 10930
rect -2320 10690 -2230 10930
rect -1990 10690 -1900 10930
rect -1660 10690 -1570 10930
rect -1330 10690 -1240 10930
rect -1000 10690 -910 10930
rect -670 10690 -580 10930
rect -340 10690 -250 10930
rect -10 10690 80 10930
rect 320 10690 410 10930
rect 650 10690 740 10930
rect 980 10690 1070 10930
rect 1310 10690 1400 10930
rect 1640 10690 1730 10930
rect 1970 10690 2060 10930
rect 2300 10690 2390 10930
rect 2630 10690 2720 10930
rect 2960 10690 3050 10930
rect 3290 10690 3380 10930
rect 3620 10690 3710 10930
rect 3950 10690 4040 10930
rect 4280 10690 4370 10930
rect 4610 10690 4700 10930
rect 4940 10690 5030 10930
rect 5270 10690 5360 10930
rect 5600 10690 5690 10930
rect 5930 10690 6020 10930
rect 6260 10690 6350 10930
rect 6590 10690 6730 10930
rect -5510 10600 6730 10690
rect -5510 10360 -5200 10600
rect -4960 10360 -4870 10600
rect -4630 10360 -4540 10600
rect -4300 10360 -4210 10600
rect -3970 10360 -3880 10600
rect -3640 10360 -3550 10600
rect -3310 10360 -3220 10600
rect -2980 10360 -2890 10600
rect -2650 10360 -2560 10600
rect -2320 10360 -2230 10600
rect -1990 10360 -1900 10600
rect -1660 10360 -1570 10600
rect -1330 10360 -1240 10600
rect -1000 10360 -910 10600
rect -670 10360 -580 10600
rect -340 10360 -250 10600
rect -10 10360 80 10600
rect 320 10360 410 10600
rect 650 10360 740 10600
rect 980 10360 1070 10600
rect 1310 10360 1400 10600
rect 1640 10360 1730 10600
rect 1970 10360 2060 10600
rect 2300 10360 2390 10600
rect 2630 10360 2720 10600
rect 2960 10360 3050 10600
rect 3290 10360 3380 10600
rect 3620 10360 3710 10600
rect 3950 10360 4040 10600
rect 4280 10360 4370 10600
rect 4610 10360 4700 10600
rect 4940 10360 5030 10600
rect 5270 10360 5360 10600
rect 5600 10360 5690 10600
rect 5930 10360 6020 10600
rect 6260 10360 6350 10600
rect 6590 10360 6730 10600
rect -5510 10270 6730 10360
rect -5510 10030 -5200 10270
rect -4960 10030 -4870 10270
rect -4630 10030 -4540 10270
rect -4300 10030 -4210 10270
rect -3970 10030 -3880 10270
rect -3640 10030 -3550 10270
rect -3310 10030 -3220 10270
rect -2980 10030 -2890 10270
rect -2650 10030 -2560 10270
rect -2320 10030 -2230 10270
rect -1990 10030 -1900 10270
rect -1660 10030 -1570 10270
rect -1330 10030 -1240 10270
rect -1000 10030 -910 10270
rect -670 10030 -580 10270
rect -340 10030 -250 10270
rect -10 10030 80 10270
rect 320 10030 410 10270
rect 650 10030 740 10270
rect 980 10030 1070 10270
rect 1310 10030 1400 10270
rect 1640 10030 1730 10270
rect 1970 10030 2060 10270
rect 2300 10030 2390 10270
rect 2630 10030 2720 10270
rect 2960 10030 3050 10270
rect 3290 10030 3380 10270
rect 3620 10030 3710 10270
rect 3950 10030 4040 10270
rect 4280 10030 4370 10270
rect 4610 10030 4700 10270
rect 4940 10030 5030 10270
rect 5270 10030 5360 10270
rect 5600 10030 5690 10270
rect 5930 10030 6020 10270
rect 6260 10030 6350 10270
rect 6590 10030 6730 10270
rect -5510 9940 6730 10030
rect -5510 9700 -5200 9940
rect -4960 9700 -4870 9940
rect -4630 9700 -4540 9940
rect -4300 9700 -4210 9940
rect -3970 9700 -3880 9940
rect -3640 9700 -3550 9940
rect -3310 9700 -3220 9940
rect -2980 9700 -2890 9940
rect -2650 9700 -2560 9940
rect -2320 9700 -2230 9940
rect -1990 9700 -1900 9940
rect -1660 9700 -1570 9940
rect -1330 9700 -1240 9940
rect -1000 9700 -910 9940
rect -670 9700 -580 9940
rect -340 9700 -250 9940
rect -10 9700 80 9940
rect 320 9700 410 9940
rect 650 9700 740 9940
rect 980 9700 1070 9940
rect 1310 9700 1400 9940
rect 1640 9700 1730 9940
rect 1970 9700 2060 9940
rect 2300 9700 2390 9940
rect 2630 9700 2720 9940
rect 2960 9700 3050 9940
rect 3290 9700 3380 9940
rect 3620 9700 3710 9940
rect 3950 9700 4040 9940
rect 4280 9700 4370 9940
rect 4610 9700 4700 9940
rect 4940 9700 5030 9940
rect 5270 9700 5360 9940
rect 5600 9700 5690 9940
rect 5930 9700 6020 9940
rect 6260 9700 6350 9940
rect 6590 9700 6730 9940
rect -5510 9610 6730 9700
rect -5510 9370 -5200 9610
rect -4960 9370 -4870 9610
rect -4630 9370 -4540 9610
rect -4300 9370 -4210 9610
rect -3970 9370 -3880 9610
rect -3640 9370 -3550 9610
rect -3310 9370 -3220 9610
rect -2980 9370 -2890 9610
rect -2650 9370 -2560 9610
rect -2320 9370 -2230 9610
rect -1990 9370 -1900 9610
rect -1660 9370 -1570 9610
rect -1330 9370 -1240 9610
rect -1000 9370 -910 9610
rect -670 9370 -580 9610
rect -340 9370 -250 9610
rect -10 9370 80 9610
rect 320 9370 410 9610
rect 650 9370 740 9610
rect 980 9370 1070 9610
rect 1310 9370 1400 9610
rect 1640 9370 1730 9610
rect 1970 9370 2060 9610
rect 2300 9370 2390 9610
rect 2630 9370 2720 9610
rect 2960 9370 3050 9610
rect 3290 9370 3380 9610
rect 3620 9370 3710 9610
rect 3950 9370 4040 9610
rect 4280 9370 4370 9610
rect 4610 9370 4700 9610
rect 4940 9370 5030 9610
rect 5270 9370 5360 9610
rect 5600 9370 5690 9610
rect 5930 9370 6020 9610
rect 6260 9370 6350 9610
rect 6590 9370 6730 9610
rect -5510 9280 6730 9370
rect -5510 9040 -5200 9280
rect -4960 9040 -4870 9280
rect -4630 9040 -4540 9280
rect -4300 9040 -4210 9280
rect -3970 9040 -3880 9280
rect -3640 9040 -3550 9280
rect -3310 9040 -3220 9280
rect -2980 9040 -2890 9280
rect -2650 9040 -2560 9280
rect -2320 9040 -2230 9280
rect -1990 9040 -1900 9280
rect -1660 9040 -1570 9280
rect -1330 9040 -1240 9280
rect -1000 9040 -910 9280
rect -670 9040 -580 9280
rect -340 9040 -250 9280
rect -10 9040 80 9280
rect 320 9040 410 9280
rect 650 9040 740 9280
rect 980 9040 1070 9280
rect 1310 9040 1400 9280
rect 1640 9040 1730 9280
rect 1970 9040 2060 9280
rect 2300 9040 2390 9280
rect 2630 9040 2720 9280
rect 2960 9040 3050 9280
rect 3290 9040 3380 9280
rect 3620 9040 3710 9280
rect 3950 9040 4040 9280
rect 4280 9040 4370 9280
rect 4610 9040 4700 9280
rect 4940 9040 5030 9280
rect 5270 9040 5360 9280
rect 5600 9040 5690 9280
rect 5930 9040 6020 9280
rect 6260 9040 6350 9280
rect 6590 9040 6730 9280
rect -5510 8720 6730 9040
rect 8170 20830 20410 20960
rect 8170 20590 8310 20830
rect 8550 20590 8640 20830
rect 8880 20590 8970 20830
rect 9210 20590 9300 20830
rect 9540 20590 9630 20830
rect 9870 20590 9960 20830
rect 10200 20590 10290 20830
rect 10530 20590 10620 20830
rect 10860 20590 10950 20830
rect 11190 20590 11280 20830
rect 11520 20590 11610 20830
rect 11850 20590 11940 20830
rect 12180 20590 12270 20830
rect 12510 20590 12600 20830
rect 12840 20590 12930 20830
rect 13170 20590 13260 20830
rect 13500 20590 13590 20830
rect 13830 20590 13920 20830
rect 14160 20590 14250 20830
rect 14490 20590 14580 20830
rect 14820 20590 14910 20830
rect 15150 20590 15240 20830
rect 15480 20590 15570 20830
rect 15810 20590 15900 20830
rect 16140 20590 16230 20830
rect 16470 20590 16560 20830
rect 16800 20590 16890 20830
rect 17130 20590 17220 20830
rect 17460 20590 17550 20830
rect 17790 20590 17880 20830
rect 18120 20590 18210 20830
rect 18450 20590 18540 20830
rect 18780 20590 18870 20830
rect 19110 20590 19200 20830
rect 19440 20590 19530 20830
rect 19770 20590 19860 20830
rect 20100 20590 20410 20830
rect 8170 20500 20410 20590
rect 8170 20260 8310 20500
rect 8550 20260 8640 20500
rect 8880 20260 8970 20500
rect 9210 20260 9300 20500
rect 9540 20260 9630 20500
rect 9870 20260 9960 20500
rect 10200 20260 10290 20500
rect 10530 20260 10620 20500
rect 10860 20260 10950 20500
rect 11190 20260 11280 20500
rect 11520 20260 11610 20500
rect 11850 20260 11940 20500
rect 12180 20260 12270 20500
rect 12510 20260 12600 20500
rect 12840 20260 12930 20500
rect 13170 20260 13260 20500
rect 13500 20260 13590 20500
rect 13830 20260 13920 20500
rect 14160 20260 14250 20500
rect 14490 20260 14580 20500
rect 14820 20260 14910 20500
rect 15150 20260 15240 20500
rect 15480 20260 15570 20500
rect 15810 20260 15900 20500
rect 16140 20260 16230 20500
rect 16470 20260 16560 20500
rect 16800 20260 16890 20500
rect 17130 20260 17220 20500
rect 17460 20260 17550 20500
rect 17790 20260 17880 20500
rect 18120 20260 18210 20500
rect 18450 20260 18540 20500
rect 18780 20260 18870 20500
rect 19110 20260 19200 20500
rect 19440 20260 19530 20500
rect 19770 20260 19860 20500
rect 20100 20260 20410 20500
rect 8170 20170 20410 20260
rect 8170 19930 8310 20170
rect 8550 19930 8640 20170
rect 8880 19930 8970 20170
rect 9210 19930 9300 20170
rect 9540 19930 9630 20170
rect 9870 19930 9960 20170
rect 10200 19930 10290 20170
rect 10530 19930 10620 20170
rect 10860 19930 10950 20170
rect 11190 19930 11280 20170
rect 11520 19930 11610 20170
rect 11850 19930 11940 20170
rect 12180 19930 12270 20170
rect 12510 19930 12600 20170
rect 12840 19930 12930 20170
rect 13170 19930 13260 20170
rect 13500 19930 13590 20170
rect 13830 19930 13920 20170
rect 14160 19930 14250 20170
rect 14490 19930 14580 20170
rect 14820 19930 14910 20170
rect 15150 19930 15240 20170
rect 15480 19930 15570 20170
rect 15810 19930 15900 20170
rect 16140 19930 16230 20170
rect 16470 19930 16560 20170
rect 16800 19930 16890 20170
rect 17130 19930 17220 20170
rect 17460 19930 17550 20170
rect 17790 19930 17880 20170
rect 18120 19930 18210 20170
rect 18450 19930 18540 20170
rect 18780 19930 18870 20170
rect 19110 19930 19200 20170
rect 19440 19930 19530 20170
rect 19770 19930 19860 20170
rect 20100 19930 20410 20170
rect 8170 19840 20410 19930
rect 8170 19600 8310 19840
rect 8550 19600 8640 19840
rect 8880 19600 8970 19840
rect 9210 19600 9300 19840
rect 9540 19600 9630 19840
rect 9870 19600 9960 19840
rect 10200 19600 10290 19840
rect 10530 19600 10620 19840
rect 10860 19600 10950 19840
rect 11190 19600 11280 19840
rect 11520 19600 11610 19840
rect 11850 19600 11940 19840
rect 12180 19600 12270 19840
rect 12510 19600 12600 19840
rect 12840 19600 12930 19840
rect 13170 19600 13260 19840
rect 13500 19600 13590 19840
rect 13830 19600 13920 19840
rect 14160 19600 14250 19840
rect 14490 19600 14580 19840
rect 14820 19600 14910 19840
rect 15150 19600 15240 19840
rect 15480 19600 15570 19840
rect 15810 19600 15900 19840
rect 16140 19600 16230 19840
rect 16470 19600 16560 19840
rect 16800 19600 16890 19840
rect 17130 19600 17220 19840
rect 17460 19600 17550 19840
rect 17790 19600 17880 19840
rect 18120 19600 18210 19840
rect 18450 19600 18540 19840
rect 18780 19600 18870 19840
rect 19110 19600 19200 19840
rect 19440 19600 19530 19840
rect 19770 19600 19860 19840
rect 20100 19600 20410 19840
rect 8170 19510 20410 19600
rect 8170 19270 8310 19510
rect 8550 19270 8640 19510
rect 8880 19270 8970 19510
rect 9210 19270 9300 19510
rect 9540 19270 9630 19510
rect 9870 19270 9960 19510
rect 10200 19270 10290 19510
rect 10530 19270 10620 19510
rect 10860 19270 10950 19510
rect 11190 19270 11280 19510
rect 11520 19270 11610 19510
rect 11850 19270 11940 19510
rect 12180 19270 12270 19510
rect 12510 19270 12600 19510
rect 12840 19270 12930 19510
rect 13170 19270 13260 19510
rect 13500 19270 13590 19510
rect 13830 19270 13920 19510
rect 14160 19270 14250 19510
rect 14490 19270 14580 19510
rect 14820 19270 14910 19510
rect 15150 19270 15240 19510
rect 15480 19270 15570 19510
rect 15810 19270 15900 19510
rect 16140 19270 16230 19510
rect 16470 19270 16560 19510
rect 16800 19270 16890 19510
rect 17130 19270 17220 19510
rect 17460 19270 17550 19510
rect 17790 19270 17880 19510
rect 18120 19270 18210 19510
rect 18450 19270 18540 19510
rect 18780 19270 18870 19510
rect 19110 19270 19200 19510
rect 19440 19270 19530 19510
rect 19770 19270 19860 19510
rect 20100 19270 20410 19510
rect 8170 19180 20410 19270
rect 8170 18940 8310 19180
rect 8550 18940 8640 19180
rect 8880 18940 8970 19180
rect 9210 18940 9300 19180
rect 9540 18940 9630 19180
rect 9870 18940 9960 19180
rect 10200 18940 10290 19180
rect 10530 18940 10620 19180
rect 10860 18940 10950 19180
rect 11190 18940 11280 19180
rect 11520 18940 11610 19180
rect 11850 18940 11940 19180
rect 12180 18940 12270 19180
rect 12510 18940 12600 19180
rect 12840 18940 12930 19180
rect 13170 18940 13260 19180
rect 13500 18940 13590 19180
rect 13830 18940 13920 19180
rect 14160 18940 14250 19180
rect 14490 18940 14580 19180
rect 14820 18940 14910 19180
rect 15150 18940 15240 19180
rect 15480 18940 15570 19180
rect 15810 18940 15900 19180
rect 16140 18940 16230 19180
rect 16470 18940 16560 19180
rect 16800 18940 16890 19180
rect 17130 18940 17220 19180
rect 17460 18940 17550 19180
rect 17790 18940 17880 19180
rect 18120 18940 18210 19180
rect 18450 18940 18540 19180
rect 18780 18940 18870 19180
rect 19110 18940 19200 19180
rect 19440 18940 19530 19180
rect 19770 18940 19860 19180
rect 20100 18940 20410 19180
rect 8170 18850 20410 18940
rect 8170 18610 8310 18850
rect 8550 18610 8640 18850
rect 8880 18610 8970 18850
rect 9210 18610 9300 18850
rect 9540 18610 9630 18850
rect 9870 18610 9960 18850
rect 10200 18610 10290 18850
rect 10530 18610 10620 18850
rect 10860 18610 10950 18850
rect 11190 18610 11280 18850
rect 11520 18610 11610 18850
rect 11850 18610 11940 18850
rect 12180 18610 12270 18850
rect 12510 18610 12600 18850
rect 12840 18610 12930 18850
rect 13170 18610 13260 18850
rect 13500 18610 13590 18850
rect 13830 18610 13920 18850
rect 14160 18610 14250 18850
rect 14490 18610 14580 18850
rect 14820 18610 14910 18850
rect 15150 18610 15240 18850
rect 15480 18610 15570 18850
rect 15810 18610 15900 18850
rect 16140 18610 16230 18850
rect 16470 18610 16560 18850
rect 16800 18610 16890 18850
rect 17130 18610 17220 18850
rect 17460 18610 17550 18850
rect 17790 18610 17880 18850
rect 18120 18610 18210 18850
rect 18450 18610 18540 18850
rect 18780 18610 18870 18850
rect 19110 18610 19200 18850
rect 19440 18610 19530 18850
rect 19770 18610 19860 18850
rect 20100 18610 20410 18850
rect 8170 18520 20410 18610
rect 8170 18280 8310 18520
rect 8550 18280 8640 18520
rect 8880 18280 8970 18520
rect 9210 18280 9300 18520
rect 9540 18280 9630 18520
rect 9870 18280 9960 18520
rect 10200 18280 10290 18520
rect 10530 18280 10620 18520
rect 10860 18280 10950 18520
rect 11190 18280 11280 18520
rect 11520 18280 11610 18520
rect 11850 18280 11940 18520
rect 12180 18280 12270 18520
rect 12510 18280 12600 18520
rect 12840 18280 12930 18520
rect 13170 18280 13260 18520
rect 13500 18280 13590 18520
rect 13830 18280 13920 18520
rect 14160 18280 14250 18520
rect 14490 18280 14580 18520
rect 14820 18280 14910 18520
rect 15150 18280 15240 18520
rect 15480 18280 15570 18520
rect 15810 18280 15900 18520
rect 16140 18280 16230 18520
rect 16470 18280 16560 18520
rect 16800 18280 16890 18520
rect 17130 18280 17220 18520
rect 17460 18280 17550 18520
rect 17790 18280 17880 18520
rect 18120 18280 18210 18520
rect 18450 18280 18540 18520
rect 18780 18280 18870 18520
rect 19110 18280 19200 18520
rect 19440 18280 19530 18520
rect 19770 18280 19860 18520
rect 20100 18280 20410 18520
rect 8170 18190 20410 18280
rect 8170 17950 8310 18190
rect 8550 17950 8640 18190
rect 8880 17950 8970 18190
rect 9210 17950 9300 18190
rect 9540 17950 9630 18190
rect 9870 17950 9960 18190
rect 10200 17950 10290 18190
rect 10530 17950 10620 18190
rect 10860 17950 10950 18190
rect 11190 17950 11280 18190
rect 11520 17950 11610 18190
rect 11850 17950 11940 18190
rect 12180 17950 12270 18190
rect 12510 17950 12600 18190
rect 12840 17950 12930 18190
rect 13170 17950 13260 18190
rect 13500 17950 13590 18190
rect 13830 17950 13920 18190
rect 14160 17950 14250 18190
rect 14490 17950 14580 18190
rect 14820 17950 14910 18190
rect 15150 17950 15240 18190
rect 15480 17950 15570 18190
rect 15810 17950 15900 18190
rect 16140 17950 16230 18190
rect 16470 17950 16560 18190
rect 16800 17950 16890 18190
rect 17130 17950 17220 18190
rect 17460 17950 17550 18190
rect 17790 17950 17880 18190
rect 18120 17950 18210 18190
rect 18450 17950 18540 18190
rect 18780 17950 18870 18190
rect 19110 17950 19200 18190
rect 19440 17950 19530 18190
rect 19770 17950 19860 18190
rect 20100 17950 20410 18190
rect 8170 17860 20410 17950
rect 8170 17620 8310 17860
rect 8550 17620 8640 17860
rect 8880 17620 8970 17860
rect 9210 17620 9300 17860
rect 9540 17620 9630 17860
rect 9870 17620 9960 17860
rect 10200 17620 10290 17860
rect 10530 17620 10620 17860
rect 10860 17620 10950 17860
rect 11190 17620 11280 17860
rect 11520 17620 11610 17860
rect 11850 17620 11940 17860
rect 12180 17620 12270 17860
rect 12510 17620 12600 17860
rect 12840 17620 12930 17860
rect 13170 17620 13260 17860
rect 13500 17620 13590 17860
rect 13830 17620 13920 17860
rect 14160 17620 14250 17860
rect 14490 17620 14580 17860
rect 14820 17620 14910 17860
rect 15150 17620 15240 17860
rect 15480 17620 15570 17860
rect 15810 17620 15900 17860
rect 16140 17620 16230 17860
rect 16470 17620 16560 17860
rect 16800 17620 16890 17860
rect 17130 17620 17220 17860
rect 17460 17620 17550 17860
rect 17790 17620 17880 17860
rect 18120 17620 18210 17860
rect 18450 17620 18540 17860
rect 18780 17620 18870 17860
rect 19110 17620 19200 17860
rect 19440 17620 19530 17860
rect 19770 17620 19860 17860
rect 20100 17620 20410 17860
rect 8170 17530 20410 17620
rect 8170 17290 8310 17530
rect 8550 17290 8640 17530
rect 8880 17290 8970 17530
rect 9210 17290 9300 17530
rect 9540 17290 9630 17530
rect 9870 17290 9960 17530
rect 10200 17290 10290 17530
rect 10530 17290 10620 17530
rect 10860 17290 10950 17530
rect 11190 17290 11280 17530
rect 11520 17290 11610 17530
rect 11850 17290 11940 17530
rect 12180 17290 12270 17530
rect 12510 17290 12600 17530
rect 12840 17290 12930 17530
rect 13170 17290 13260 17530
rect 13500 17290 13590 17530
rect 13830 17290 13920 17530
rect 14160 17290 14250 17530
rect 14490 17290 14580 17530
rect 14820 17290 14910 17530
rect 15150 17290 15240 17530
rect 15480 17290 15570 17530
rect 15810 17290 15900 17530
rect 16140 17290 16230 17530
rect 16470 17290 16560 17530
rect 16800 17290 16890 17530
rect 17130 17290 17220 17530
rect 17460 17290 17550 17530
rect 17790 17290 17880 17530
rect 18120 17290 18210 17530
rect 18450 17290 18540 17530
rect 18780 17290 18870 17530
rect 19110 17290 19200 17530
rect 19440 17290 19530 17530
rect 19770 17290 19860 17530
rect 20100 17290 20410 17530
rect 8170 17200 20410 17290
rect 8170 16960 8310 17200
rect 8550 16960 8640 17200
rect 8880 16960 8970 17200
rect 9210 16960 9300 17200
rect 9540 16960 9630 17200
rect 9870 16960 9960 17200
rect 10200 16960 10290 17200
rect 10530 16960 10620 17200
rect 10860 16960 10950 17200
rect 11190 16960 11280 17200
rect 11520 16960 11610 17200
rect 11850 16960 11940 17200
rect 12180 16960 12270 17200
rect 12510 16960 12600 17200
rect 12840 16960 12930 17200
rect 13170 16960 13260 17200
rect 13500 16960 13590 17200
rect 13830 16960 13920 17200
rect 14160 16960 14250 17200
rect 14490 16960 14580 17200
rect 14820 16960 14910 17200
rect 15150 16960 15240 17200
rect 15480 16960 15570 17200
rect 15810 16960 15900 17200
rect 16140 16960 16230 17200
rect 16470 16960 16560 17200
rect 16800 16960 16890 17200
rect 17130 16960 17220 17200
rect 17460 16960 17550 17200
rect 17790 16960 17880 17200
rect 18120 16960 18210 17200
rect 18450 16960 18540 17200
rect 18780 16960 18870 17200
rect 19110 16960 19200 17200
rect 19440 16960 19530 17200
rect 19770 16960 19860 17200
rect 20100 16960 20410 17200
rect 8170 16870 20410 16960
rect 8170 16630 8310 16870
rect 8550 16630 8640 16870
rect 8880 16630 8970 16870
rect 9210 16630 9300 16870
rect 9540 16630 9630 16870
rect 9870 16630 9960 16870
rect 10200 16630 10290 16870
rect 10530 16630 10620 16870
rect 10860 16630 10950 16870
rect 11190 16630 11280 16870
rect 11520 16630 11610 16870
rect 11850 16630 11940 16870
rect 12180 16630 12270 16870
rect 12510 16630 12600 16870
rect 12840 16630 12930 16870
rect 13170 16630 13260 16870
rect 13500 16630 13590 16870
rect 13830 16630 13920 16870
rect 14160 16630 14250 16870
rect 14490 16630 14580 16870
rect 14820 16630 14910 16870
rect 15150 16630 15240 16870
rect 15480 16630 15570 16870
rect 15810 16630 15900 16870
rect 16140 16630 16230 16870
rect 16470 16630 16560 16870
rect 16800 16630 16890 16870
rect 17130 16630 17220 16870
rect 17460 16630 17550 16870
rect 17790 16630 17880 16870
rect 18120 16630 18210 16870
rect 18450 16630 18540 16870
rect 18780 16630 18870 16870
rect 19110 16630 19200 16870
rect 19440 16630 19530 16870
rect 19770 16630 19860 16870
rect 20100 16630 20410 16870
rect 8170 16540 20410 16630
rect 8170 16300 8310 16540
rect 8550 16300 8640 16540
rect 8880 16300 8970 16540
rect 9210 16300 9300 16540
rect 9540 16300 9630 16540
rect 9870 16300 9960 16540
rect 10200 16300 10290 16540
rect 10530 16300 10620 16540
rect 10860 16300 10950 16540
rect 11190 16300 11280 16540
rect 11520 16300 11610 16540
rect 11850 16300 11940 16540
rect 12180 16300 12270 16540
rect 12510 16300 12600 16540
rect 12840 16300 12930 16540
rect 13170 16300 13260 16540
rect 13500 16300 13590 16540
rect 13830 16300 13920 16540
rect 14160 16300 14250 16540
rect 14490 16300 14580 16540
rect 14820 16300 14910 16540
rect 15150 16300 15240 16540
rect 15480 16300 15570 16540
rect 15810 16300 15900 16540
rect 16140 16300 16230 16540
rect 16470 16300 16560 16540
rect 16800 16300 16890 16540
rect 17130 16300 17220 16540
rect 17460 16300 17550 16540
rect 17790 16300 17880 16540
rect 18120 16300 18210 16540
rect 18450 16300 18540 16540
rect 18780 16300 18870 16540
rect 19110 16300 19200 16540
rect 19440 16300 19530 16540
rect 19770 16300 19860 16540
rect 20100 16300 20410 16540
rect 8170 16210 20410 16300
rect 8170 15970 8310 16210
rect 8550 15970 8640 16210
rect 8880 15970 8970 16210
rect 9210 15970 9300 16210
rect 9540 15970 9630 16210
rect 9870 15970 9960 16210
rect 10200 15970 10290 16210
rect 10530 15970 10620 16210
rect 10860 15970 10950 16210
rect 11190 15970 11280 16210
rect 11520 15970 11610 16210
rect 11850 15970 11940 16210
rect 12180 15970 12270 16210
rect 12510 15970 12600 16210
rect 12840 15970 12930 16210
rect 13170 15970 13260 16210
rect 13500 15970 13590 16210
rect 13830 15970 13920 16210
rect 14160 15970 14250 16210
rect 14490 15970 14580 16210
rect 14820 15970 14910 16210
rect 15150 15970 15240 16210
rect 15480 15970 15570 16210
rect 15810 15970 15900 16210
rect 16140 15970 16230 16210
rect 16470 15970 16560 16210
rect 16800 15970 16890 16210
rect 17130 15970 17220 16210
rect 17460 15970 17550 16210
rect 17790 15970 17880 16210
rect 18120 15970 18210 16210
rect 18450 15970 18540 16210
rect 18780 15970 18870 16210
rect 19110 15970 19200 16210
rect 19440 15970 19530 16210
rect 19770 15970 19860 16210
rect 20100 15970 20410 16210
rect 8170 15880 20410 15970
rect 8170 15640 8310 15880
rect 8550 15640 8640 15880
rect 8880 15640 8970 15880
rect 9210 15640 9300 15880
rect 9540 15640 9630 15880
rect 9870 15640 9960 15880
rect 10200 15640 10290 15880
rect 10530 15640 10620 15880
rect 10860 15640 10950 15880
rect 11190 15640 11280 15880
rect 11520 15640 11610 15880
rect 11850 15640 11940 15880
rect 12180 15640 12270 15880
rect 12510 15640 12600 15880
rect 12840 15640 12930 15880
rect 13170 15640 13260 15880
rect 13500 15640 13590 15880
rect 13830 15640 13920 15880
rect 14160 15640 14250 15880
rect 14490 15640 14580 15880
rect 14820 15640 14910 15880
rect 15150 15640 15240 15880
rect 15480 15640 15570 15880
rect 15810 15640 15900 15880
rect 16140 15640 16230 15880
rect 16470 15640 16560 15880
rect 16800 15640 16890 15880
rect 17130 15640 17220 15880
rect 17460 15640 17550 15880
rect 17790 15640 17880 15880
rect 18120 15640 18210 15880
rect 18450 15640 18540 15880
rect 18780 15640 18870 15880
rect 19110 15640 19200 15880
rect 19440 15640 19530 15880
rect 19770 15640 19860 15880
rect 20100 15640 20410 15880
rect 8170 15550 20410 15640
rect 8170 15310 8310 15550
rect 8550 15310 8640 15550
rect 8880 15310 8970 15550
rect 9210 15310 9300 15550
rect 9540 15310 9630 15550
rect 9870 15310 9960 15550
rect 10200 15310 10290 15550
rect 10530 15310 10620 15550
rect 10860 15310 10950 15550
rect 11190 15310 11280 15550
rect 11520 15310 11610 15550
rect 11850 15310 11940 15550
rect 12180 15310 12270 15550
rect 12510 15310 12600 15550
rect 12840 15310 12930 15550
rect 13170 15310 13260 15550
rect 13500 15310 13590 15550
rect 13830 15310 13920 15550
rect 14160 15310 14250 15550
rect 14490 15310 14580 15550
rect 14820 15310 14910 15550
rect 15150 15310 15240 15550
rect 15480 15310 15570 15550
rect 15810 15310 15900 15550
rect 16140 15310 16230 15550
rect 16470 15310 16560 15550
rect 16800 15310 16890 15550
rect 17130 15310 17220 15550
rect 17460 15310 17550 15550
rect 17790 15310 17880 15550
rect 18120 15310 18210 15550
rect 18450 15310 18540 15550
rect 18780 15310 18870 15550
rect 19110 15310 19200 15550
rect 19440 15310 19530 15550
rect 19770 15310 19860 15550
rect 20100 15310 20410 15550
rect 8170 15220 20410 15310
rect 8170 14980 8310 15220
rect 8550 14980 8640 15220
rect 8880 14980 8970 15220
rect 9210 14980 9300 15220
rect 9540 14980 9630 15220
rect 9870 14980 9960 15220
rect 10200 14980 10290 15220
rect 10530 14980 10620 15220
rect 10860 14980 10950 15220
rect 11190 14980 11280 15220
rect 11520 14980 11610 15220
rect 11850 14980 11940 15220
rect 12180 14980 12270 15220
rect 12510 14980 12600 15220
rect 12840 14980 12930 15220
rect 13170 14980 13260 15220
rect 13500 14980 13590 15220
rect 13830 14980 13920 15220
rect 14160 14980 14250 15220
rect 14490 14980 14580 15220
rect 14820 14980 14910 15220
rect 15150 14980 15240 15220
rect 15480 14980 15570 15220
rect 15810 14980 15900 15220
rect 16140 14980 16230 15220
rect 16470 14980 16560 15220
rect 16800 14980 16890 15220
rect 17130 14980 17220 15220
rect 17460 14980 17550 15220
rect 17790 14980 17880 15220
rect 18120 14980 18210 15220
rect 18450 14980 18540 15220
rect 18780 14980 18870 15220
rect 19110 14980 19200 15220
rect 19440 14980 19530 15220
rect 19770 14980 19860 15220
rect 20100 14980 20410 15220
rect 8170 14890 20410 14980
rect 8170 14650 8310 14890
rect 8550 14650 8640 14890
rect 8880 14650 8970 14890
rect 9210 14650 9300 14890
rect 9540 14650 9630 14890
rect 9870 14650 9960 14890
rect 10200 14650 10290 14890
rect 10530 14650 10620 14890
rect 10860 14650 10950 14890
rect 11190 14650 11280 14890
rect 11520 14650 11610 14890
rect 11850 14650 11940 14890
rect 12180 14650 12270 14890
rect 12510 14650 12600 14890
rect 12840 14650 12930 14890
rect 13170 14650 13260 14890
rect 13500 14650 13590 14890
rect 13830 14650 13920 14890
rect 14160 14650 14250 14890
rect 14490 14650 14580 14890
rect 14820 14650 14910 14890
rect 15150 14650 15240 14890
rect 15480 14650 15570 14890
rect 15810 14650 15900 14890
rect 16140 14650 16230 14890
rect 16470 14650 16560 14890
rect 16800 14650 16890 14890
rect 17130 14650 17220 14890
rect 17460 14650 17550 14890
rect 17790 14650 17880 14890
rect 18120 14650 18210 14890
rect 18450 14650 18540 14890
rect 18780 14650 18870 14890
rect 19110 14650 19200 14890
rect 19440 14650 19530 14890
rect 19770 14650 19860 14890
rect 20100 14650 20410 14890
rect 8170 14560 20410 14650
rect 8170 14320 8310 14560
rect 8550 14320 8640 14560
rect 8880 14320 8970 14560
rect 9210 14320 9300 14560
rect 9540 14320 9630 14560
rect 9870 14320 9960 14560
rect 10200 14320 10290 14560
rect 10530 14320 10620 14560
rect 10860 14320 10950 14560
rect 11190 14320 11280 14560
rect 11520 14320 11610 14560
rect 11850 14320 11940 14560
rect 12180 14320 12270 14560
rect 12510 14320 12600 14560
rect 12840 14320 12930 14560
rect 13170 14320 13260 14560
rect 13500 14320 13590 14560
rect 13830 14320 13920 14560
rect 14160 14320 14250 14560
rect 14490 14320 14580 14560
rect 14820 14320 14910 14560
rect 15150 14320 15240 14560
rect 15480 14320 15570 14560
rect 15810 14320 15900 14560
rect 16140 14320 16230 14560
rect 16470 14320 16560 14560
rect 16800 14320 16890 14560
rect 17130 14320 17220 14560
rect 17460 14320 17550 14560
rect 17790 14320 17880 14560
rect 18120 14320 18210 14560
rect 18450 14320 18540 14560
rect 18780 14320 18870 14560
rect 19110 14320 19200 14560
rect 19440 14320 19530 14560
rect 19770 14320 19860 14560
rect 20100 14320 20410 14560
rect 8170 14230 20410 14320
rect 8170 13990 8310 14230
rect 8550 13990 8640 14230
rect 8880 13990 8970 14230
rect 9210 13990 9300 14230
rect 9540 13990 9630 14230
rect 9870 13990 9960 14230
rect 10200 13990 10290 14230
rect 10530 13990 10620 14230
rect 10860 13990 10950 14230
rect 11190 13990 11280 14230
rect 11520 13990 11610 14230
rect 11850 13990 11940 14230
rect 12180 13990 12270 14230
rect 12510 13990 12600 14230
rect 12840 13990 12930 14230
rect 13170 13990 13260 14230
rect 13500 13990 13590 14230
rect 13830 13990 13920 14230
rect 14160 13990 14250 14230
rect 14490 13990 14580 14230
rect 14820 13990 14910 14230
rect 15150 13990 15240 14230
rect 15480 13990 15570 14230
rect 15810 13990 15900 14230
rect 16140 13990 16230 14230
rect 16470 13990 16560 14230
rect 16800 13990 16890 14230
rect 17130 13990 17220 14230
rect 17460 13990 17550 14230
rect 17790 13990 17880 14230
rect 18120 13990 18210 14230
rect 18450 13990 18540 14230
rect 18780 13990 18870 14230
rect 19110 13990 19200 14230
rect 19440 13990 19530 14230
rect 19770 13990 19860 14230
rect 20100 13990 20410 14230
rect 8170 13900 20410 13990
rect 8170 13660 8310 13900
rect 8550 13660 8640 13900
rect 8880 13660 8970 13900
rect 9210 13660 9300 13900
rect 9540 13660 9630 13900
rect 9870 13660 9960 13900
rect 10200 13660 10290 13900
rect 10530 13660 10620 13900
rect 10860 13660 10950 13900
rect 11190 13660 11280 13900
rect 11520 13660 11610 13900
rect 11850 13660 11940 13900
rect 12180 13660 12270 13900
rect 12510 13660 12600 13900
rect 12840 13660 12930 13900
rect 13170 13660 13260 13900
rect 13500 13660 13590 13900
rect 13830 13660 13920 13900
rect 14160 13660 14250 13900
rect 14490 13660 14580 13900
rect 14820 13660 14910 13900
rect 15150 13660 15240 13900
rect 15480 13660 15570 13900
rect 15810 13660 15900 13900
rect 16140 13660 16230 13900
rect 16470 13660 16560 13900
rect 16800 13660 16890 13900
rect 17130 13660 17220 13900
rect 17460 13660 17550 13900
rect 17790 13660 17880 13900
rect 18120 13660 18210 13900
rect 18450 13660 18540 13900
rect 18780 13660 18870 13900
rect 19110 13660 19200 13900
rect 19440 13660 19530 13900
rect 19770 13660 19860 13900
rect 20100 13660 20410 13900
rect 8170 13570 20410 13660
rect 8170 13330 8310 13570
rect 8550 13330 8640 13570
rect 8880 13330 8970 13570
rect 9210 13330 9300 13570
rect 9540 13330 9630 13570
rect 9870 13330 9960 13570
rect 10200 13330 10290 13570
rect 10530 13330 10620 13570
rect 10860 13330 10950 13570
rect 11190 13330 11280 13570
rect 11520 13330 11610 13570
rect 11850 13330 11940 13570
rect 12180 13330 12270 13570
rect 12510 13330 12600 13570
rect 12840 13330 12930 13570
rect 13170 13330 13260 13570
rect 13500 13330 13590 13570
rect 13830 13330 13920 13570
rect 14160 13330 14250 13570
rect 14490 13330 14580 13570
rect 14820 13330 14910 13570
rect 15150 13330 15240 13570
rect 15480 13330 15570 13570
rect 15810 13330 15900 13570
rect 16140 13330 16230 13570
rect 16470 13330 16560 13570
rect 16800 13330 16890 13570
rect 17130 13330 17220 13570
rect 17460 13330 17550 13570
rect 17790 13330 17880 13570
rect 18120 13330 18210 13570
rect 18450 13330 18540 13570
rect 18780 13330 18870 13570
rect 19110 13330 19200 13570
rect 19440 13330 19530 13570
rect 19770 13330 19860 13570
rect 20100 13330 20410 13570
rect 8170 13240 20410 13330
rect 8170 13000 8310 13240
rect 8550 13000 8640 13240
rect 8880 13000 8970 13240
rect 9210 13000 9300 13240
rect 9540 13000 9630 13240
rect 9870 13000 9960 13240
rect 10200 13000 10290 13240
rect 10530 13000 10620 13240
rect 10860 13000 10950 13240
rect 11190 13000 11280 13240
rect 11520 13000 11610 13240
rect 11850 13000 11940 13240
rect 12180 13000 12270 13240
rect 12510 13000 12600 13240
rect 12840 13000 12930 13240
rect 13170 13000 13260 13240
rect 13500 13000 13590 13240
rect 13830 13000 13920 13240
rect 14160 13000 14250 13240
rect 14490 13000 14580 13240
rect 14820 13000 14910 13240
rect 15150 13000 15240 13240
rect 15480 13000 15570 13240
rect 15810 13000 15900 13240
rect 16140 13000 16230 13240
rect 16470 13000 16560 13240
rect 16800 13000 16890 13240
rect 17130 13000 17220 13240
rect 17460 13000 17550 13240
rect 17790 13000 17880 13240
rect 18120 13000 18210 13240
rect 18450 13000 18540 13240
rect 18780 13000 18870 13240
rect 19110 13000 19200 13240
rect 19440 13000 19530 13240
rect 19770 13000 19860 13240
rect 20100 13000 20410 13240
rect 8170 12910 20410 13000
rect 8170 12670 8310 12910
rect 8550 12670 8640 12910
rect 8880 12670 8970 12910
rect 9210 12670 9300 12910
rect 9540 12670 9630 12910
rect 9870 12670 9960 12910
rect 10200 12670 10290 12910
rect 10530 12670 10620 12910
rect 10860 12670 10950 12910
rect 11190 12670 11280 12910
rect 11520 12670 11610 12910
rect 11850 12670 11940 12910
rect 12180 12670 12270 12910
rect 12510 12670 12600 12910
rect 12840 12670 12930 12910
rect 13170 12670 13260 12910
rect 13500 12670 13590 12910
rect 13830 12670 13920 12910
rect 14160 12670 14250 12910
rect 14490 12670 14580 12910
rect 14820 12670 14910 12910
rect 15150 12670 15240 12910
rect 15480 12670 15570 12910
rect 15810 12670 15900 12910
rect 16140 12670 16230 12910
rect 16470 12670 16560 12910
rect 16800 12670 16890 12910
rect 17130 12670 17220 12910
rect 17460 12670 17550 12910
rect 17790 12670 17880 12910
rect 18120 12670 18210 12910
rect 18450 12670 18540 12910
rect 18780 12670 18870 12910
rect 19110 12670 19200 12910
rect 19440 12670 19530 12910
rect 19770 12670 19860 12910
rect 20100 12670 20410 12910
rect 8170 12580 20410 12670
rect 8170 12340 8310 12580
rect 8550 12340 8640 12580
rect 8880 12340 8970 12580
rect 9210 12340 9300 12580
rect 9540 12340 9630 12580
rect 9870 12340 9960 12580
rect 10200 12340 10290 12580
rect 10530 12340 10620 12580
rect 10860 12340 10950 12580
rect 11190 12340 11280 12580
rect 11520 12340 11610 12580
rect 11850 12340 11940 12580
rect 12180 12340 12270 12580
rect 12510 12340 12600 12580
rect 12840 12340 12930 12580
rect 13170 12340 13260 12580
rect 13500 12340 13590 12580
rect 13830 12340 13920 12580
rect 14160 12340 14250 12580
rect 14490 12340 14580 12580
rect 14820 12340 14910 12580
rect 15150 12340 15240 12580
rect 15480 12340 15570 12580
rect 15810 12340 15900 12580
rect 16140 12340 16230 12580
rect 16470 12340 16560 12580
rect 16800 12340 16890 12580
rect 17130 12340 17220 12580
rect 17460 12340 17550 12580
rect 17790 12340 17880 12580
rect 18120 12340 18210 12580
rect 18450 12340 18540 12580
rect 18780 12340 18870 12580
rect 19110 12340 19200 12580
rect 19440 12340 19530 12580
rect 19770 12340 19860 12580
rect 20100 12340 20410 12580
rect 8170 12250 20410 12340
rect 8170 12010 8310 12250
rect 8550 12010 8640 12250
rect 8880 12010 8970 12250
rect 9210 12010 9300 12250
rect 9540 12010 9630 12250
rect 9870 12010 9960 12250
rect 10200 12010 10290 12250
rect 10530 12010 10620 12250
rect 10860 12010 10950 12250
rect 11190 12010 11280 12250
rect 11520 12010 11610 12250
rect 11850 12010 11940 12250
rect 12180 12010 12270 12250
rect 12510 12010 12600 12250
rect 12840 12010 12930 12250
rect 13170 12010 13260 12250
rect 13500 12010 13590 12250
rect 13830 12010 13920 12250
rect 14160 12010 14250 12250
rect 14490 12010 14580 12250
rect 14820 12010 14910 12250
rect 15150 12010 15240 12250
rect 15480 12010 15570 12250
rect 15810 12010 15900 12250
rect 16140 12010 16230 12250
rect 16470 12010 16560 12250
rect 16800 12010 16890 12250
rect 17130 12010 17220 12250
rect 17460 12010 17550 12250
rect 17790 12010 17880 12250
rect 18120 12010 18210 12250
rect 18450 12010 18540 12250
rect 18780 12010 18870 12250
rect 19110 12010 19200 12250
rect 19440 12010 19530 12250
rect 19770 12010 19860 12250
rect 20100 12010 20410 12250
rect 8170 11920 20410 12010
rect 8170 11680 8310 11920
rect 8550 11680 8640 11920
rect 8880 11680 8970 11920
rect 9210 11680 9300 11920
rect 9540 11680 9630 11920
rect 9870 11680 9960 11920
rect 10200 11680 10290 11920
rect 10530 11680 10620 11920
rect 10860 11680 10950 11920
rect 11190 11680 11280 11920
rect 11520 11680 11610 11920
rect 11850 11680 11940 11920
rect 12180 11680 12270 11920
rect 12510 11680 12600 11920
rect 12840 11680 12930 11920
rect 13170 11680 13260 11920
rect 13500 11680 13590 11920
rect 13830 11680 13920 11920
rect 14160 11680 14250 11920
rect 14490 11680 14580 11920
rect 14820 11680 14910 11920
rect 15150 11680 15240 11920
rect 15480 11680 15570 11920
rect 15810 11680 15900 11920
rect 16140 11680 16230 11920
rect 16470 11680 16560 11920
rect 16800 11680 16890 11920
rect 17130 11680 17220 11920
rect 17460 11680 17550 11920
rect 17790 11680 17880 11920
rect 18120 11680 18210 11920
rect 18450 11680 18540 11920
rect 18780 11680 18870 11920
rect 19110 11680 19200 11920
rect 19440 11680 19530 11920
rect 19770 11680 19860 11920
rect 20100 11680 20410 11920
rect 8170 11590 20410 11680
rect 8170 11350 8310 11590
rect 8550 11350 8640 11590
rect 8880 11350 8970 11590
rect 9210 11350 9300 11590
rect 9540 11350 9630 11590
rect 9870 11350 9960 11590
rect 10200 11350 10290 11590
rect 10530 11350 10620 11590
rect 10860 11350 10950 11590
rect 11190 11350 11280 11590
rect 11520 11350 11610 11590
rect 11850 11350 11940 11590
rect 12180 11350 12270 11590
rect 12510 11350 12600 11590
rect 12840 11350 12930 11590
rect 13170 11350 13260 11590
rect 13500 11350 13590 11590
rect 13830 11350 13920 11590
rect 14160 11350 14250 11590
rect 14490 11350 14580 11590
rect 14820 11350 14910 11590
rect 15150 11350 15240 11590
rect 15480 11350 15570 11590
rect 15810 11350 15900 11590
rect 16140 11350 16230 11590
rect 16470 11350 16560 11590
rect 16800 11350 16890 11590
rect 17130 11350 17220 11590
rect 17460 11350 17550 11590
rect 17790 11350 17880 11590
rect 18120 11350 18210 11590
rect 18450 11350 18540 11590
rect 18780 11350 18870 11590
rect 19110 11350 19200 11590
rect 19440 11350 19530 11590
rect 19770 11350 19860 11590
rect 20100 11350 20410 11590
rect 8170 11260 20410 11350
rect 8170 11020 8310 11260
rect 8550 11020 8640 11260
rect 8880 11020 8970 11260
rect 9210 11020 9300 11260
rect 9540 11020 9630 11260
rect 9870 11020 9960 11260
rect 10200 11020 10290 11260
rect 10530 11020 10620 11260
rect 10860 11020 10950 11260
rect 11190 11020 11280 11260
rect 11520 11020 11610 11260
rect 11850 11020 11940 11260
rect 12180 11020 12270 11260
rect 12510 11020 12600 11260
rect 12840 11020 12930 11260
rect 13170 11020 13260 11260
rect 13500 11020 13590 11260
rect 13830 11020 13920 11260
rect 14160 11020 14250 11260
rect 14490 11020 14580 11260
rect 14820 11020 14910 11260
rect 15150 11020 15240 11260
rect 15480 11020 15570 11260
rect 15810 11020 15900 11260
rect 16140 11020 16230 11260
rect 16470 11020 16560 11260
rect 16800 11020 16890 11260
rect 17130 11020 17220 11260
rect 17460 11020 17550 11260
rect 17790 11020 17880 11260
rect 18120 11020 18210 11260
rect 18450 11020 18540 11260
rect 18780 11020 18870 11260
rect 19110 11020 19200 11260
rect 19440 11020 19530 11260
rect 19770 11020 19860 11260
rect 20100 11020 20410 11260
rect 8170 10930 20410 11020
rect 8170 10690 8310 10930
rect 8550 10690 8640 10930
rect 8880 10690 8970 10930
rect 9210 10690 9300 10930
rect 9540 10690 9630 10930
rect 9870 10690 9960 10930
rect 10200 10690 10290 10930
rect 10530 10690 10620 10930
rect 10860 10690 10950 10930
rect 11190 10690 11280 10930
rect 11520 10690 11610 10930
rect 11850 10690 11940 10930
rect 12180 10690 12270 10930
rect 12510 10690 12600 10930
rect 12840 10690 12930 10930
rect 13170 10690 13260 10930
rect 13500 10690 13590 10930
rect 13830 10690 13920 10930
rect 14160 10690 14250 10930
rect 14490 10690 14580 10930
rect 14820 10690 14910 10930
rect 15150 10690 15240 10930
rect 15480 10690 15570 10930
rect 15810 10690 15900 10930
rect 16140 10690 16230 10930
rect 16470 10690 16560 10930
rect 16800 10690 16890 10930
rect 17130 10690 17220 10930
rect 17460 10690 17550 10930
rect 17790 10690 17880 10930
rect 18120 10690 18210 10930
rect 18450 10690 18540 10930
rect 18780 10690 18870 10930
rect 19110 10690 19200 10930
rect 19440 10690 19530 10930
rect 19770 10690 19860 10930
rect 20100 10690 20410 10930
rect 8170 10600 20410 10690
rect 8170 10360 8310 10600
rect 8550 10360 8640 10600
rect 8880 10360 8970 10600
rect 9210 10360 9300 10600
rect 9540 10360 9630 10600
rect 9870 10360 9960 10600
rect 10200 10360 10290 10600
rect 10530 10360 10620 10600
rect 10860 10360 10950 10600
rect 11190 10360 11280 10600
rect 11520 10360 11610 10600
rect 11850 10360 11940 10600
rect 12180 10360 12270 10600
rect 12510 10360 12600 10600
rect 12840 10360 12930 10600
rect 13170 10360 13260 10600
rect 13500 10360 13590 10600
rect 13830 10360 13920 10600
rect 14160 10360 14250 10600
rect 14490 10360 14580 10600
rect 14820 10360 14910 10600
rect 15150 10360 15240 10600
rect 15480 10360 15570 10600
rect 15810 10360 15900 10600
rect 16140 10360 16230 10600
rect 16470 10360 16560 10600
rect 16800 10360 16890 10600
rect 17130 10360 17220 10600
rect 17460 10360 17550 10600
rect 17790 10360 17880 10600
rect 18120 10360 18210 10600
rect 18450 10360 18540 10600
rect 18780 10360 18870 10600
rect 19110 10360 19200 10600
rect 19440 10360 19530 10600
rect 19770 10360 19860 10600
rect 20100 10360 20410 10600
rect 8170 10270 20410 10360
rect 8170 10030 8310 10270
rect 8550 10030 8640 10270
rect 8880 10030 8970 10270
rect 9210 10030 9300 10270
rect 9540 10030 9630 10270
rect 9870 10030 9960 10270
rect 10200 10030 10290 10270
rect 10530 10030 10620 10270
rect 10860 10030 10950 10270
rect 11190 10030 11280 10270
rect 11520 10030 11610 10270
rect 11850 10030 11940 10270
rect 12180 10030 12270 10270
rect 12510 10030 12600 10270
rect 12840 10030 12930 10270
rect 13170 10030 13260 10270
rect 13500 10030 13590 10270
rect 13830 10030 13920 10270
rect 14160 10030 14250 10270
rect 14490 10030 14580 10270
rect 14820 10030 14910 10270
rect 15150 10030 15240 10270
rect 15480 10030 15570 10270
rect 15810 10030 15900 10270
rect 16140 10030 16230 10270
rect 16470 10030 16560 10270
rect 16800 10030 16890 10270
rect 17130 10030 17220 10270
rect 17460 10030 17550 10270
rect 17790 10030 17880 10270
rect 18120 10030 18210 10270
rect 18450 10030 18540 10270
rect 18780 10030 18870 10270
rect 19110 10030 19200 10270
rect 19440 10030 19530 10270
rect 19770 10030 19860 10270
rect 20100 10030 20410 10270
rect 8170 9940 20410 10030
rect 8170 9700 8310 9940
rect 8550 9700 8640 9940
rect 8880 9700 8970 9940
rect 9210 9700 9300 9940
rect 9540 9700 9630 9940
rect 9870 9700 9960 9940
rect 10200 9700 10290 9940
rect 10530 9700 10620 9940
rect 10860 9700 10950 9940
rect 11190 9700 11280 9940
rect 11520 9700 11610 9940
rect 11850 9700 11940 9940
rect 12180 9700 12270 9940
rect 12510 9700 12600 9940
rect 12840 9700 12930 9940
rect 13170 9700 13260 9940
rect 13500 9700 13590 9940
rect 13830 9700 13920 9940
rect 14160 9700 14250 9940
rect 14490 9700 14580 9940
rect 14820 9700 14910 9940
rect 15150 9700 15240 9940
rect 15480 9700 15570 9940
rect 15810 9700 15900 9940
rect 16140 9700 16230 9940
rect 16470 9700 16560 9940
rect 16800 9700 16890 9940
rect 17130 9700 17220 9940
rect 17460 9700 17550 9940
rect 17790 9700 17880 9940
rect 18120 9700 18210 9940
rect 18450 9700 18540 9940
rect 18780 9700 18870 9940
rect 19110 9700 19200 9940
rect 19440 9700 19530 9940
rect 19770 9700 19860 9940
rect 20100 9700 20410 9940
rect 8170 9610 20410 9700
rect 8170 9370 8310 9610
rect 8550 9370 8640 9610
rect 8880 9370 8970 9610
rect 9210 9370 9300 9610
rect 9540 9370 9630 9610
rect 9870 9370 9960 9610
rect 10200 9370 10290 9610
rect 10530 9370 10620 9610
rect 10860 9370 10950 9610
rect 11190 9370 11280 9610
rect 11520 9370 11610 9610
rect 11850 9370 11940 9610
rect 12180 9370 12270 9610
rect 12510 9370 12600 9610
rect 12840 9370 12930 9610
rect 13170 9370 13260 9610
rect 13500 9370 13590 9610
rect 13830 9370 13920 9610
rect 14160 9370 14250 9610
rect 14490 9370 14580 9610
rect 14820 9370 14910 9610
rect 15150 9370 15240 9610
rect 15480 9370 15570 9610
rect 15810 9370 15900 9610
rect 16140 9370 16230 9610
rect 16470 9370 16560 9610
rect 16800 9370 16890 9610
rect 17130 9370 17220 9610
rect 17460 9370 17550 9610
rect 17790 9370 17880 9610
rect 18120 9370 18210 9610
rect 18450 9370 18540 9610
rect 18780 9370 18870 9610
rect 19110 9370 19200 9610
rect 19440 9370 19530 9610
rect 19770 9370 19860 9610
rect 20100 9370 20410 9610
rect 8170 9280 20410 9370
rect 8170 9040 8310 9280
rect 8550 9040 8640 9280
rect 8880 9040 8970 9280
rect 9210 9040 9300 9280
rect 9540 9040 9630 9280
rect 9870 9040 9960 9280
rect 10200 9040 10290 9280
rect 10530 9040 10620 9280
rect 10860 9040 10950 9280
rect 11190 9040 11280 9280
rect 11520 9040 11610 9280
rect 11850 9040 11940 9280
rect 12180 9040 12270 9280
rect 12510 9040 12600 9280
rect 12840 9040 12930 9280
rect 13170 9040 13260 9280
rect 13500 9040 13590 9280
rect 13830 9040 13920 9280
rect 14160 9040 14250 9280
rect 14490 9040 14580 9280
rect 14820 9040 14910 9280
rect 15150 9040 15240 9280
rect 15480 9040 15570 9280
rect 15810 9040 15900 9280
rect 16140 9040 16230 9280
rect 16470 9040 16560 9280
rect 16800 9040 16890 9280
rect 17130 9040 17220 9280
rect 17460 9040 17550 9280
rect 17790 9040 17880 9280
rect 18120 9040 18210 9280
rect 18450 9040 18540 9280
rect 18780 9040 18870 9280
rect 19110 9040 19200 9280
rect 19440 9040 19530 9280
rect 19770 9040 19860 9280
rect 20100 9040 20410 9280
rect 8170 8720 20410 9040
rect 31130 7830 37830 7880
rect 31130 7590 31180 7830
rect 31420 7590 31510 7830
rect 31750 7590 31840 7830
rect 32080 7590 32170 7830
rect 32410 7590 32500 7830
rect 32740 7590 32830 7830
rect 33070 7590 33160 7830
rect 33400 7590 33490 7830
rect 33730 7590 33820 7830
rect 34060 7590 34150 7830
rect 34390 7590 34480 7830
rect 34720 7590 34810 7830
rect 35050 7590 35140 7830
rect 35380 7590 35470 7830
rect 35710 7590 35800 7830
rect 36040 7590 36130 7830
rect 36370 7590 36460 7830
rect 36700 7590 36790 7830
rect 37030 7590 37120 7830
rect 37360 7590 37450 7830
rect 37690 7590 37830 7830
rect 31130 7500 37830 7590
rect 31130 7260 31180 7500
rect 31420 7260 31510 7500
rect 31750 7260 31840 7500
rect 32080 7260 32170 7500
rect 32410 7260 32500 7500
rect 32740 7260 32830 7500
rect 33070 7260 33160 7500
rect 33400 7260 33490 7500
rect 33730 7260 33820 7500
rect 34060 7260 34150 7500
rect 34390 7260 34480 7500
rect 34720 7260 34810 7500
rect 35050 7260 35140 7500
rect 35380 7260 35470 7500
rect 35710 7260 35800 7500
rect 36040 7260 36130 7500
rect 36370 7260 36460 7500
rect 36700 7260 36790 7500
rect 37030 7260 37120 7500
rect 37360 7260 37450 7500
rect 37690 7260 37830 7500
rect 31130 7170 37830 7260
rect 31130 6930 31180 7170
rect 31420 6930 31510 7170
rect 31750 6930 31840 7170
rect 32080 6930 32170 7170
rect 32410 6930 32500 7170
rect 32740 6930 32830 7170
rect 33070 6930 33160 7170
rect 33400 6930 33490 7170
rect 33730 6930 33820 7170
rect 34060 6930 34150 7170
rect 34390 6930 34480 7170
rect 34720 6930 34810 7170
rect 35050 6930 35140 7170
rect 35380 6930 35470 7170
rect 35710 6930 35800 7170
rect 36040 6930 36130 7170
rect 36370 6930 36460 7170
rect 36700 6930 36790 7170
rect 37030 6930 37120 7170
rect 37360 6930 37450 7170
rect 37690 6930 37830 7170
rect 31130 6840 37830 6930
rect 31130 6600 31180 6840
rect 31420 6600 31510 6840
rect 31750 6600 31840 6840
rect 32080 6600 32170 6840
rect 32410 6600 32500 6840
rect 32740 6600 32830 6840
rect 33070 6600 33160 6840
rect 33400 6600 33490 6840
rect 33730 6600 33820 6840
rect 34060 6600 34150 6840
rect 34390 6600 34480 6840
rect 34720 6600 34810 6840
rect 35050 6600 35140 6840
rect 35380 6600 35470 6840
rect 35710 6600 35800 6840
rect 36040 6600 36130 6840
rect 36370 6600 36460 6840
rect 36700 6600 36790 6840
rect 37030 6600 37120 6840
rect 37360 6600 37450 6840
rect 37690 6600 37830 6840
rect 31130 6510 37830 6600
rect 31130 6270 31180 6510
rect 31420 6270 31510 6510
rect 31750 6270 31840 6510
rect 32080 6270 32170 6510
rect 32410 6270 32500 6510
rect 32740 6270 32830 6510
rect 33070 6270 33160 6510
rect 33400 6270 33490 6510
rect 33730 6270 33820 6510
rect 34060 6270 34150 6510
rect 34390 6270 34480 6510
rect 34720 6270 34810 6510
rect 35050 6270 35140 6510
rect 35380 6270 35470 6510
rect 35710 6270 35800 6510
rect 36040 6270 36130 6510
rect 36370 6270 36460 6510
rect 36700 6270 36790 6510
rect 37030 6270 37120 6510
rect 37360 6270 37450 6510
rect 37690 6270 37830 6510
rect 31130 6180 37830 6270
rect 31130 5940 31180 6180
rect 31420 5940 31510 6180
rect 31750 5940 31840 6180
rect 32080 5940 32170 6180
rect 32410 5940 32500 6180
rect 32740 5940 32830 6180
rect 33070 5940 33160 6180
rect 33400 5940 33490 6180
rect 33730 5940 33820 6180
rect 34060 5940 34150 6180
rect 34390 5940 34480 6180
rect 34720 5940 34810 6180
rect 35050 5940 35140 6180
rect 35380 5940 35470 6180
rect 35710 5940 35800 6180
rect 36040 5940 36130 6180
rect 36370 5940 36460 6180
rect 36700 5940 36790 6180
rect 37030 5940 37120 6180
rect 37360 5940 37450 6180
rect 37690 5940 37830 6180
rect 31130 5850 37830 5940
rect 31130 5610 31180 5850
rect 31420 5610 31510 5850
rect 31750 5610 31840 5850
rect 32080 5610 32170 5850
rect 32410 5610 32500 5850
rect 32740 5610 32830 5850
rect 33070 5610 33160 5850
rect 33400 5610 33490 5850
rect 33730 5610 33820 5850
rect 34060 5610 34150 5850
rect 34390 5610 34480 5850
rect 34720 5610 34810 5850
rect 35050 5610 35140 5850
rect 35380 5610 35470 5850
rect 35710 5610 35800 5850
rect 36040 5610 36130 5850
rect 36370 5610 36460 5850
rect 36700 5610 36790 5850
rect 37030 5610 37120 5850
rect 37360 5610 37450 5850
rect 37690 5610 37830 5850
rect 31130 5520 37830 5610
rect 31130 5280 31180 5520
rect 31420 5280 31510 5520
rect 31750 5280 31840 5520
rect 32080 5280 32170 5520
rect 32410 5280 32500 5520
rect 32740 5280 32830 5520
rect 33070 5280 33160 5520
rect 33400 5280 33490 5520
rect 33730 5280 33820 5520
rect 34060 5280 34150 5520
rect 34390 5280 34480 5520
rect 34720 5280 34810 5520
rect 35050 5280 35140 5520
rect 35380 5280 35470 5520
rect 35710 5280 35800 5520
rect 36040 5280 36130 5520
rect 36370 5280 36460 5520
rect 36700 5280 36790 5520
rect 37030 5280 37120 5520
rect 37360 5280 37450 5520
rect 37690 5280 37830 5520
rect 31130 5190 37830 5280
rect 31130 4950 31180 5190
rect 31420 4950 31510 5190
rect 31750 4950 31840 5190
rect 32080 4950 32170 5190
rect 32410 4950 32500 5190
rect 32740 4950 32830 5190
rect 33070 4950 33160 5190
rect 33400 4950 33490 5190
rect 33730 4950 33820 5190
rect 34060 4950 34150 5190
rect 34390 4950 34480 5190
rect 34720 4950 34810 5190
rect 35050 4950 35140 5190
rect 35380 4950 35470 5190
rect 35710 4950 35800 5190
rect 36040 4950 36130 5190
rect 36370 4950 36460 5190
rect 36700 4950 36790 5190
rect 37030 4950 37120 5190
rect 37360 4950 37450 5190
rect 37690 4950 37830 5190
rect 31130 4860 37830 4950
rect 31130 4620 31180 4860
rect 31420 4620 31510 4860
rect 31750 4620 31840 4860
rect 32080 4620 32170 4860
rect 32410 4620 32500 4860
rect 32740 4620 32830 4860
rect 33070 4620 33160 4860
rect 33400 4620 33490 4860
rect 33730 4620 33820 4860
rect 34060 4620 34150 4860
rect 34390 4620 34480 4860
rect 34720 4620 34810 4860
rect 35050 4620 35140 4860
rect 35380 4620 35470 4860
rect 35710 4620 35800 4860
rect 36040 4620 36130 4860
rect 36370 4620 36460 4860
rect 36700 4620 36790 4860
rect 37030 4620 37120 4860
rect 37360 4620 37450 4860
rect 37690 4620 37830 4860
rect 31130 4530 37830 4620
rect 31130 4290 31180 4530
rect 31420 4290 31510 4530
rect 31750 4290 31840 4530
rect 32080 4290 32170 4530
rect 32410 4290 32500 4530
rect 32740 4290 32830 4530
rect 33070 4290 33160 4530
rect 33400 4290 33490 4530
rect 33730 4290 33820 4530
rect 34060 4290 34150 4530
rect 34390 4290 34480 4530
rect 34720 4290 34810 4530
rect 35050 4290 35140 4530
rect 35380 4290 35470 4530
rect 35710 4290 35800 4530
rect 36040 4290 36130 4530
rect 36370 4290 36460 4530
rect 36700 4290 36790 4530
rect 37030 4290 37120 4530
rect 37360 4290 37450 4530
rect 37690 4290 37830 4530
rect 31130 4200 37830 4290
rect 31130 3960 31180 4200
rect 31420 3960 31510 4200
rect 31750 3960 31840 4200
rect 32080 3960 32170 4200
rect 32410 3960 32500 4200
rect 32740 3960 32830 4200
rect 33070 3960 33160 4200
rect 33400 3960 33490 4200
rect 33730 3960 33820 4200
rect 34060 3960 34150 4200
rect 34390 3960 34480 4200
rect 34720 3960 34810 4200
rect 35050 3960 35140 4200
rect 35380 3960 35470 4200
rect 35710 3960 35800 4200
rect 36040 3960 36130 4200
rect 36370 3960 36460 4200
rect 36700 3960 36790 4200
rect 37030 3960 37120 4200
rect 37360 3960 37450 4200
rect 37690 3960 37830 4200
rect 31130 3870 37830 3960
rect 31130 3630 31180 3870
rect 31420 3630 31510 3870
rect 31750 3630 31840 3870
rect 32080 3630 32170 3870
rect 32410 3630 32500 3870
rect 32740 3630 32830 3870
rect 33070 3630 33160 3870
rect 33400 3630 33490 3870
rect 33730 3630 33820 3870
rect 34060 3630 34150 3870
rect 34390 3630 34480 3870
rect 34720 3630 34810 3870
rect 35050 3630 35140 3870
rect 35380 3630 35470 3870
rect 35710 3630 35800 3870
rect 36040 3630 36130 3870
rect 36370 3630 36460 3870
rect 36700 3630 36790 3870
rect 37030 3630 37120 3870
rect 37360 3630 37450 3870
rect 37690 3630 37830 3870
rect 31130 3540 37830 3630
rect 31130 3300 31180 3540
rect 31420 3300 31510 3540
rect 31750 3300 31840 3540
rect 32080 3300 32170 3540
rect 32410 3300 32500 3540
rect 32740 3300 32830 3540
rect 33070 3300 33160 3540
rect 33400 3300 33490 3540
rect 33730 3300 33820 3540
rect 34060 3300 34150 3540
rect 34390 3300 34480 3540
rect 34720 3300 34810 3540
rect 35050 3300 35140 3540
rect 35380 3300 35470 3540
rect 35710 3300 35800 3540
rect 36040 3300 36130 3540
rect 36370 3300 36460 3540
rect 36700 3300 36790 3540
rect 37030 3300 37120 3540
rect 37360 3300 37450 3540
rect 37690 3300 37830 3540
rect 31130 3210 37830 3300
rect 31130 2970 31180 3210
rect 31420 2970 31510 3210
rect 31750 2970 31840 3210
rect 32080 2970 32170 3210
rect 32410 2970 32500 3210
rect 32740 2970 32830 3210
rect 33070 2970 33160 3210
rect 33400 2970 33490 3210
rect 33730 2970 33820 3210
rect 34060 2970 34150 3210
rect 34390 2970 34480 3210
rect 34720 2970 34810 3210
rect 35050 2970 35140 3210
rect 35380 2970 35470 3210
rect 35710 2970 35800 3210
rect 36040 2970 36130 3210
rect 36370 2970 36460 3210
rect 36700 2970 36790 3210
rect 37030 2970 37120 3210
rect 37360 2970 37450 3210
rect 37690 2970 37830 3210
rect 31130 2880 37830 2970
rect 31130 2640 31180 2880
rect 31420 2640 31510 2880
rect 31750 2640 31840 2880
rect 32080 2640 32170 2880
rect 32410 2640 32500 2880
rect 32740 2640 32830 2880
rect 33070 2640 33160 2880
rect 33400 2640 33490 2880
rect 33730 2640 33820 2880
rect 34060 2640 34150 2880
rect 34390 2640 34480 2880
rect 34720 2640 34810 2880
rect 35050 2640 35140 2880
rect 35380 2640 35470 2880
rect 35710 2640 35800 2880
rect 36040 2640 36130 2880
rect 36370 2640 36460 2880
rect 36700 2640 36790 2880
rect 37030 2640 37120 2880
rect 37360 2640 37450 2880
rect 37690 2640 37830 2880
rect 31130 2550 37830 2640
rect 31130 2310 31180 2550
rect 31420 2310 31510 2550
rect 31750 2310 31840 2550
rect 32080 2310 32170 2550
rect 32410 2310 32500 2550
rect 32740 2310 32830 2550
rect 33070 2310 33160 2550
rect 33400 2310 33490 2550
rect 33730 2310 33820 2550
rect 34060 2310 34150 2550
rect 34390 2310 34480 2550
rect 34720 2310 34810 2550
rect 35050 2310 35140 2550
rect 35380 2310 35470 2550
rect 35710 2310 35800 2550
rect 36040 2310 36130 2550
rect 36370 2310 36460 2550
rect 36700 2310 36790 2550
rect 37030 2310 37120 2550
rect 37360 2310 37450 2550
rect 37690 2310 37830 2550
rect 31130 2220 37830 2310
rect 31130 1980 31180 2220
rect 31420 1980 31510 2220
rect 31750 1980 31840 2220
rect 32080 1980 32170 2220
rect 32410 1980 32500 2220
rect 32740 1980 32830 2220
rect 33070 1980 33160 2220
rect 33400 1980 33490 2220
rect 33730 1980 33820 2220
rect 34060 1980 34150 2220
rect 34390 1980 34480 2220
rect 34720 1980 34810 2220
rect 35050 1980 35140 2220
rect 35380 1980 35470 2220
rect 35710 1980 35800 2220
rect 36040 1980 36130 2220
rect 36370 1980 36460 2220
rect 36700 1980 36790 2220
rect 37030 1980 37120 2220
rect 37360 1980 37450 2220
rect 37690 1980 37830 2220
rect 31130 1890 37830 1980
rect 31130 1650 31180 1890
rect 31420 1650 31510 1890
rect 31750 1650 31840 1890
rect 32080 1650 32170 1890
rect 32410 1650 32500 1890
rect 32740 1650 32830 1890
rect 33070 1650 33160 1890
rect 33400 1650 33490 1890
rect 33730 1650 33820 1890
rect 34060 1650 34150 1890
rect 34390 1650 34480 1890
rect 34720 1650 34810 1890
rect 35050 1650 35140 1890
rect 35380 1650 35470 1890
rect 35710 1650 35800 1890
rect 36040 1650 36130 1890
rect 36370 1650 36460 1890
rect 36700 1650 36790 1890
rect 37030 1650 37120 1890
rect 37360 1650 37450 1890
rect 37690 1650 37830 1890
rect 31130 1560 37830 1650
rect 31130 1320 31180 1560
rect 31420 1320 31510 1560
rect 31750 1320 31840 1560
rect 32080 1320 32170 1560
rect 32410 1320 32500 1560
rect 32740 1320 32830 1560
rect 33070 1320 33160 1560
rect 33400 1320 33490 1560
rect 33730 1320 33820 1560
rect 34060 1320 34150 1560
rect 34390 1320 34480 1560
rect 34720 1320 34810 1560
rect 35050 1320 35140 1560
rect 35380 1320 35470 1560
rect 35710 1320 35800 1560
rect 36040 1320 36130 1560
rect 36370 1320 36460 1560
rect 36700 1320 36790 1560
rect 37030 1320 37120 1560
rect 37360 1320 37450 1560
rect 37690 1320 37830 1560
rect 31130 1180 37830 1320
rect 31130 230 37830 280
rect 31130 -10 31180 230
rect 31420 -10 31510 230
rect 31750 -10 31840 230
rect 32080 -10 32170 230
rect 32410 -10 32500 230
rect 32740 -10 32830 230
rect 33070 -10 33160 230
rect 33400 -10 33490 230
rect 33730 -10 33820 230
rect 34060 -10 34150 230
rect 34390 -10 34480 230
rect 34720 -10 34810 230
rect 35050 -10 35140 230
rect 35380 -10 35470 230
rect 35710 -10 35800 230
rect 36040 -10 36130 230
rect 36370 -10 36460 230
rect 36700 -10 36790 230
rect 37030 -10 37120 230
rect 37360 -10 37450 230
rect 37690 -10 37830 230
rect 31130 -100 37830 -10
rect 31130 -340 31180 -100
rect 31420 -340 31510 -100
rect 31750 -340 31840 -100
rect 32080 -340 32170 -100
rect 32410 -340 32500 -100
rect 32740 -340 32830 -100
rect 33070 -340 33160 -100
rect 33400 -340 33490 -100
rect 33730 -340 33820 -100
rect 34060 -340 34150 -100
rect 34390 -340 34480 -100
rect 34720 -340 34810 -100
rect 35050 -340 35140 -100
rect 35380 -340 35470 -100
rect 35710 -340 35800 -100
rect 36040 -340 36130 -100
rect 36370 -340 36460 -100
rect 36700 -340 36790 -100
rect 37030 -340 37120 -100
rect 37360 -340 37450 -100
rect 37690 -340 37830 -100
rect 31130 -430 37830 -340
rect 31130 -670 31180 -430
rect 31420 -670 31510 -430
rect 31750 -670 31840 -430
rect 32080 -670 32170 -430
rect 32410 -670 32500 -430
rect 32740 -670 32830 -430
rect 33070 -670 33160 -430
rect 33400 -670 33490 -430
rect 33730 -670 33820 -430
rect 34060 -670 34150 -430
rect 34390 -670 34480 -430
rect 34720 -670 34810 -430
rect 35050 -670 35140 -430
rect 35380 -670 35470 -430
rect 35710 -670 35800 -430
rect 36040 -670 36130 -430
rect 36370 -670 36460 -430
rect 36700 -670 36790 -430
rect 37030 -670 37120 -430
rect 37360 -670 37450 -430
rect 37690 -670 37830 -430
rect 31130 -760 37830 -670
rect 31130 -1000 31180 -760
rect 31420 -1000 31510 -760
rect 31750 -1000 31840 -760
rect 32080 -1000 32170 -760
rect 32410 -1000 32500 -760
rect 32740 -1000 32830 -760
rect 33070 -1000 33160 -760
rect 33400 -1000 33490 -760
rect 33730 -1000 33820 -760
rect 34060 -1000 34150 -760
rect 34390 -1000 34480 -760
rect 34720 -1000 34810 -760
rect 35050 -1000 35140 -760
rect 35380 -1000 35470 -760
rect 35710 -1000 35800 -760
rect 36040 -1000 36130 -760
rect 36370 -1000 36460 -760
rect 36700 -1000 36790 -760
rect 37030 -1000 37120 -760
rect 37360 -1000 37450 -760
rect 37690 -1000 37830 -760
rect 31130 -1090 37830 -1000
rect 31130 -1330 31180 -1090
rect 31420 -1330 31510 -1090
rect 31750 -1330 31840 -1090
rect 32080 -1330 32170 -1090
rect 32410 -1330 32500 -1090
rect 32740 -1330 32830 -1090
rect 33070 -1330 33160 -1090
rect 33400 -1330 33490 -1090
rect 33730 -1330 33820 -1090
rect 34060 -1330 34150 -1090
rect 34390 -1330 34480 -1090
rect 34720 -1330 34810 -1090
rect 35050 -1330 35140 -1090
rect 35380 -1330 35470 -1090
rect 35710 -1330 35800 -1090
rect 36040 -1330 36130 -1090
rect 36370 -1330 36460 -1090
rect 36700 -1330 36790 -1090
rect 37030 -1330 37120 -1090
rect 37360 -1330 37450 -1090
rect 37690 -1330 37830 -1090
rect 31130 -1420 37830 -1330
rect 31130 -1660 31180 -1420
rect 31420 -1660 31510 -1420
rect 31750 -1660 31840 -1420
rect 32080 -1660 32170 -1420
rect 32410 -1660 32500 -1420
rect 32740 -1660 32830 -1420
rect 33070 -1660 33160 -1420
rect 33400 -1660 33490 -1420
rect 33730 -1660 33820 -1420
rect 34060 -1660 34150 -1420
rect 34390 -1660 34480 -1420
rect 34720 -1660 34810 -1420
rect 35050 -1660 35140 -1420
rect 35380 -1660 35470 -1420
rect 35710 -1660 35800 -1420
rect 36040 -1660 36130 -1420
rect 36370 -1660 36460 -1420
rect 36700 -1660 36790 -1420
rect 37030 -1660 37120 -1420
rect 37360 -1660 37450 -1420
rect 37690 -1660 37830 -1420
rect 31130 -1750 37830 -1660
rect 31130 -1990 31180 -1750
rect 31420 -1990 31510 -1750
rect 31750 -1990 31840 -1750
rect 32080 -1990 32170 -1750
rect 32410 -1990 32500 -1750
rect 32740 -1990 32830 -1750
rect 33070 -1990 33160 -1750
rect 33400 -1990 33490 -1750
rect 33730 -1990 33820 -1750
rect 34060 -1990 34150 -1750
rect 34390 -1990 34480 -1750
rect 34720 -1990 34810 -1750
rect 35050 -1990 35140 -1750
rect 35380 -1990 35470 -1750
rect 35710 -1990 35800 -1750
rect 36040 -1990 36130 -1750
rect 36370 -1990 36460 -1750
rect 36700 -1990 36790 -1750
rect 37030 -1990 37120 -1750
rect 37360 -1990 37450 -1750
rect 37690 -1990 37830 -1750
rect 31130 -2080 37830 -1990
rect 31130 -2320 31180 -2080
rect 31420 -2320 31510 -2080
rect 31750 -2320 31840 -2080
rect 32080 -2320 32170 -2080
rect 32410 -2320 32500 -2080
rect 32740 -2320 32830 -2080
rect 33070 -2320 33160 -2080
rect 33400 -2320 33490 -2080
rect 33730 -2320 33820 -2080
rect 34060 -2320 34150 -2080
rect 34390 -2320 34480 -2080
rect 34720 -2320 34810 -2080
rect 35050 -2320 35140 -2080
rect 35380 -2320 35470 -2080
rect 35710 -2320 35800 -2080
rect 36040 -2320 36130 -2080
rect 36370 -2320 36460 -2080
rect 36700 -2320 36790 -2080
rect 37030 -2320 37120 -2080
rect 37360 -2320 37450 -2080
rect 37690 -2320 37830 -2080
rect 31130 -2410 37830 -2320
rect 31130 -2650 31180 -2410
rect 31420 -2650 31510 -2410
rect 31750 -2650 31840 -2410
rect 32080 -2650 32170 -2410
rect 32410 -2650 32500 -2410
rect 32740 -2650 32830 -2410
rect 33070 -2650 33160 -2410
rect 33400 -2650 33490 -2410
rect 33730 -2650 33820 -2410
rect 34060 -2650 34150 -2410
rect 34390 -2650 34480 -2410
rect 34720 -2650 34810 -2410
rect 35050 -2650 35140 -2410
rect 35380 -2650 35470 -2410
rect 35710 -2650 35800 -2410
rect 36040 -2650 36130 -2410
rect 36370 -2650 36460 -2410
rect 36700 -2650 36790 -2410
rect 37030 -2650 37120 -2410
rect 37360 -2650 37450 -2410
rect 37690 -2650 37830 -2410
rect 31130 -2740 37830 -2650
rect 31130 -2980 31180 -2740
rect 31420 -2980 31510 -2740
rect 31750 -2980 31840 -2740
rect 32080 -2980 32170 -2740
rect 32410 -2980 32500 -2740
rect 32740 -2980 32830 -2740
rect 33070 -2980 33160 -2740
rect 33400 -2980 33490 -2740
rect 33730 -2980 33820 -2740
rect 34060 -2980 34150 -2740
rect 34390 -2980 34480 -2740
rect 34720 -2980 34810 -2740
rect 35050 -2980 35140 -2740
rect 35380 -2980 35470 -2740
rect 35710 -2980 35800 -2740
rect 36040 -2980 36130 -2740
rect 36370 -2980 36460 -2740
rect 36700 -2980 36790 -2740
rect 37030 -2980 37120 -2740
rect 37360 -2980 37450 -2740
rect 37690 -2980 37830 -2740
rect 31130 -3070 37830 -2980
rect 31130 -3310 31180 -3070
rect 31420 -3310 31510 -3070
rect 31750 -3310 31840 -3070
rect 32080 -3310 32170 -3070
rect 32410 -3310 32500 -3070
rect 32740 -3310 32830 -3070
rect 33070 -3310 33160 -3070
rect 33400 -3310 33490 -3070
rect 33730 -3310 33820 -3070
rect 34060 -3310 34150 -3070
rect 34390 -3310 34480 -3070
rect 34720 -3310 34810 -3070
rect 35050 -3310 35140 -3070
rect 35380 -3310 35470 -3070
rect 35710 -3310 35800 -3070
rect 36040 -3310 36130 -3070
rect 36370 -3310 36460 -3070
rect 36700 -3310 36790 -3070
rect 37030 -3310 37120 -3070
rect 37360 -3310 37450 -3070
rect 37690 -3310 37830 -3070
rect 31130 -3400 37830 -3310
rect 31130 -3640 31180 -3400
rect 31420 -3640 31510 -3400
rect 31750 -3640 31840 -3400
rect 32080 -3640 32170 -3400
rect 32410 -3640 32500 -3400
rect 32740 -3640 32830 -3400
rect 33070 -3640 33160 -3400
rect 33400 -3640 33490 -3400
rect 33730 -3640 33820 -3400
rect 34060 -3640 34150 -3400
rect 34390 -3640 34480 -3400
rect 34720 -3640 34810 -3400
rect 35050 -3640 35140 -3400
rect 35380 -3640 35470 -3400
rect 35710 -3640 35800 -3400
rect 36040 -3640 36130 -3400
rect 36370 -3640 36460 -3400
rect 36700 -3640 36790 -3400
rect 37030 -3640 37120 -3400
rect 37360 -3640 37450 -3400
rect 37690 -3640 37830 -3400
rect 31130 -3730 37830 -3640
rect 31130 -3970 31180 -3730
rect 31420 -3970 31510 -3730
rect 31750 -3970 31840 -3730
rect 32080 -3970 32170 -3730
rect 32410 -3970 32500 -3730
rect 32740 -3970 32830 -3730
rect 33070 -3970 33160 -3730
rect 33400 -3970 33490 -3730
rect 33730 -3970 33820 -3730
rect 34060 -3970 34150 -3730
rect 34390 -3970 34480 -3730
rect 34720 -3970 34810 -3730
rect 35050 -3970 35140 -3730
rect 35380 -3970 35470 -3730
rect 35710 -3970 35800 -3730
rect 36040 -3970 36130 -3730
rect 36370 -3970 36460 -3730
rect 36700 -3970 36790 -3730
rect 37030 -3970 37120 -3730
rect 37360 -3970 37450 -3730
rect 37690 -3970 37830 -3730
rect 31130 -4060 37830 -3970
rect 31130 -4300 31180 -4060
rect 31420 -4300 31510 -4060
rect 31750 -4300 31840 -4060
rect 32080 -4300 32170 -4060
rect 32410 -4300 32500 -4060
rect 32740 -4300 32830 -4060
rect 33070 -4300 33160 -4060
rect 33400 -4300 33490 -4060
rect 33730 -4300 33820 -4060
rect 34060 -4300 34150 -4060
rect 34390 -4300 34480 -4060
rect 34720 -4300 34810 -4060
rect 35050 -4300 35140 -4060
rect 35380 -4300 35470 -4060
rect 35710 -4300 35800 -4060
rect 36040 -4300 36130 -4060
rect 36370 -4300 36460 -4060
rect 36700 -4300 36790 -4060
rect 37030 -4300 37120 -4060
rect 37360 -4300 37450 -4060
rect 37690 -4300 37830 -4060
rect 31130 -4390 37830 -4300
rect 31130 -4630 31180 -4390
rect 31420 -4630 31510 -4390
rect 31750 -4630 31840 -4390
rect 32080 -4630 32170 -4390
rect 32410 -4630 32500 -4390
rect 32740 -4630 32830 -4390
rect 33070 -4630 33160 -4390
rect 33400 -4630 33490 -4390
rect 33730 -4630 33820 -4390
rect 34060 -4630 34150 -4390
rect 34390 -4630 34480 -4390
rect 34720 -4630 34810 -4390
rect 35050 -4630 35140 -4390
rect 35380 -4630 35470 -4390
rect 35710 -4630 35800 -4390
rect 36040 -4630 36130 -4390
rect 36370 -4630 36460 -4390
rect 36700 -4630 36790 -4390
rect 37030 -4630 37120 -4390
rect 37360 -4630 37450 -4390
rect 37690 -4630 37830 -4390
rect -1320 -4840 230 -4660
rect -1320 -5080 -1180 -4840
rect -940 -5080 -850 -4840
rect -610 -5080 -520 -4840
rect -280 -5080 -190 -4840
rect 50 -5080 230 -4840
rect -1320 -5170 230 -5080
rect -1320 -5410 -1180 -5170
rect -940 -5410 -850 -5170
rect -610 -5410 -520 -5170
rect -280 -5410 -190 -5170
rect 50 -5410 230 -5170
rect -1320 -5500 230 -5410
rect -1320 -5740 -1180 -5500
rect -940 -5740 -850 -5500
rect -610 -5740 -520 -5500
rect -280 -5740 -190 -5500
rect 50 -5740 230 -5500
rect -1320 -5830 230 -5740
rect -1320 -6070 -1180 -5830
rect -940 -6070 -850 -5830
rect -610 -6070 -520 -5830
rect -280 -6070 -190 -5830
rect 50 -6070 230 -5830
rect -1320 -6210 230 -6070
rect 14550 -4840 16100 -4660
rect 14550 -5080 14730 -4840
rect 14970 -5080 15060 -4840
rect 15300 -5080 15390 -4840
rect 15630 -5080 15720 -4840
rect 15960 -5080 16100 -4840
rect 14550 -5170 16100 -5080
rect 14550 -5410 14730 -5170
rect 14970 -5410 15060 -5170
rect 15300 -5410 15390 -5170
rect 15630 -5410 15720 -5170
rect 15960 -5410 16100 -5170
rect 14550 -5500 16100 -5410
rect 14550 -5740 14730 -5500
rect 14970 -5740 15060 -5500
rect 15300 -5740 15390 -5500
rect 15630 -5740 15720 -5500
rect 15960 -5740 16100 -5500
rect 14550 -5830 16100 -5740
rect 14550 -6070 14730 -5830
rect 14970 -6070 15060 -5830
rect 15300 -6070 15390 -5830
rect 15630 -6070 15720 -5830
rect 15960 -6070 16100 -5830
rect 14550 -6210 16100 -6070
rect 31130 -4720 37830 -4630
rect 31130 -4960 31180 -4720
rect 31420 -4960 31510 -4720
rect 31750 -4960 31840 -4720
rect 32080 -4960 32170 -4720
rect 32410 -4960 32500 -4720
rect 32740 -4960 32830 -4720
rect 33070 -4960 33160 -4720
rect 33400 -4960 33490 -4720
rect 33730 -4960 33820 -4720
rect 34060 -4960 34150 -4720
rect 34390 -4960 34480 -4720
rect 34720 -4960 34810 -4720
rect 35050 -4960 35140 -4720
rect 35380 -4960 35470 -4720
rect 35710 -4960 35800 -4720
rect 36040 -4960 36130 -4720
rect 36370 -4960 36460 -4720
rect 36700 -4960 36790 -4720
rect 37030 -4960 37120 -4720
rect 37360 -4960 37450 -4720
rect 37690 -4960 37830 -4720
rect 31130 -5050 37830 -4960
rect 31130 -5290 31180 -5050
rect 31420 -5290 31510 -5050
rect 31750 -5290 31840 -5050
rect 32080 -5290 32170 -5050
rect 32410 -5290 32500 -5050
rect 32740 -5290 32830 -5050
rect 33070 -5290 33160 -5050
rect 33400 -5290 33490 -5050
rect 33730 -5290 33820 -5050
rect 34060 -5290 34150 -5050
rect 34390 -5290 34480 -5050
rect 34720 -5290 34810 -5050
rect 35050 -5290 35140 -5050
rect 35380 -5290 35470 -5050
rect 35710 -5290 35800 -5050
rect 36040 -5290 36130 -5050
rect 36370 -5290 36460 -5050
rect 36700 -5290 36790 -5050
rect 37030 -5290 37120 -5050
rect 37360 -5290 37450 -5050
rect 37690 -5290 37830 -5050
rect 31130 -5380 37830 -5290
rect 31130 -5620 31180 -5380
rect 31420 -5620 31510 -5380
rect 31750 -5620 31840 -5380
rect 32080 -5620 32170 -5380
rect 32410 -5620 32500 -5380
rect 32740 -5620 32830 -5380
rect 33070 -5620 33160 -5380
rect 33400 -5620 33490 -5380
rect 33730 -5620 33820 -5380
rect 34060 -5620 34150 -5380
rect 34390 -5620 34480 -5380
rect 34720 -5620 34810 -5380
rect 35050 -5620 35140 -5380
rect 35380 -5620 35470 -5380
rect 35710 -5620 35800 -5380
rect 36040 -5620 36130 -5380
rect 36370 -5620 36460 -5380
rect 36700 -5620 36790 -5380
rect 37030 -5620 37120 -5380
rect 37360 -5620 37450 -5380
rect 37690 -5620 37830 -5380
rect 31130 -5710 37830 -5620
rect 31130 -5950 31180 -5710
rect 31420 -5950 31510 -5710
rect 31750 -5950 31840 -5710
rect 32080 -5950 32170 -5710
rect 32410 -5950 32500 -5710
rect 32740 -5950 32830 -5710
rect 33070 -5950 33160 -5710
rect 33400 -5950 33490 -5710
rect 33730 -5950 33820 -5710
rect 34060 -5950 34150 -5710
rect 34390 -5950 34480 -5710
rect 34720 -5950 34810 -5710
rect 35050 -5950 35140 -5710
rect 35380 -5950 35470 -5710
rect 35710 -5950 35800 -5710
rect 36040 -5950 36130 -5710
rect 36370 -5950 36460 -5710
rect 36700 -5950 36790 -5710
rect 37030 -5950 37120 -5710
rect 37360 -5950 37450 -5710
rect 37690 -5950 37830 -5710
rect 31130 -6040 37830 -5950
rect 31130 -6280 31180 -6040
rect 31420 -6280 31510 -6040
rect 31750 -6280 31840 -6040
rect 32080 -6280 32170 -6040
rect 32410 -6280 32500 -6040
rect 32740 -6280 32830 -6040
rect 33070 -6280 33160 -6040
rect 33400 -6280 33490 -6040
rect 33730 -6280 33820 -6040
rect 34060 -6280 34150 -6040
rect 34390 -6280 34480 -6040
rect 34720 -6280 34810 -6040
rect 35050 -6280 35140 -6040
rect 35380 -6280 35470 -6040
rect 35710 -6280 35800 -6040
rect 36040 -6280 36130 -6040
rect 36370 -6280 36460 -6040
rect 36700 -6280 36790 -6040
rect 37030 -6280 37120 -6040
rect 37360 -6280 37450 -6040
rect 37690 -6280 37830 -6040
rect 31130 -6420 37830 -6280
<< mimcap2contact >>
rect -5200 20590 -4960 20830
rect -4870 20590 -4630 20830
rect -4540 20590 -4300 20830
rect -4210 20590 -3970 20830
rect -3880 20590 -3640 20830
rect -3550 20590 -3310 20830
rect -3220 20590 -2980 20830
rect -2890 20590 -2650 20830
rect -2560 20590 -2320 20830
rect -2230 20590 -1990 20830
rect -1900 20590 -1660 20830
rect -1570 20590 -1330 20830
rect -1240 20590 -1000 20830
rect -910 20590 -670 20830
rect -580 20590 -340 20830
rect -250 20590 -10 20830
rect 80 20590 320 20830
rect 410 20590 650 20830
rect 740 20590 980 20830
rect 1070 20590 1310 20830
rect 1400 20590 1640 20830
rect 1730 20590 1970 20830
rect 2060 20590 2300 20830
rect 2390 20590 2630 20830
rect 2720 20590 2960 20830
rect 3050 20590 3290 20830
rect 3380 20590 3620 20830
rect 3710 20590 3950 20830
rect 4040 20590 4280 20830
rect 4370 20590 4610 20830
rect 4700 20590 4940 20830
rect 5030 20590 5270 20830
rect 5360 20590 5600 20830
rect 5690 20590 5930 20830
rect 6020 20590 6260 20830
rect 6350 20590 6590 20830
rect -5200 20260 -4960 20500
rect -4870 20260 -4630 20500
rect -4540 20260 -4300 20500
rect -4210 20260 -3970 20500
rect -3880 20260 -3640 20500
rect -3550 20260 -3310 20500
rect -3220 20260 -2980 20500
rect -2890 20260 -2650 20500
rect -2560 20260 -2320 20500
rect -2230 20260 -1990 20500
rect -1900 20260 -1660 20500
rect -1570 20260 -1330 20500
rect -1240 20260 -1000 20500
rect -910 20260 -670 20500
rect -580 20260 -340 20500
rect -250 20260 -10 20500
rect 80 20260 320 20500
rect 410 20260 650 20500
rect 740 20260 980 20500
rect 1070 20260 1310 20500
rect 1400 20260 1640 20500
rect 1730 20260 1970 20500
rect 2060 20260 2300 20500
rect 2390 20260 2630 20500
rect 2720 20260 2960 20500
rect 3050 20260 3290 20500
rect 3380 20260 3620 20500
rect 3710 20260 3950 20500
rect 4040 20260 4280 20500
rect 4370 20260 4610 20500
rect 4700 20260 4940 20500
rect 5030 20260 5270 20500
rect 5360 20260 5600 20500
rect 5690 20260 5930 20500
rect 6020 20260 6260 20500
rect 6350 20260 6590 20500
rect -5200 19930 -4960 20170
rect -4870 19930 -4630 20170
rect -4540 19930 -4300 20170
rect -4210 19930 -3970 20170
rect -3880 19930 -3640 20170
rect -3550 19930 -3310 20170
rect -3220 19930 -2980 20170
rect -2890 19930 -2650 20170
rect -2560 19930 -2320 20170
rect -2230 19930 -1990 20170
rect -1900 19930 -1660 20170
rect -1570 19930 -1330 20170
rect -1240 19930 -1000 20170
rect -910 19930 -670 20170
rect -580 19930 -340 20170
rect -250 19930 -10 20170
rect 80 19930 320 20170
rect 410 19930 650 20170
rect 740 19930 980 20170
rect 1070 19930 1310 20170
rect 1400 19930 1640 20170
rect 1730 19930 1970 20170
rect 2060 19930 2300 20170
rect 2390 19930 2630 20170
rect 2720 19930 2960 20170
rect 3050 19930 3290 20170
rect 3380 19930 3620 20170
rect 3710 19930 3950 20170
rect 4040 19930 4280 20170
rect 4370 19930 4610 20170
rect 4700 19930 4940 20170
rect 5030 19930 5270 20170
rect 5360 19930 5600 20170
rect 5690 19930 5930 20170
rect 6020 19930 6260 20170
rect 6350 19930 6590 20170
rect -5200 19600 -4960 19840
rect -4870 19600 -4630 19840
rect -4540 19600 -4300 19840
rect -4210 19600 -3970 19840
rect -3880 19600 -3640 19840
rect -3550 19600 -3310 19840
rect -3220 19600 -2980 19840
rect -2890 19600 -2650 19840
rect -2560 19600 -2320 19840
rect -2230 19600 -1990 19840
rect -1900 19600 -1660 19840
rect -1570 19600 -1330 19840
rect -1240 19600 -1000 19840
rect -910 19600 -670 19840
rect -580 19600 -340 19840
rect -250 19600 -10 19840
rect 80 19600 320 19840
rect 410 19600 650 19840
rect 740 19600 980 19840
rect 1070 19600 1310 19840
rect 1400 19600 1640 19840
rect 1730 19600 1970 19840
rect 2060 19600 2300 19840
rect 2390 19600 2630 19840
rect 2720 19600 2960 19840
rect 3050 19600 3290 19840
rect 3380 19600 3620 19840
rect 3710 19600 3950 19840
rect 4040 19600 4280 19840
rect 4370 19600 4610 19840
rect 4700 19600 4940 19840
rect 5030 19600 5270 19840
rect 5360 19600 5600 19840
rect 5690 19600 5930 19840
rect 6020 19600 6260 19840
rect 6350 19600 6590 19840
rect -5200 19270 -4960 19510
rect -4870 19270 -4630 19510
rect -4540 19270 -4300 19510
rect -4210 19270 -3970 19510
rect -3880 19270 -3640 19510
rect -3550 19270 -3310 19510
rect -3220 19270 -2980 19510
rect -2890 19270 -2650 19510
rect -2560 19270 -2320 19510
rect -2230 19270 -1990 19510
rect -1900 19270 -1660 19510
rect -1570 19270 -1330 19510
rect -1240 19270 -1000 19510
rect -910 19270 -670 19510
rect -580 19270 -340 19510
rect -250 19270 -10 19510
rect 80 19270 320 19510
rect 410 19270 650 19510
rect 740 19270 980 19510
rect 1070 19270 1310 19510
rect 1400 19270 1640 19510
rect 1730 19270 1970 19510
rect 2060 19270 2300 19510
rect 2390 19270 2630 19510
rect 2720 19270 2960 19510
rect 3050 19270 3290 19510
rect 3380 19270 3620 19510
rect 3710 19270 3950 19510
rect 4040 19270 4280 19510
rect 4370 19270 4610 19510
rect 4700 19270 4940 19510
rect 5030 19270 5270 19510
rect 5360 19270 5600 19510
rect 5690 19270 5930 19510
rect 6020 19270 6260 19510
rect 6350 19270 6590 19510
rect -5200 18940 -4960 19180
rect -4870 18940 -4630 19180
rect -4540 18940 -4300 19180
rect -4210 18940 -3970 19180
rect -3880 18940 -3640 19180
rect -3550 18940 -3310 19180
rect -3220 18940 -2980 19180
rect -2890 18940 -2650 19180
rect -2560 18940 -2320 19180
rect -2230 18940 -1990 19180
rect -1900 18940 -1660 19180
rect -1570 18940 -1330 19180
rect -1240 18940 -1000 19180
rect -910 18940 -670 19180
rect -580 18940 -340 19180
rect -250 18940 -10 19180
rect 80 18940 320 19180
rect 410 18940 650 19180
rect 740 18940 980 19180
rect 1070 18940 1310 19180
rect 1400 18940 1640 19180
rect 1730 18940 1970 19180
rect 2060 18940 2300 19180
rect 2390 18940 2630 19180
rect 2720 18940 2960 19180
rect 3050 18940 3290 19180
rect 3380 18940 3620 19180
rect 3710 18940 3950 19180
rect 4040 18940 4280 19180
rect 4370 18940 4610 19180
rect 4700 18940 4940 19180
rect 5030 18940 5270 19180
rect 5360 18940 5600 19180
rect 5690 18940 5930 19180
rect 6020 18940 6260 19180
rect 6350 18940 6590 19180
rect -5200 18610 -4960 18850
rect -4870 18610 -4630 18850
rect -4540 18610 -4300 18850
rect -4210 18610 -3970 18850
rect -3880 18610 -3640 18850
rect -3550 18610 -3310 18850
rect -3220 18610 -2980 18850
rect -2890 18610 -2650 18850
rect -2560 18610 -2320 18850
rect -2230 18610 -1990 18850
rect -1900 18610 -1660 18850
rect -1570 18610 -1330 18850
rect -1240 18610 -1000 18850
rect -910 18610 -670 18850
rect -580 18610 -340 18850
rect -250 18610 -10 18850
rect 80 18610 320 18850
rect 410 18610 650 18850
rect 740 18610 980 18850
rect 1070 18610 1310 18850
rect 1400 18610 1640 18850
rect 1730 18610 1970 18850
rect 2060 18610 2300 18850
rect 2390 18610 2630 18850
rect 2720 18610 2960 18850
rect 3050 18610 3290 18850
rect 3380 18610 3620 18850
rect 3710 18610 3950 18850
rect 4040 18610 4280 18850
rect 4370 18610 4610 18850
rect 4700 18610 4940 18850
rect 5030 18610 5270 18850
rect 5360 18610 5600 18850
rect 5690 18610 5930 18850
rect 6020 18610 6260 18850
rect 6350 18610 6590 18850
rect -5200 18280 -4960 18520
rect -4870 18280 -4630 18520
rect -4540 18280 -4300 18520
rect -4210 18280 -3970 18520
rect -3880 18280 -3640 18520
rect -3550 18280 -3310 18520
rect -3220 18280 -2980 18520
rect -2890 18280 -2650 18520
rect -2560 18280 -2320 18520
rect -2230 18280 -1990 18520
rect -1900 18280 -1660 18520
rect -1570 18280 -1330 18520
rect -1240 18280 -1000 18520
rect -910 18280 -670 18520
rect -580 18280 -340 18520
rect -250 18280 -10 18520
rect 80 18280 320 18520
rect 410 18280 650 18520
rect 740 18280 980 18520
rect 1070 18280 1310 18520
rect 1400 18280 1640 18520
rect 1730 18280 1970 18520
rect 2060 18280 2300 18520
rect 2390 18280 2630 18520
rect 2720 18280 2960 18520
rect 3050 18280 3290 18520
rect 3380 18280 3620 18520
rect 3710 18280 3950 18520
rect 4040 18280 4280 18520
rect 4370 18280 4610 18520
rect 4700 18280 4940 18520
rect 5030 18280 5270 18520
rect 5360 18280 5600 18520
rect 5690 18280 5930 18520
rect 6020 18280 6260 18520
rect 6350 18280 6590 18520
rect -5200 17950 -4960 18190
rect -4870 17950 -4630 18190
rect -4540 17950 -4300 18190
rect -4210 17950 -3970 18190
rect -3880 17950 -3640 18190
rect -3550 17950 -3310 18190
rect -3220 17950 -2980 18190
rect -2890 17950 -2650 18190
rect -2560 17950 -2320 18190
rect -2230 17950 -1990 18190
rect -1900 17950 -1660 18190
rect -1570 17950 -1330 18190
rect -1240 17950 -1000 18190
rect -910 17950 -670 18190
rect -580 17950 -340 18190
rect -250 17950 -10 18190
rect 80 17950 320 18190
rect 410 17950 650 18190
rect 740 17950 980 18190
rect 1070 17950 1310 18190
rect 1400 17950 1640 18190
rect 1730 17950 1970 18190
rect 2060 17950 2300 18190
rect 2390 17950 2630 18190
rect 2720 17950 2960 18190
rect 3050 17950 3290 18190
rect 3380 17950 3620 18190
rect 3710 17950 3950 18190
rect 4040 17950 4280 18190
rect 4370 17950 4610 18190
rect 4700 17950 4940 18190
rect 5030 17950 5270 18190
rect 5360 17950 5600 18190
rect 5690 17950 5930 18190
rect 6020 17950 6260 18190
rect 6350 17950 6590 18190
rect -5200 17620 -4960 17860
rect -4870 17620 -4630 17860
rect -4540 17620 -4300 17860
rect -4210 17620 -3970 17860
rect -3880 17620 -3640 17860
rect -3550 17620 -3310 17860
rect -3220 17620 -2980 17860
rect -2890 17620 -2650 17860
rect -2560 17620 -2320 17860
rect -2230 17620 -1990 17860
rect -1900 17620 -1660 17860
rect -1570 17620 -1330 17860
rect -1240 17620 -1000 17860
rect -910 17620 -670 17860
rect -580 17620 -340 17860
rect -250 17620 -10 17860
rect 80 17620 320 17860
rect 410 17620 650 17860
rect 740 17620 980 17860
rect 1070 17620 1310 17860
rect 1400 17620 1640 17860
rect 1730 17620 1970 17860
rect 2060 17620 2300 17860
rect 2390 17620 2630 17860
rect 2720 17620 2960 17860
rect 3050 17620 3290 17860
rect 3380 17620 3620 17860
rect 3710 17620 3950 17860
rect 4040 17620 4280 17860
rect 4370 17620 4610 17860
rect 4700 17620 4940 17860
rect 5030 17620 5270 17860
rect 5360 17620 5600 17860
rect 5690 17620 5930 17860
rect 6020 17620 6260 17860
rect 6350 17620 6590 17860
rect -5200 17290 -4960 17530
rect -4870 17290 -4630 17530
rect -4540 17290 -4300 17530
rect -4210 17290 -3970 17530
rect -3880 17290 -3640 17530
rect -3550 17290 -3310 17530
rect -3220 17290 -2980 17530
rect -2890 17290 -2650 17530
rect -2560 17290 -2320 17530
rect -2230 17290 -1990 17530
rect -1900 17290 -1660 17530
rect -1570 17290 -1330 17530
rect -1240 17290 -1000 17530
rect -910 17290 -670 17530
rect -580 17290 -340 17530
rect -250 17290 -10 17530
rect 80 17290 320 17530
rect 410 17290 650 17530
rect 740 17290 980 17530
rect 1070 17290 1310 17530
rect 1400 17290 1640 17530
rect 1730 17290 1970 17530
rect 2060 17290 2300 17530
rect 2390 17290 2630 17530
rect 2720 17290 2960 17530
rect 3050 17290 3290 17530
rect 3380 17290 3620 17530
rect 3710 17290 3950 17530
rect 4040 17290 4280 17530
rect 4370 17290 4610 17530
rect 4700 17290 4940 17530
rect 5030 17290 5270 17530
rect 5360 17290 5600 17530
rect 5690 17290 5930 17530
rect 6020 17290 6260 17530
rect 6350 17290 6590 17530
rect -5200 16960 -4960 17200
rect -4870 16960 -4630 17200
rect -4540 16960 -4300 17200
rect -4210 16960 -3970 17200
rect -3880 16960 -3640 17200
rect -3550 16960 -3310 17200
rect -3220 16960 -2980 17200
rect -2890 16960 -2650 17200
rect -2560 16960 -2320 17200
rect -2230 16960 -1990 17200
rect -1900 16960 -1660 17200
rect -1570 16960 -1330 17200
rect -1240 16960 -1000 17200
rect -910 16960 -670 17200
rect -580 16960 -340 17200
rect -250 16960 -10 17200
rect 80 16960 320 17200
rect 410 16960 650 17200
rect 740 16960 980 17200
rect 1070 16960 1310 17200
rect 1400 16960 1640 17200
rect 1730 16960 1970 17200
rect 2060 16960 2300 17200
rect 2390 16960 2630 17200
rect 2720 16960 2960 17200
rect 3050 16960 3290 17200
rect 3380 16960 3620 17200
rect 3710 16960 3950 17200
rect 4040 16960 4280 17200
rect 4370 16960 4610 17200
rect 4700 16960 4940 17200
rect 5030 16960 5270 17200
rect 5360 16960 5600 17200
rect 5690 16960 5930 17200
rect 6020 16960 6260 17200
rect 6350 16960 6590 17200
rect -5200 16630 -4960 16870
rect -4870 16630 -4630 16870
rect -4540 16630 -4300 16870
rect -4210 16630 -3970 16870
rect -3880 16630 -3640 16870
rect -3550 16630 -3310 16870
rect -3220 16630 -2980 16870
rect -2890 16630 -2650 16870
rect -2560 16630 -2320 16870
rect -2230 16630 -1990 16870
rect -1900 16630 -1660 16870
rect -1570 16630 -1330 16870
rect -1240 16630 -1000 16870
rect -910 16630 -670 16870
rect -580 16630 -340 16870
rect -250 16630 -10 16870
rect 80 16630 320 16870
rect 410 16630 650 16870
rect 740 16630 980 16870
rect 1070 16630 1310 16870
rect 1400 16630 1640 16870
rect 1730 16630 1970 16870
rect 2060 16630 2300 16870
rect 2390 16630 2630 16870
rect 2720 16630 2960 16870
rect 3050 16630 3290 16870
rect 3380 16630 3620 16870
rect 3710 16630 3950 16870
rect 4040 16630 4280 16870
rect 4370 16630 4610 16870
rect 4700 16630 4940 16870
rect 5030 16630 5270 16870
rect 5360 16630 5600 16870
rect 5690 16630 5930 16870
rect 6020 16630 6260 16870
rect 6350 16630 6590 16870
rect -5200 16300 -4960 16540
rect -4870 16300 -4630 16540
rect -4540 16300 -4300 16540
rect -4210 16300 -3970 16540
rect -3880 16300 -3640 16540
rect -3550 16300 -3310 16540
rect -3220 16300 -2980 16540
rect -2890 16300 -2650 16540
rect -2560 16300 -2320 16540
rect -2230 16300 -1990 16540
rect -1900 16300 -1660 16540
rect -1570 16300 -1330 16540
rect -1240 16300 -1000 16540
rect -910 16300 -670 16540
rect -580 16300 -340 16540
rect -250 16300 -10 16540
rect 80 16300 320 16540
rect 410 16300 650 16540
rect 740 16300 980 16540
rect 1070 16300 1310 16540
rect 1400 16300 1640 16540
rect 1730 16300 1970 16540
rect 2060 16300 2300 16540
rect 2390 16300 2630 16540
rect 2720 16300 2960 16540
rect 3050 16300 3290 16540
rect 3380 16300 3620 16540
rect 3710 16300 3950 16540
rect 4040 16300 4280 16540
rect 4370 16300 4610 16540
rect 4700 16300 4940 16540
rect 5030 16300 5270 16540
rect 5360 16300 5600 16540
rect 5690 16300 5930 16540
rect 6020 16300 6260 16540
rect 6350 16300 6590 16540
rect -5200 15970 -4960 16210
rect -4870 15970 -4630 16210
rect -4540 15970 -4300 16210
rect -4210 15970 -3970 16210
rect -3880 15970 -3640 16210
rect -3550 15970 -3310 16210
rect -3220 15970 -2980 16210
rect -2890 15970 -2650 16210
rect -2560 15970 -2320 16210
rect -2230 15970 -1990 16210
rect -1900 15970 -1660 16210
rect -1570 15970 -1330 16210
rect -1240 15970 -1000 16210
rect -910 15970 -670 16210
rect -580 15970 -340 16210
rect -250 15970 -10 16210
rect 80 15970 320 16210
rect 410 15970 650 16210
rect 740 15970 980 16210
rect 1070 15970 1310 16210
rect 1400 15970 1640 16210
rect 1730 15970 1970 16210
rect 2060 15970 2300 16210
rect 2390 15970 2630 16210
rect 2720 15970 2960 16210
rect 3050 15970 3290 16210
rect 3380 15970 3620 16210
rect 3710 15970 3950 16210
rect 4040 15970 4280 16210
rect 4370 15970 4610 16210
rect 4700 15970 4940 16210
rect 5030 15970 5270 16210
rect 5360 15970 5600 16210
rect 5690 15970 5930 16210
rect 6020 15970 6260 16210
rect 6350 15970 6590 16210
rect -5200 15640 -4960 15880
rect -4870 15640 -4630 15880
rect -4540 15640 -4300 15880
rect -4210 15640 -3970 15880
rect -3880 15640 -3640 15880
rect -3550 15640 -3310 15880
rect -3220 15640 -2980 15880
rect -2890 15640 -2650 15880
rect -2560 15640 -2320 15880
rect -2230 15640 -1990 15880
rect -1900 15640 -1660 15880
rect -1570 15640 -1330 15880
rect -1240 15640 -1000 15880
rect -910 15640 -670 15880
rect -580 15640 -340 15880
rect -250 15640 -10 15880
rect 80 15640 320 15880
rect 410 15640 650 15880
rect 740 15640 980 15880
rect 1070 15640 1310 15880
rect 1400 15640 1640 15880
rect 1730 15640 1970 15880
rect 2060 15640 2300 15880
rect 2390 15640 2630 15880
rect 2720 15640 2960 15880
rect 3050 15640 3290 15880
rect 3380 15640 3620 15880
rect 3710 15640 3950 15880
rect 4040 15640 4280 15880
rect 4370 15640 4610 15880
rect 4700 15640 4940 15880
rect 5030 15640 5270 15880
rect 5360 15640 5600 15880
rect 5690 15640 5930 15880
rect 6020 15640 6260 15880
rect 6350 15640 6590 15880
rect -5200 15310 -4960 15550
rect -4870 15310 -4630 15550
rect -4540 15310 -4300 15550
rect -4210 15310 -3970 15550
rect -3880 15310 -3640 15550
rect -3550 15310 -3310 15550
rect -3220 15310 -2980 15550
rect -2890 15310 -2650 15550
rect -2560 15310 -2320 15550
rect -2230 15310 -1990 15550
rect -1900 15310 -1660 15550
rect -1570 15310 -1330 15550
rect -1240 15310 -1000 15550
rect -910 15310 -670 15550
rect -580 15310 -340 15550
rect -250 15310 -10 15550
rect 80 15310 320 15550
rect 410 15310 650 15550
rect 740 15310 980 15550
rect 1070 15310 1310 15550
rect 1400 15310 1640 15550
rect 1730 15310 1970 15550
rect 2060 15310 2300 15550
rect 2390 15310 2630 15550
rect 2720 15310 2960 15550
rect 3050 15310 3290 15550
rect 3380 15310 3620 15550
rect 3710 15310 3950 15550
rect 4040 15310 4280 15550
rect 4370 15310 4610 15550
rect 4700 15310 4940 15550
rect 5030 15310 5270 15550
rect 5360 15310 5600 15550
rect 5690 15310 5930 15550
rect 6020 15310 6260 15550
rect 6350 15310 6590 15550
rect -5200 14980 -4960 15220
rect -4870 14980 -4630 15220
rect -4540 14980 -4300 15220
rect -4210 14980 -3970 15220
rect -3880 14980 -3640 15220
rect -3550 14980 -3310 15220
rect -3220 14980 -2980 15220
rect -2890 14980 -2650 15220
rect -2560 14980 -2320 15220
rect -2230 14980 -1990 15220
rect -1900 14980 -1660 15220
rect -1570 14980 -1330 15220
rect -1240 14980 -1000 15220
rect -910 14980 -670 15220
rect -580 14980 -340 15220
rect -250 14980 -10 15220
rect 80 14980 320 15220
rect 410 14980 650 15220
rect 740 14980 980 15220
rect 1070 14980 1310 15220
rect 1400 14980 1640 15220
rect 1730 14980 1970 15220
rect 2060 14980 2300 15220
rect 2390 14980 2630 15220
rect 2720 14980 2960 15220
rect 3050 14980 3290 15220
rect 3380 14980 3620 15220
rect 3710 14980 3950 15220
rect 4040 14980 4280 15220
rect 4370 14980 4610 15220
rect 4700 14980 4940 15220
rect 5030 14980 5270 15220
rect 5360 14980 5600 15220
rect 5690 14980 5930 15220
rect 6020 14980 6260 15220
rect 6350 14980 6590 15220
rect -5200 14650 -4960 14890
rect -4870 14650 -4630 14890
rect -4540 14650 -4300 14890
rect -4210 14650 -3970 14890
rect -3880 14650 -3640 14890
rect -3550 14650 -3310 14890
rect -3220 14650 -2980 14890
rect -2890 14650 -2650 14890
rect -2560 14650 -2320 14890
rect -2230 14650 -1990 14890
rect -1900 14650 -1660 14890
rect -1570 14650 -1330 14890
rect -1240 14650 -1000 14890
rect -910 14650 -670 14890
rect -580 14650 -340 14890
rect -250 14650 -10 14890
rect 80 14650 320 14890
rect 410 14650 650 14890
rect 740 14650 980 14890
rect 1070 14650 1310 14890
rect 1400 14650 1640 14890
rect 1730 14650 1970 14890
rect 2060 14650 2300 14890
rect 2390 14650 2630 14890
rect 2720 14650 2960 14890
rect 3050 14650 3290 14890
rect 3380 14650 3620 14890
rect 3710 14650 3950 14890
rect 4040 14650 4280 14890
rect 4370 14650 4610 14890
rect 4700 14650 4940 14890
rect 5030 14650 5270 14890
rect 5360 14650 5600 14890
rect 5690 14650 5930 14890
rect 6020 14650 6260 14890
rect 6350 14650 6590 14890
rect -5200 14320 -4960 14560
rect -4870 14320 -4630 14560
rect -4540 14320 -4300 14560
rect -4210 14320 -3970 14560
rect -3880 14320 -3640 14560
rect -3550 14320 -3310 14560
rect -3220 14320 -2980 14560
rect -2890 14320 -2650 14560
rect -2560 14320 -2320 14560
rect -2230 14320 -1990 14560
rect -1900 14320 -1660 14560
rect -1570 14320 -1330 14560
rect -1240 14320 -1000 14560
rect -910 14320 -670 14560
rect -580 14320 -340 14560
rect -250 14320 -10 14560
rect 80 14320 320 14560
rect 410 14320 650 14560
rect 740 14320 980 14560
rect 1070 14320 1310 14560
rect 1400 14320 1640 14560
rect 1730 14320 1970 14560
rect 2060 14320 2300 14560
rect 2390 14320 2630 14560
rect 2720 14320 2960 14560
rect 3050 14320 3290 14560
rect 3380 14320 3620 14560
rect 3710 14320 3950 14560
rect 4040 14320 4280 14560
rect 4370 14320 4610 14560
rect 4700 14320 4940 14560
rect 5030 14320 5270 14560
rect 5360 14320 5600 14560
rect 5690 14320 5930 14560
rect 6020 14320 6260 14560
rect 6350 14320 6590 14560
rect -5200 13990 -4960 14230
rect -4870 13990 -4630 14230
rect -4540 13990 -4300 14230
rect -4210 13990 -3970 14230
rect -3880 13990 -3640 14230
rect -3550 13990 -3310 14230
rect -3220 13990 -2980 14230
rect -2890 13990 -2650 14230
rect -2560 13990 -2320 14230
rect -2230 13990 -1990 14230
rect -1900 13990 -1660 14230
rect -1570 13990 -1330 14230
rect -1240 13990 -1000 14230
rect -910 13990 -670 14230
rect -580 13990 -340 14230
rect -250 13990 -10 14230
rect 80 13990 320 14230
rect 410 13990 650 14230
rect 740 13990 980 14230
rect 1070 13990 1310 14230
rect 1400 13990 1640 14230
rect 1730 13990 1970 14230
rect 2060 13990 2300 14230
rect 2390 13990 2630 14230
rect 2720 13990 2960 14230
rect 3050 13990 3290 14230
rect 3380 13990 3620 14230
rect 3710 13990 3950 14230
rect 4040 13990 4280 14230
rect 4370 13990 4610 14230
rect 4700 13990 4940 14230
rect 5030 13990 5270 14230
rect 5360 13990 5600 14230
rect 5690 13990 5930 14230
rect 6020 13990 6260 14230
rect 6350 13990 6590 14230
rect -5200 13660 -4960 13900
rect -4870 13660 -4630 13900
rect -4540 13660 -4300 13900
rect -4210 13660 -3970 13900
rect -3880 13660 -3640 13900
rect -3550 13660 -3310 13900
rect -3220 13660 -2980 13900
rect -2890 13660 -2650 13900
rect -2560 13660 -2320 13900
rect -2230 13660 -1990 13900
rect -1900 13660 -1660 13900
rect -1570 13660 -1330 13900
rect -1240 13660 -1000 13900
rect -910 13660 -670 13900
rect -580 13660 -340 13900
rect -250 13660 -10 13900
rect 80 13660 320 13900
rect 410 13660 650 13900
rect 740 13660 980 13900
rect 1070 13660 1310 13900
rect 1400 13660 1640 13900
rect 1730 13660 1970 13900
rect 2060 13660 2300 13900
rect 2390 13660 2630 13900
rect 2720 13660 2960 13900
rect 3050 13660 3290 13900
rect 3380 13660 3620 13900
rect 3710 13660 3950 13900
rect 4040 13660 4280 13900
rect 4370 13660 4610 13900
rect 4700 13660 4940 13900
rect 5030 13660 5270 13900
rect 5360 13660 5600 13900
rect 5690 13660 5930 13900
rect 6020 13660 6260 13900
rect 6350 13660 6590 13900
rect -5200 13330 -4960 13570
rect -4870 13330 -4630 13570
rect -4540 13330 -4300 13570
rect -4210 13330 -3970 13570
rect -3880 13330 -3640 13570
rect -3550 13330 -3310 13570
rect -3220 13330 -2980 13570
rect -2890 13330 -2650 13570
rect -2560 13330 -2320 13570
rect -2230 13330 -1990 13570
rect -1900 13330 -1660 13570
rect -1570 13330 -1330 13570
rect -1240 13330 -1000 13570
rect -910 13330 -670 13570
rect -580 13330 -340 13570
rect -250 13330 -10 13570
rect 80 13330 320 13570
rect 410 13330 650 13570
rect 740 13330 980 13570
rect 1070 13330 1310 13570
rect 1400 13330 1640 13570
rect 1730 13330 1970 13570
rect 2060 13330 2300 13570
rect 2390 13330 2630 13570
rect 2720 13330 2960 13570
rect 3050 13330 3290 13570
rect 3380 13330 3620 13570
rect 3710 13330 3950 13570
rect 4040 13330 4280 13570
rect 4370 13330 4610 13570
rect 4700 13330 4940 13570
rect 5030 13330 5270 13570
rect 5360 13330 5600 13570
rect 5690 13330 5930 13570
rect 6020 13330 6260 13570
rect 6350 13330 6590 13570
rect -5200 13000 -4960 13240
rect -4870 13000 -4630 13240
rect -4540 13000 -4300 13240
rect -4210 13000 -3970 13240
rect -3880 13000 -3640 13240
rect -3550 13000 -3310 13240
rect -3220 13000 -2980 13240
rect -2890 13000 -2650 13240
rect -2560 13000 -2320 13240
rect -2230 13000 -1990 13240
rect -1900 13000 -1660 13240
rect -1570 13000 -1330 13240
rect -1240 13000 -1000 13240
rect -910 13000 -670 13240
rect -580 13000 -340 13240
rect -250 13000 -10 13240
rect 80 13000 320 13240
rect 410 13000 650 13240
rect 740 13000 980 13240
rect 1070 13000 1310 13240
rect 1400 13000 1640 13240
rect 1730 13000 1970 13240
rect 2060 13000 2300 13240
rect 2390 13000 2630 13240
rect 2720 13000 2960 13240
rect 3050 13000 3290 13240
rect 3380 13000 3620 13240
rect 3710 13000 3950 13240
rect 4040 13000 4280 13240
rect 4370 13000 4610 13240
rect 4700 13000 4940 13240
rect 5030 13000 5270 13240
rect 5360 13000 5600 13240
rect 5690 13000 5930 13240
rect 6020 13000 6260 13240
rect 6350 13000 6590 13240
rect -5200 12670 -4960 12910
rect -4870 12670 -4630 12910
rect -4540 12670 -4300 12910
rect -4210 12670 -3970 12910
rect -3880 12670 -3640 12910
rect -3550 12670 -3310 12910
rect -3220 12670 -2980 12910
rect -2890 12670 -2650 12910
rect -2560 12670 -2320 12910
rect -2230 12670 -1990 12910
rect -1900 12670 -1660 12910
rect -1570 12670 -1330 12910
rect -1240 12670 -1000 12910
rect -910 12670 -670 12910
rect -580 12670 -340 12910
rect -250 12670 -10 12910
rect 80 12670 320 12910
rect 410 12670 650 12910
rect 740 12670 980 12910
rect 1070 12670 1310 12910
rect 1400 12670 1640 12910
rect 1730 12670 1970 12910
rect 2060 12670 2300 12910
rect 2390 12670 2630 12910
rect 2720 12670 2960 12910
rect 3050 12670 3290 12910
rect 3380 12670 3620 12910
rect 3710 12670 3950 12910
rect 4040 12670 4280 12910
rect 4370 12670 4610 12910
rect 4700 12670 4940 12910
rect 5030 12670 5270 12910
rect 5360 12670 5600 12910
rect 5690 12670 5930 12910
rect 6020 12670 6260 12910
rect 6350 12670 6590 12910
rect -5200 12340 -4960 12580
rect -4870 12340 -4630 12580
rect -4540 12340 -4300 12580
rect -4210 12340 -3970 12580
rect -3880 12340 -3640 12580
rect -3550 12340 -3310 12580
rect -3220 12340 -2980 12580
rect -2890 12340 -2650 12580
rect -2560 12340 -2320 12580
rect -2230 12340 -1990 12580
rect -1900 12340 -1660 12580
rect -1570 12340 -1330 12580
rect -1240 12340 -1000 12580
rect -910 12340 -670 12580
rect -580 12340 -340 12580
rect -250 12340 -10 12580
rect 80 12340 320 12580
rect 410 12340 650 12580
rect 740 12340 980 12580
rect 1070 12340 1310 12580
rect 1400 12340 1640 12580
rect 1730 12340 1970 12580
rect 2060 12340 2300 12580
rect 2390 12340 2630 12580
rect 2720 12340 2960 12580
rect 3050 12340 3290 12580
rect 3380 12340 3620 12580
rect 3710 12340 3950 12580
rect 4040 12340 4280 12580
rect 4370 12340 4610 12580
rect 4700 12340 4940 12580
rect 5030 12340 5270 12580
rect 5360 12340 5600 12580
rect 5690 12340 5930 12580
rect 6020 12340 6260 12580
rect 6350 12340 6590 12580
rect -5200 12010 -4960 12250
rect -4870 12010 -4630 12250
rect -4540 12010 -4300 12250
rect -4210 12010 -3970 12250
rect -3880 12010 -3640 12250
rect -3550 12010 -3310 12250
rect -3220 12010 -2980 12250
rect -2890 12010 -2650 12250
rect -2560 12010 -2320 12250
rect -2230 12010 -1990 12250
rect -1900 12010 -1660 12250
rect -1570 12010 -1330 12250
rect -1240 12010 -1000 12250
rect -910 12010 -670 12250
rect -580 12010 -340 12250
rect -250 12010 -10 12250
rect 80 12010 320 12250
rect 410 12010 650 12250
rect 740 12010 980 12250
rect 1070 12010 1310 12250
rect 1400 12010 1640 12250
rect 1730 12010 1970 12250
rect 2060 12010 2300 12250
rect 2390 12010 2630 12250
rect 2720 12010 2960 12250
rect 3050 12010 3290 12250
rect 3380 12010 3620 12250
rect 3710 12010 3950 12250
rect 4040 12010 4280 12250
rect 4370 12010 4610 12250
rect 4700 12010 4940 12250
rect 5030 12010 5270 12250
rect 5360 12010 5600 12250
rect 5690 12010 5930 12250
rect 6020 12010 6260 12250
rect 6350 12010 6590 12250
rect -5200 11680 -4960 11920
rect -4870 11680 -4630 11920
rect -4540 11680 -4300 11920
rect -4210 11680 -3970 11920
rect -3880 11680 -3640 11920
rect -3550 11680 -3310 11920
rect -3220 11680 -2980 11920
rect -2890 11680 -2650 11920
rect -2560 11680 -2320 11920
rect -2230 11680 -1990 11920
rect -1900 11680 -1660 11920
rect -1570 11680 -1330 11920
rect -1240 11680 -1000 11920
rect -910 11680 -670 11920
rect -580 11680 -340 11920
rect -250 11680 -10 11920
rect 80 11680 320 11920
rect 410 11680 650 11920
rect 740 11680 980 11920
rect 1070 11680 1310 11920
rect 1400 11680 1640 11920
rect 1730 11680 1970 11920
rect 2060 11680 2300 11920
rect 2390 11680 2630 11920
rect 2720 11680 2960 11920
rect 3050 11680 3290 11920
rect 3380 11680 3620 11920
rect 3710 11680 3950 11920
rect 4040 11680 4280 11920
rect 4370 11680 4610 11920
rect 4700 11680 4940 11920
rect 5030 11680 5270 11920
rect 5360 11680 5600 11920
rect 5690 11680 5930 11920
rect 6020 11680 6260 11920
rect 6350 11680 6590 11920
rect -5200 11350 -4960 11590
rect -4870 11350 -4630 11590
rect -4540 11350 -4300 11590
rect -4210 11350 -3970 11590
rect -3880 11350 -3640 11590
rect -3550 11350 -3310 11590
rect -3220 11350 -2980 11590
rect -2890 11350 -2650 11590
rect -2560 11350 -2320 11590
rect -2230 11350 -1990 11590
rect -1900 11350 -1660 11590
rect -1570 11350 -1330 11590
rect -1240 11350 -1000 11590
rect -910 11350 -670 11590
rect -580 11350 -340 11590
rect -250 11350 -10 11590
rect 80 11350 320 11590
rect 410 11350 650 11590
rect 740 11350 980 11590
rect 1070 11350 1310 11590
rect 1400 11350 1640 11590
rect 1730 11350 1970 11590
rect 2060 11350 2300 11590
rect 2390 11350 2630 11590
rect 2720 11350 2960 11590
rect 3050 11350 3290 11590
rect 3380 11350 3620 11590
rect 3710 11350 3950 11590
rect 4040 11350 4280 11590
rect 4370 11350 4610 11590
rect 4700 11350 4940 11590
rect 5030 11350 5270 11590
rect 5360 11350 5600 11590
rect 5690 11350 5930 11590
rect 6020 11350 6260 11590
rect 6350 11350 6590 11590
rect -5200 11020 -4960 11260
rect -4870 11020 -4630 11260
rect -4540 11020 -4300 11260
rect -4210 11020 -3970 11260
rect -3880 11020 -3640 11260
rect -3550 11020 -3310 11260
rect -3220 11020 -2980 11260
rect -2890 11020 -2650 11260
rect -2560 11020 -2320 11260
rect -2230 11020 -1990 11260
rect -1900 11020 -1660 11260
rect -1570 11020 -1330 11260
rect -1240 11020 -1000 11260
rect -910 11020 -670 11260
rect -580 11020 -340 11260
rect -250 11020 -10 11260
rect 80 11020 320 11260
rect 410 11020 650 11260
rect 740 11020 980 11260
rect 1070 11020 1310 11260
rect 1400 11020 1640 11260
rect 1730 11020 1970 11260
rect 2060 11020 2300 11260
rect 2390 11020 2630 11260
rect 2720 11020 2960 11260
rect 3050 11020 3290 11260
rect 3380 11020 3620 11260
rect 3710 11020 3950 11260
rect 4040 11020 4280 11260
rect 4370 11020 4610 11260
rect 4700 11020 4940 11260
rect 5030 11020 5270 11260
rect 5360 11020 5600 11260
rect 5690 11020 5930 11260
rect 6020 11020 6260 11260
rect 6350 11020 6590 11260
rect -5200 10690 -4960 10930
rect -4870 10690 -4630 10930
rect -4540 10690 -4300 10930
rect -4210 10690 -3970 10930
rect -3880 10690 -3640 10930
rect -3550 10690 -3310 10930
rect -3220 10690 -2980 10930
rect -2890 10690 -2650 10930
rect -2560 10690 -2320 10930
rect -2230 10690 -1990 10930
rect -1900 10690 -1660 10930
rect -1570 10690 -1330 10930
rect -1240 10690 -1000 10930
rect -910 10690 -670 10930
rect -580 10690 -340 10930
rect -250 10690 -10 10930
rect 80 10690 320 10930
rect 410 10690 650 10930
rect 740 10690 980 10930
rect 1070 10690 1310 10930
rect 1400 10690 1640 10930
rect 1730 10690 1970 10930
rect 2060 10690 2300 10930
rect 2390 10690 2630 10930
rect 2720 10690 2960 10930
rect 3050 10690 3290 10930
rect 3380 10690 3620 10930
rect 3710 10690 3950 10930
rect 4040 10690 4280 10930
rect 4370 10690 4610 10930
rect 4700 10690 4940 10930
rect 5030 10690 5270 10930
rect 5360 10690 5600 10930
rect 5690 10690 5930 10930
rect 6020 10690 6260 10930
rect 6350 10690 6590 10930
rect -5200 10360 -4960 10600
rect -4870 10360 -4630 10600
rect -4540 10360 -4300 10600
rect -4210 10360 -3970 10600
rect -3880 10360 -3640 10600
rect -3550 10360 -3310 10600
rect -3220 10360 -2980 10600
rect -2890 10360 -2650 10600
rect -2560 10360 -2320 10600
rect -2230 10360 -1990 10600
rect -1900 10360 -1660 10600
rect -1570 10360 -1330 10600
rect -1240 10360 -1000 10600
rect -910 10360 -670 10600
rect -580 10360 -340 10600
rect -250 10360 -10 10600
rect 80 10360 320 10600
rect 410 10360 650 10600
rect 740 10360 980 10600
rect 1070 10360 1310 10600
rect 1400 10360 1640 10600
rect 1730 10360 1970 10600
rect 2060 10360 2300 10600
rect 2390 10360 2630 10600
rect 2720 10360 2960 10600
rect 3050 10360 3290 10600
rect 3380 10360 3620 10600
rect 3710 10360 3950 10600
rect 4040 10360 4280 10600
rect 4370 10360 4610 10600
rect 4700 10360 4940 10600
rect 5030 10360 5270 10600
rect 5360 10360 5600 10600
rect 5690 10360 5930 10600
rect 6020 10360 6260 10600
rect 6350 10360 6590 10600
rect -5200 10030 -4960 10270
rect -4870 10030 -4630 10270
rect -4540 10030 -4300 10270
rect -4210 10030 -3970 10270
rect -3880 10030 -3640 10270
rect -3550 10030 -3310 10270
rect -3220 10030 -2980 10270
rect -2890 10030 -2650 10270
rect -2560 10030 -2320 10270
rect -2230 10030 -1990 10270
rect -1900 10030 -1660 10270
rect -1570 10030 -1330 10270
rect -1240 10030 -1000 10270
rect -910 10030 -670 10270
rect -580 10030 -340 10270
rect -250 10030 -10 10270
rect 80 10030 320 10270
rect 410 10030 650 10270
rect 740 10030 980 10270
rect 1070 10030 1310 10270
rect 1400 10030 1640 10270
rect 1730 10030 1970 10270
rect 2060 10030 2300 10270
rect 2390 10030 2630 10270
rect 2720 10030 2960 10270
rect 3050 10030 3290 10270
rect 3380 10030 3620 10270
rect 3710 10030 3950 10270
rect 4040 10030 4280 10270
rect 4370 10030 4610 10270
rect 4700 10030 4940 10270
rect 5030 10030 5270 10270
rect 5360 10030 5600 10270
rect 5690 10030 5930 10270
rect 6020 10030 6260 10270
rect 6350 10030 6590 10270
rect -5200 9700 -4960 9940
rect -4870 9700 -4630 9940
rect -4540 9700 -4300 9940
rect -4210 9700 -3970 9940
rect -3880 9700 -3640 9940
rect -3550 9700 -3310 9940
rect -3220 9700 -2980 9940
rect -2890 9700 -2650 9940
rect -2560 9700 -2320 9940
rect -2230 9700 -1990 9940
rect -1900 9700 -1660 9940
rect -1570 9700 -1330 9940
rect -1240 9700 -1000 9940
rect -910 9700 -670 9940
rect -580 9700 -340 9940
rect -250 9700 -10 9940
rect 80 9700 320 9940
rect 410 9700 650 9940
rect 740 9700 980 9940
rect 1070 9700 1310 9940
rect 1400 9700 1640 9940
rect 1730 9700 1970 9940
rect 2060 9700 2300 9940
rect 2390 9700 2630 9940
rect 2720 9700 2960 9940
rect 3050 9700 3290 9940
rect 3380 9700 3620 9940
rect 3710 9700 3950 9940
rect 4040 9700 4280 9940
rect 4370 9700 4610 9940
rect 4700 9700 4940 9940
rect 5030 9700 5270 9940
rect 5360 9700 5600 9940
rect 5690 9700 5930 9940
rect 6020 9700 6260 9940
rect 6350 9700 6590 9940
rect -5200 9370 -4960 9610
rect -4870 9370 -4630 9610
rect -4540 9370 -4300 9610
rect -4210 9370 -3970 9610
rect -3880 9370 -3640 9610
rect -3550 9370 -3310 9610
rect -3220 9370 -2980 9610
rect -2890 9370 -2650 9610
rect -2560 9370 -2320 9610
rect -2230 9370 -1990 9610
rect -1900 9370 -1660 9610
rect -1570 9370 -1330 9610
rect -1240 9370 -1000 9610
rect -910 9370 -670 9610
rect -580 9370 -340 9610
rect -250 9370 -10 9610
rect 80 9370 320 9610
rect 410 9370 650 9610
rect 740 9370 980 9610
rect 1070 9370 1310 9610
rect 1400 9370 1640 9610
rect 1730 9370 1970 9610
rect 2060 9370 2300 9610
rect 2390 9370 2630 9610
rect 2720 9370 2960 9610
rect 3050 9370 3290 9610
rect 3380 9370 3620 9610
rect 3710 9370 3950 9610
rect 4040 9370 4280 9610
rect 4370 9370 4610 9610
rect 4700 9370 4940 9610
rect 5030 9370 5270 9610
rect 5360 9370 5600 9610
rect 5690 9370 5930 9610
rect 6020 9370 6260 9610
rect 6350 9370 6590 9610
rect -5200 9040 -4960 9280
rect -4870 9040 -4630 9280
rect -4540 9040 -4300 9280
rect -4210 9040 -3970 9280
rect -3880 9040 -3640 9280
rect -3550 9040 -3310 9280
rect -3220 9040 -2980 9280
rect -2890 9040 -2650 9280
rect -2560 9040 -2320 9280
rect -2230 9040 -1990 9280
rect -1900 9040 -1660 9280
rect -1570 9040 -1330 9280
rect -1240 9040 -1000 9280
rect -910 9040 -670 9280
rect -580 9040 -340 9280
rect -250 9040 -10 9280
rect 80 9040 320 9280
rect 410 9040 650 9280
rect 740 9040 980 9280
rect 1070 9040 1310 9280
rect 1400 9040 1640 9280
rect 1730 9040 1970 9280
rect 2060 9040 2300 9280
rect 2390 9040 2630 9280
rect 2720 9040 2960 9280
rect 3050 9040 3290 9280
rect 3380 9040 3620 9280
rect 3710 9040 3950 9280
rect 4040 9040 4280 9280
rect 4370 9040 4610 9280
rect 4700 9040 4940 9280
rect 5030 9040 5270 9280
rect 5360 9040 5600 9280
rect 5690 9040 5930 9280
rect 6020 9040 6260 9280
rect 6350 9040 6590 9280
rect 8310 20590 8550 20830
rect 8640 20590 8880 20830
rect 8970 20590 9210 20830
rect 9300 20590 9540 20830
rect 9630 20590 9870 20830
rect 9960 20590 10200 20830
rect 10290 20590 10530 20830
rect 10620 20590 10860 20830
rect 10950 20590 11190 20830
rect 11280 20590 11520 20830
rect 11610 20590 11850 20830
rect 11940 20590 12180 20830
rect 12270 20590 12510 20830
rect 12600 20590 12840 20830
rect 12930 20590 13170 20830
rect 13260 20590 13500 20830
rect 13590 20590 13830 20830
rect 13920 20590 14160 20830
rect 14250 20590 14490 20830
rect 14580 20590 14820 20830
rect 14910 20590 15150 20830
rect 15240 20590 15480 20830
rect 15570 20590 15810 20830
rect 15900 20590 16140 20830
rect 16230 20590 16470 20830
rect 16560 20590 16800 20830
rect 16890 20590 17130 20830
rect 17220 20590 17460 20830
rect 17550 20590 17790 20830
rect 17880 20590 18120 20830
rect 18210 20590 18450 20830
rect 18540 20590 18780 20830
rect 18870 20590 19110 20830
rect 19200 20590 19440 20830
rect 19530 20590 19770 20830
rect 19860 20590 20100 20830
rect 8310 20260 8550 20500
rect 8640 20260 8880 20500
rect 8970 20260 9210 20500
rect 9300 20260 9540 20500
rect 9630 20260 9870 20500
rect 9960 20260 10200 20500
rect 10290 20260 10530 20500
rect 10620 20260 10860 20500
rect 10950 20260 11190 20500
rect 11280 20260 11520 20500
rect 11610 20260 11850 20500
rect 11940 20260 12180 20500
rect 12270 20260 12510 20500
rect 12600 20260 12840 20500
rect 12930 20260 13170 20500
rect 13260 20260 13500 20500
rect 13590 20260 13830 20500
rect 13920 20260 14160 20500
rect 14250 20260 14490 20500
rect 14580 20260 14820 20500
rect 14910 20260 15150 20500
rect 15240 20260 15480 20500
rect 15570 20260 15810 20500
rect 15900 20260 16140 20500
rect 16230 20260 16470 20500
rect 16560 20260 16800 20500
rect 16890 20260 17130 20500
rect 17220 20260 17460 20500
rect 17550 20260 17790 20500
rect 17880 20260 18120 20500
rect 18210 20260 18450 20500
rect 18540 20260 18780 20500
rect 18870 20260 19110 20500
rect 19200 20260 19440 20500
rect 19530 20260 19770 20500
rect 19860 20260 20100 20500
rect 8310 19930 8550 20170
rect 8640 19930 8880 20170
rect 8970 19930 9210 20170
rect 9300 19930 9540 20170
rect 9630 19930 9870 20170
rect 9960 19930 10200 20170
rect 10290 19930 10530 20170
rect 10620 19930 10860 20170
rect 10950 19930 11190 20170
rect 11280 19930 11520 20170
rect 11610 19930 11850 20170
rect 11940 19930 12180 20170
rect 12270 19930 12510 20170
rect 12600 19930 12840 20170
rect 12930 19930 13170 20170
rect 13260 19930 13500 20170
rect 13590 19930 13830 20170
rect 13920 19930 14160 20170
rect 14250 19930 14490 20170
rect 14580 19930 14820 20170
rect 14910 19930 15150 20170
rect 15240 19930 15480 20170
rect 15570 19930 15810 20170
rect 15900 19930 16140 20170
rect 16230 19930 16470 20170
rect 16560 19930 16800 20170
rect 16890 19930 17130 20170
rect 17220 19930 17460 20170
rect 17550 19930 17790 20170
rect 17880 19930 18120 20170
rect 18210 19930 18450 20170
rect 18540 19930 18780 20170
rect 18870 19930 19110 20170
rect 19200 19930 19440 20170
rect 19530 19930 19770 20170
rect 19860 19930 20100 20170
rect 8310 19600 8550 19840
rect 8640 19600 8880 19840
rect 8970 19600 9210 19840
rect 9300 19600 9540 19840
rect 9630 19600 9870 19840
rect 9960 19600 10200 19840
rect 10290 19600 10530 19840
rect 10620 19600 10860 19840
rect 10950 19600 11190 19840
rect 11280 19600 11520 19840
rect 11610 19600 11850 19840
rect 11940 19600 12180 19840
rect 12270 19600 12510 19840
rect 12600 19600 12840 19840
rect 12930 19600 13170 19840
rect 13260 19600 13500 19840
rect 13590 19600 13830 19840
rect 13920 19600 14160 19840
rect 14250 19600 14490 19840
rect 14580 19600 14820 19840
rect 14910 19600 15150 19840
rect 15240 19600 15480 19840
rect 15570 19600 15810 19840
rect 15900 19600 16140 19840
rect 16230 19600 16470 19840
rect 16560 19600 16800 19840
rect 16890 19600 17130 19840
rect 17220 19600 17460 19840
rect 17550 19600 17790 19840
rect 17880 19600 18120 19840
rect 18210 19600 18450 19840
rect 18540 19600 18780 19840
rect 18870 19600 19110 19840
rect 19200 19600 19440 19840
rect 19530 19600 19770 19840
rect 19860 19600 20100 19840
rect 8310 19270 8550 19510
rect 8640 19270 8880 19510
rect 8970 19270 9210 19510
rect 9300 19270 9540 19510
rect 9630 19270 9870 19510
rect 9960 19270 10200 19510
rect 10290 19270 10530 19510
rect 10620 19270 10860 19510
rect 10950 19270 11190 19510
rect 11280 19270 11520 19510
rect 11610 19270 11850 19510
rect 11940 19270 12180 19510
rect 12270 19270 12510 19510
rect 12600 19270 12840 19510
rect 12930 19270 13170 19510
rect 13260 19270 13500 19510
rect 13590 19270 13830 19510
rect 13920 19270 14160 19510
rect 14250 19270 14490 19510
rect 14580 19270 14820 19510
rect 14910 19270 15150 19510
rect 15240 19270 15480 19510
rect 15570 19270 15810 19510
rect 15900 19270 16140 19510
rect 16230 19270 16470 19510
rect 16560 19270 16800 19510
rect 16890 19270 17130 19510
rect 17220 19270 17460 19510
rect 17550 19270 17790 19510
rect 17880 19270 18120 19510
rect 18210 19270 18450 19510
rect 18540 19270 18780 19510
rect 18870 19270 19110 19510
rect 19200 19270 19440 19510
rect 19530 19270 19770 19510
rect 19860 19270 20100 19510
rect 8310 18940 8550 19180
rect 8640 18940 8880 19180
rect 8970 18940 9210 19180
rect 9300 18940 9540 19180
rect 9630 18940 9870 19180
rect 9960 18940 10200 19180
rect 10290 18940 10530 19180
rect 10620 18940 10860 19180
rect 10950 18940 11190 19180
rect 11280 18940 11520 19180
rect 11610 18940 11850 19180
rect 11940 18940 12180 19180
rect 12270 18940 12510 19180
rect 12600 18940 12840 19180
rect 12930 18940 13170 19180
rect 13260 18940 13500 19180
rect 13590 18940 13830 19180
rect 13920 18940 14160 19180
rect 14250 18940 14490 19180
rect 14580 18940 14820 19180
rect 14910 18940 15150 19180
rect 15240 18940 15480 19180
rect 15570 18940 15810 19180
rect 15900 18940 16140 19180
rect 16230 18940 16470 19180
rect 16560 18940 16800 19180
rect 16890 18940 17130 19180
rect 17220 18940 17460 19180
rect 17550 18940 17790 19180
rect 17880 18940 18120 19180
rect 18210 18940 18450 19180
rect 18540 18940 18780 19180
rect 18870 18940 19110 19180
rect 19200 18940 19440 19180
rect 19530 18940 19770 19180
rect 19860 18940 20100 19180
rect 8310 18610 8550 18850
rect 8640 18610 8880 18850
rect 8970 18610 9210 18850
rect 9300 18610 9540 18850
rect 9630 18610 9870 18850
rect 9960 18610 10200 18850
rect 10290 18610 10530 18850
rect 10620 18610 10860 18850
rect 10950 18610 11190 18850
rect 11280 18610 11520 18850
rect 11610 18610 11850 18850
rect 11940 18610 12180 18850
rect 12270 18610 12510 18850
rect 12600 18610 12840 18850
rect 12930 18610 13170 18850
rect 13260 18610 13500 18850
rect 13590 18610 13830 18850
rect 13920 18610 14160 18850
rect 14250 18610 14490 18850
rect 14580 18610 14820 18850
rect 14910 18610 15150 18850
rect 15240 18610 15480 18850
rect 15570 18610 15810 18850
rect 15900 18610 16140 18850
rect 16230 18610 16470 18850
rect 16560 18610 16800 18850
rect 16890 18610 17130 18850
rect 17220 18610 17460 18850
rect 17550 18610 17790 18850
rect 17880 18610 18120 18850
rect 18210 18610 18450 18850
rect 18540 18610 18780 18850
rect 18870 18610 19110 18850
rect 19200 18610 19440 18850
rect 19530 18610 19770 18850
rect 19860 18610 20100 18850
rect 8310 18280 8550 18520
rect 8640 18280 8880 18520
rect 8970 18280 9210 18520
rect 9300 18280 9540 18520
rect 9630 18280 9870 18520
rect 9960 18280 10200 18520
rect 10290 18280 10530 18520
rect 10620 18280 10860 18520
rect 10950 18280 11190 18520
rect 11280 18280 11520 18520
rect 11610 18280 11850 18520
rect 11940 18280 12180 18520
rect 12270 18280 12510 18520
rect 12600 18280 12840 18520
rect 12930 18280 13170 18520
rect 13260 18280 13500 18520
rect 13590 18280 13830 18520
rect 13920 18280 14160 18520
rect 14250 18280 14490 18520
rect 14580 18280 14820 18520
rect 14910 18280 15150 18520
rect 15240 18280 15480 18520
rect 15570 18280 15810 18520
rect 15900 18280 16140 18520
rect 16230 18280 16470 18520
rect 16560 18280 16800 18520
rect 16890 18280 17130 18520
rect 17220 18280 17460 18520
rect 17550 18280 17790 18520
rect 17880 18280 18120 18520
rect 18210 18280 18450 18520
rect 18540 18280 18780 18520
rect 18870 18280 19110 18520
rect 19200 18280 19440 18520
rect 19530 18280 19770 18520
rect 19860 18280 20100 18520
rect 8310 17950 8550 18190
rect 8640 17950 8880 18190
rect 8970 17950 9210 18190
rect 9300 17950 9540 18190
rect 9630 17950 9870 18190
rect 9960 17950 10200 18190
rect 10290 17950 10530 18190
rect 10620 17950 10860 18190
rect 10950 17950 11190 18190
rect 11280 17950 11520 18190
rect 11610 17950 11850 18190
rect 11940 17950 12180 18190
rect 12270 17950 12510 18190
rect 12600 17950 12840 18190
rect 12930 17950 13170 18190
rect 13260 17950 13500 18190
rect 13590 17950 13830 18190
rect 13920 17950 14160 18190
rect 14250 17950 14490 18190
rect 14580 17950 14820 18190
rect 14910 17950 15150 18190
rect 15240 17950 15480 18190
rect 15570 17950 15810 18190
rect 15900 17950 16140 18190
rect 16230 17950 16470 18190
rect 16560 17950 16800 18190
rect 16890 17950 17130 18190
rect 17220 17950 17460 18190
rect 17550 17950 17790 18190
rect 17880 17950 18120 18190
rect 18210 17950 18450 18190
rect 18540 17950 18780 18190
rect 18870 17950 19110 18190
rect 19200 17950 19440 18190
rect 19530 17950 19770 18190
rect 19860 17950 20100 18190
rect 8310 17620 8550 17860
rect 8640 17620 8880 17860
rect 8970 17620 9210 17860
rect 9300 17620 9540 17860
rect 9630 17620 9870 17860
rect 9960 17620 10200 17860
rect 10290 17620 10530 17860
rect 10620 17620 10860 17860
rect 10950 17620 11190 17860
rect 11280 17620 11520 17860
rect 11610 17620 11850 17860
rect 11940 17620 12180 17860
rect 12270 17620 12510 17860
rect 12600 17620 12840 17860
rect 12930 17620 13170 17860
rect 13260 17620 13500 17860
rect 13590 17620 13830 17860
rect 13920 17620 14160 17860
rect 14250 17620 14490 17860
rect 14580 17620 14820 17860
rect 14910 17620 15150 17860
rect 15240 17620 15480 17860
rect 15570 17620 15810 17860
rect 15900 17620 16140 17860
rect 16230 17620 16470 17860
rect 16560 17620 16800 17860
rect 16890 17620 17130 17860
rect 17220 17620 17460 17860
rect 17550 17620 17790 17860
rect 17880 17620 18120 17860
rect 18210 17620 18450 17860
rect 18540 17620 18780 17860
rect 18870 17620 19110 17860
rect 19200 17620 19440 17860
rect 19530 17620 19770 17860
rect 19860 17620 20100 17860
rect 8310 17290 8550 17530
rect 8640 17290 8880 17530
rect 8970 17290 9210 17530
rect 9300 17290 9540 17530
rect 9630 17290 9870 17530
rect 9960 17290 10200 17530
rect 10290 17290 10530 17530
rect 10620 17290 10860 17530
rect 10950 17290 11190 17530
rect 11280 17290 11520 17530
rect 11610 17290 11850 17530
rect 11940 17290 12180 17530
rect 12270 17290 12510 17530
rect 12600 17290 12840 17530
rect 12930 17290 13170 17530
rect 13260 17290 13500 17530
rect 13590 17290 13830 17530
rect 13920 17290 14160 17530
rect 14250 17290 14490 17530
rect 14580 17290 14820 17530
rect 14910 17290 15150 17530
rect 15240 17290 15480 17530
rect 15570 17290 15810 17530
rect 15900 17290 16140 17530
rect 16230 17290 16470 17530
rect 16560 17290 16800 17530
rect 16890 17290 17130 17530
rect 17220 17290 17460 17530
rect 17550 17290 17790 17530
rect 17880 17290 18120 17530
rect 18210 17290 18450 17530
rect 18540 17290 18780 17530
rect 18870 17290 19110 17530
rect 19200 17290 19440 17530
rect 19530 17290 19770 17530
rect 19860 17290 20100 17530
rect 8310 16960 8550 17200
rect 8640 16960 8880 17200
rect 8970 16960 9210 17200
rect 9300 16960 9540 17200
rect 9630 16960 9870 17200
rect 9960 16960 10200 17200
rect 10290 16960 10530 17200
rect 10620 16960 10860 17200
rect 10950 16960 11190 17200
rect 11280 16960 11520 17200
rect 11610 16960 11850 17200
rect 11940 16960 12180 17200
rect 12270 16960 12510 17200
rect 12600 16960 12840 17200
rect 12930 16960 13170 17200
rect 13260 16960 13500 17200
rect 13590 16960 13830 17200
rect 13920 16960 14160 17200
rect 14250 16960 14490 17200
rect 14580 16960 14820 17200
rect 14910 16960 15150 17200
rect 15240 16960 15480 17200
rect 15570 16960 15810 17200
rect 15900 16960 16140 17200
rect 16230 16960 16470 17200
rect 16560 16960 16800 17200
rect 16890 16960 17130 17200
rect 17220 16960 17460 17200
rect 17550 16960 17790 17200
rect 17880 16960 18120 17200
rect 18210 16960 18450 17200
rect 18540 16960 18780 17200
rect 18870 16960 19110 17200
rect 19200 16960 19440 17200
rect 19530 16960 19770 17200
rect 19860 16960 20100 17200
rect 8310 16630 8550 16870
rect 8640 16630 8880 16870
rect 8970 16630 9210 16870
rect 9300 16630 9540 16870
rect 9630 16630 9870 16870
rect 9960 16630 10200 16870
rect 10290 16630 10530 16870
rect 10620 16630 10860 16870
rect 10950 16630 11190 16870
rect 11280 16630 11520 16870
rect 11610 16630 11850 16870
rect 11940 16630 12180 16870
rect 12270 16630 12510 16870
rect 12600 16630 12840 16870
rect 12930 16630 13170 16870
rect 13260 16630 13500 16870
rect 13590 16630 13830 16870
rect 13920 16630 14160 16870
rect 14250 16630 14490 16870
rect 14580 16630 14820 16870
rect 14910 16630 15150 16870
rect 15240 16630 15480 16870
rect 15570 16630 15810 16870
rect 15900 16630 16140 16870
rect 16230 16630 16470 16870
rect 16560 16630 16800 16870
rect 16890 16630 17130 16870
rect 17220 16630 17460 16870
rect 17550 16630 17790 16870
rect 17880 16630 18120 16870
rect 18210 16630 18450 16870
rect 18540 16630 18780 16870
rect 18870 16630 19110 16870
rect 19200 16630 19440 16870
rect 19530 16630 19770 16870
rect 19860 16630 20100 16870
rect 8310 16300 8550 16540
rect 8640 16300 8880 16540
rect 8970 16300 9210 16540
rect 9300 16300 9540 16540
rect 9630 16300 9870 16540
rect 9960 16300 10200 16540
rect 10290 16300 10530 16540
rect 10620 16300 10860 16540
rect 10950 16300 11190 16540
rect 11280 16300 11520 16540
rect 11610 16300 11850 16540
rect 11940 16300 12180 16540
rect 12270 16300 12510 16540
rect 12600 16300 12840 16540
rect 12930 16300 13170 16540
rect 13260 16300 13500 16540
rect 13590 16300 13830 16540
rect 13920 16300 14160 16540
rect 14250 16300 14490 16540
rect 14580 16300 14820 16540
rect 14910 16300 15150 16540
rect 15240 16300 15480 16540
rect 15570 16300 15810 16540
rect 15900 16300 16140 16540
rect 16230 16300 16470 16540
rect 16560 16300 16800 16540
rect 16890 16300 17130 16540
rect 17220 16300 17460 16540
rect 17550 16300 17790 16540
rect 17880 16300 18120 16540
rect 18210 16300 18450 16540
rect 18540 16300 18780 16540
rect 18870 16300 19110 16540
rect 19200 16300 19440 16540
rect 19530 16300 19770 16540
rect 19860 16300 20100 16540
rect 8310 15970 8550 16210
rect 8640 15970 8880 16210
rect 8970 15970 9210 16210
rect 9300 15970 9540 16210
rect 9630 15970 9870 16210
rect 9960 15970 10200 16210
rect 10290 15970 10530 16210
rect 10620 15970 10860 16210
rect 10950 15970 11190 16210
rect 11280 15970 11520 16210
rect 11610 15970 11850 16210
rect 11940 15970 12180 16210
rect 12270 15970 12510 16210
rect 12600 15970 12840 16210
rect 12930 15970 13170 16210
rect 13260 15970 13500 16210
rect 13590 15970 13830 16210
rect 13920 15970 14160 16210
rect 14250 15970 14490 16210
rect 14580 15970 14820 16210
rect 14910 15970 15150 16210
rect 15240 15970 15480 16210
rect 15570 15970 15810 16210
rect 15900 15970 16140 16210
rect 16230 15970 16470 16210
rect 16560 15970 16800 16210
rect 16890 15970 17130 16210
rect 17220 15970 17460 16210
rect 17550 15970 17790 16210
rect 17880 15970 18120 16210
rect 18210 15970 18450 16210
rect 18540 15970 18780 16210
rect 18870 15970 19110 16210
rect 19200 15970 19440 16210
rect 19530 15970 19770 16210
rect 19860 15970 20100 16210
rect 8310 15640 8550 15880
rect 8640 15640 8880 15880
rect 8970 15640 9210 15880
rect 9300 15640 9540 15880
rect 9630 15640 9870 15880
rect 9960 15640 10200 15880
rect 10290 15640 10530 15880
rect 10620 15640 10860 15880
rect 10950 15640 11190 15880
rect 11280 15640 11520 15880
rect 11610 15640 11850 15880
rect 11940 15640 12180 15880
rect 12270 15640 12510 15880
rect 12600 15640 12840 15880
rect 12930 15640 13170 15880
rect 13260 15640 13500 15880
rect 13590 15640 13830 15880
rect 13920 15640 14160 15880
rect 14250 15640 14490 15880
rect 14580 15640 14820 15880
rect 14910 15640 15150 15880
rect 15240 15640 15480 15880
rect 15570 15640 15810 15880
rect 15900 15640 16140 15880
rect 16230 15640 16470 15880
rect 16560 15640 16800 15880
rect 16890 15640 17130 15880
rect 17220 15640 17460 15880
rect 17550 15640 17790 15880
rect 17880 15640 18120 15880
rect 18210 15640 18450 15880
rect 18540 15640 18780 15880
rect 18870 15640 19110 15880
rect 19200 15640 19440 15880
rect 19530 15640 19770 15880
rect 19860 15640 20100 15880
rect 8310 15310 8550 15550
rect 8640 15310 8880 15550
rect 8970 15310 9210 15550
rect 9300 15310 9540 15550
rect 9630 15310 9870 15550
rect 9960 15310 10200 15550
rect 10290 15310 10530 15550
rect 10620 15310 10860 15550
rect 10950 15310 11190 15550
rect 11280 15310 11520 15550
rect 11610 15310 11850 15550
rect 11940 15310 12180 15550
rect 12270 15310 12510 15550
rect 12600 15310 12840 15550
rect 12930 15310 13170 15550
rect 13260 15310 13500 15550
rect 13590 15310 13830 15550
rect 13920 15310 14160 15550
rect 14250 15310 14490 15550
rect 14580 15310 14820 15550
rect 14910 15310 15150 15550
rect 15240 15310 15480 15550
rect 15570 15310 15810 15550
rect 15900 15310 16140 15550
rect 16230 15310 16470 15550
rect 16560 15310 16800 15550
rect 16890 15310 17130 15550
rect 17220 15310 17460 15550
rect 17550 15310 17790 15550
rect 17880 15310 18120 15550
rect 18210 15310 18450 15550
rect 18540 15310 18780 15550
rect 18870 15310 19110 15550
rect 19200 15310 19440 15550
rect 19530 15310 19770 15550
rect 19860 15310 20100 15550
rect 8310 14980 8550 15220
rect 8640 14980 8880 15220
rect 8970 14980 9210 15220
rect 9300 14980 9540 15220
rect 9630 14980 9870 15220
rect 9960 14980 10200 15220
rect 10290 14980 10530 15220
rect 10620 14980 10860 15220
rect 10950 14980 11190 15220
rect 11280 14980 11520 15220
rect 11610 14980 11850 15220
rect 11940 14980 12180 15220
rect 12270 14980 12510 15220
rect 12600 14980 12840 15220
rect 12930 14980 13170 15220
rect 13260 14980 13500 15220
rect 13590 14980 13830 15220
rect 13920 14980 14160 15220
rect 14250 14980 14490 15220
rect 14580 14980 14820 15220
rect 14910 14980 15150 15220
rect 15240 14980 15480 15220
rect 15570 14980 15810 15220
rect 15900 14980 16140 15220
rect 16230 14980 16470 15220
rect 16560 14980 16800 15220
rect 16890 14980 17130 15220
rect 17220 14980 17460 15220
rect 17550 14980 17790 15220
rect 17880 14980 18120 15220
rect 18210 14980 18450 15220
rect 18540 14980 18780 15220
rect 18870 14980 19110 15220
rect 19200 14980 19440 15220
rect 19530 14980 19770 15220
rect 19860 14980 20100 15220
rect 8310 14650 8550 14890
rect 8640 14650 8880 14890
rect 8970 14650 9210 14890
rect 9300 14650 9540 14890
rect 9630 14650 9870 14890
rect 9960 14650 10200 14890
rect 10290 14650 10530 14890
rect 10620 14650 10860 14890
rect 10950 14650 11190 14890
rect 11280 14650 11520 14890
rect 11610 14650 11850 14890
rect 11940 14650 12180 14890
rect 12270 14650 12510 14890
rect 12600 14650 12840 14890
rect 12930 14650 13170 14890
rect 13260 14650 13500 14890
rect 13590 14650 13830 14890
rect 13920 14650 14160 14890
rect 14250 14650 14490 14890
rect 14580 14650 14820 14890
rect 14910 14650 15150 14890
rect 15240 14650 15480 14890
rect 15570 14650 15810 14890
rect 15900 14650 16140 14890
rect 16230 14650 16470 14890
rect 16560 14650 16800 14890
rect 16890 14650 17130 14890
rect 17220 14650 17460 14890
rect 17550 14650 17790 14890
rect 17880 14650 18120 14890
rect 18210 14650 18450 14890
rect 18540 14650 18780 14890
rect 18870 14650 19110 14890
rect 19200 14650 19440 14890
rect 19530 14650 19770 14890
rect 19860 14650 20100 14890
rect 8310 14320 8550 14560
rect 8640 14320 8880 14560
rect 8970 14320 9210 14560
rect 9300 14320 9540 14560
rect 9630 14320 9870 14560
rect 9960 14320 10200 14560
rect 10290 14320 10530 14560
rect 10620 14320 10860 14560
rect 10950 14320 11190 14560
rect 11280 14320 11520 14560
rect 11610 14320 11850 14560
rect 11940 14320 12180 14560
rect 12270 14320 12510 14560
rect 12600 14320 12840 14560
rect 12930 14320 13170 14560
rect 13260 14320 13500 14560
rect 13590 14320 13830 14560
rect 13920 14320 14160 14560
rect 14250 14320 14490 14560
rect 14580 14320 14820 14560
rect 14910 14320 15150 14560
rect 15240 14320 15480 14560
rect 15570 14320 15810 14560
rect 15900 14320 16140 14560
rect 16230 14320 16470 14560
rect 16560 14320 16800 14560
rect 16890 14320 17130 14560
rect 17220 14320 17460 14560
rect 17550 14320 17790 14560
rect 17880 14320 18120 14560
rect 18210 14320 18450 14560
rect 18540 14320 18780 14560
rect 18870 14320 19110 14560
rect 19200 14320 19440 14560
rect 19530 14320 19770 14560
rect 19860 14320 20100 14560
rect 8310 13990 8550 14230
rect 8640 13990 8880 14230
rect 8970 13990 9210 14230
rect 9300 13990 9540 14230
rect 9630 13990 9870 14230
rect 9960 13990 10200 14230
rect 10290 13990 10530 14230
rect 10620 13990 10860 14230
rect 10950 13990 11190 14230
rect 11280 13990 11520 14230
rect 11610 13990 11850 14230
rect 11940 13990 12180 14230
rect 12270 13990 12510 14230
rect 12600 13990 12840 14230
rect 12930 13990 13170 14230
rect 13260 13990 13500 14230
rect 13590 13990 13830 14230
rect 13920 13990 14160 14230
rect 14250 13990 14490 14230
rect 14580 13990 14820 14230
rect 14910 13990 15150 14230
rect 15240 13990 15480 14230
rect 15570 13990 15810 14230
rect 15900 13990 16140 14230
rect 16230 13990 16470 14230
rect 16560 13990 16800 14230
rect 16890 13990 17130 14230
rect 17220 13990 17460 14230
rect 17550 13990 17790 14230
rect 17880 13990 18120 14230
rect 18210 13990 18450 14230
rect 18540 13990 18780 14230
rect 18870 13990 19110 14230
rect 19200 13990 19440 14230
rect 19530 13990 19770 14230
rect 19860 13990 20100 14230
rect 8310 13660 8550 13900
rect 8640 13660 8880 13900
rect 8970 13660 9210 13900
rect 9300 13660 9540 13900
rect 9630 13660 9870 13900
rect 9960 13660 10200 13900
rect 10290 13660 10530 13900
rect 10620 13660 10860 13900
rect 10950 13660 11190 13900
rect 11280 13660 11520 13900
rect 11610 13660 11850 13900
rect 11940 13660 12180 13900
rect 12270 13660 12510 13900
rect 12600 13660 12840 13900
rect 12930 13660 13170 13900
rect 13260 13660 13500 13900
rect 13590 13660 13830 13900
rect 13920 13660 14160 13900
rect 14250 13660 14490 13900
rect 14580 13660 14820 13900
rect 14910 13660 15150 13900
rect 15240 13660 15480 13900
rect 15570 13660 15810 13900
rect 15900 13660 16140 13900
rect 16230 13660 16470 13900
rect 16560 13660 16800 13900
rect 16890 13660 17130 13900
rect 17220 13660 17460 13900
rect 17550 13660 17790 13900
rect 17880 13660 18120 13900
rect 18210 13660 18450 13900
rect 18540 13660 18780 13900
rect 18870 13660 19110 13900
rect 19200 13660 19440 13900
rect 19530 13660 19770 13900
rect 19860 13660 20100 13900
rect 8310 13330 8550 13570
rect 8640 13330 8880 13570
rect 8970 13330 9210 13570
rect 9300 13330 9540 13570
rect 9630 13330 9870 13570
rect 9960 13330 10200 13570
rect 10290 13330 10530 13570
rect 10620 13330 10860 13570
rect 10950 13330 11190 13570
rect 11280 13330 11520 13570
rect 11610 13330 11850 13570
rect 11940 13330 12180 13570
rect 12270 13330 12510 13570
rect 12600 13330 12840 13570
rect 12930 13330 13170 13570
rect 13260 13330 13500 13570
rect 13590 13330 13830 13570
rect 13920 13330 14160 13570
rect 14250 13330 14490 13570
rect 14580 13330 14820 13570
rect 14910 13330 15150 13570
rect 15240 13330 15480 13570
rect 15570 13330 15810 13570
rect 15900 13330 16140 13570
rect 16230 13330 16470 13570
rect 16560 13330 16800 13570
rect 16890 13330 17130 13570
rect 17220 13330 17460 13570
rect 17550 13330 17790 13570
rect 17880 13330 18120 13570
rect 18210 13330 18450 13570
rect 18540 13330 18780 13570
rect 18870 13330 19110 13570
rect 19200 13330 19440 13570
rect 19530 13330 19770 13570
rect 19860 13330 20100 13570
rect 8310 13000 8550 13240
rect 8640 13000 8880 13240
rect 8970 13000 9210 13240
rect 9300 13000 9540 13240
rect 9630 13000 9870 13240
rect 9960 13000 10200 13240
rect 10290 13000 10530 13240
rect 10620 13000 10860 13240
rect 10950 13000 11190 13240
rect 11280 13000 11520 13240
rect 11610 13000 11850 13240
rect 11940 13000 12180 13240
rect 12270 13000 12510 13240
rect 12600 13000 12840 13240
rect 12930 13000 13170 13240
rect 13260 13000 13500 13240
rect 13590 13000 13830 13240
rect 13920 13000 14160 13240
rect 14250 13000 14490 13240
rect 14580 13000 14820 13240
rect 14910 13000 15150 13240
rect 15240 13000 15480 13240
rect 15570 13000 15810 13240
rect 15900 13000 16140 13240
rect 16230 13000 16470 13240
rect 16560 13000 16800 13240
rect 16890 13000 17130 13240
rect 17220 13000 17460 13240
rect 17550 13000 17790 13240
rect 17880 13000 18120 13240
rect 18210 13000 18450 13240
rect 18540 13000 18780 13240
rect 18870 13000 19110 13240
rect 19200 13000 19440 13240
rect 19530 13000 19770 13240
rect 19860 13000 20100 13240
rect 8310 12670 8550 12910
rect 8640 12670 8880 12910
rect 8970 12670 9210 12910
rect 9300 12670 9540 12910
rect 9630 12670 9870 12910
rect 9960 12670 10200 12910
rect 10290 12670 10530 12910
rect 10620 12670 10860 12910
rect 10950 12670 11190 12910
rect 11280 12670 11520 12910
rect 11610 12670 11850 12910
rect 11940 12670 12180 12910
rect 12270 12670 12510 12910
rect 12600 12670 12840 12910
rect 12930 12670 13170 12910
rect 13260 12670 13500 12910
rect 13590 12670 13830 12910
rect 13920 12670 14160 12910
rect 14250 12670 14490 12910
rect 14580 12670 14820 12910
rect 14910 12670 15150 12910
rect 15240 12670 15480 12910
rect 15570 12670 15810 12910
rect 15900 12670 16140 12910
rect 16230 12670 16470 12910
rect 16560 12670 16800 12910
rect 16890 12670 17130 12910
rect 17220 12670 17460 12910
rect 17550 12670 17790 12910
rect 17880 12670 18120 12910
rect 18210 12670 18450 12910
rect 18540 12670 18780 12910
rect 18870 12670 19110 12910
rect 19200 12670 19440 12910
rect 19530 12670 19770 12910
rect 19860 12670 20100 12910
rect 8310 12340 8550 12580
rect 8640 12340 8880 12580
rect 8970 12340 9210 12580
rect 9300 12340 9540 12580
rect 9630 12340 9870 12580
rect 9960 12340 10200 12580
rect 10290 12340 10530 12580
rect 10620 12340 10860 12580
rect 10950 12340 11190 12580
rect 11280 12340 11520 12580
rect 11610 12340 11850 12580
rect 11940 12340 12180 12580
rect 12270 12340 12510 12580
rect 12600 12340 12840 12580
rect 12930 12340 13170 12580
rect 13260 12340 13500 12580
rect 13590 12340 13830 12580
rect 13920 12340 14160 12580
rect 14250 12340 14490 12580
rect 14580 12340 14820 12580
rect 14910 12340 15150 12580
rect 15240 12340 15480 12580
rect 15570 12340 15810 12580
rect 15900 12340 16140 12580
rect 16230 12340 16470 12580
rect 16560 12340 16800 12580
rect 16890 12340 17130 12580
rect 17220 12340 17460 12580
rect 17550 12340 17790 12580
rect 17880 12340 18120 12580
rect 18210 12340 18450 12580
rect 18540 12340 18780 12580
rect 18870 12340 19110 12580
rect 19200 12340 19440 12580
rect 19530 12340 19770 12580
rect 19860 12340 20100 12580
rect 8310 12010 8550 12250
rect 8640 12010 8880 12250
rect 8970 12010 9210 12250
rect 9300 12010 9540 12250
rect 9630 12010 9870 12250
rect 9960 12010 10200 12250
rect 10290 12010 10530 12250
rect 10620 12010 10860 12250
rect 10950 12010 11190 12250
rect 11280 12010 11520 12250
rect 11610 12010 11850 12250
rect 11940 12010 12180 12250
rect 12270 12010 12510 12250
rect 12600 12010 12840 12250
rect 12930 12010 13170 12250
rect 13260 12010 13500 12250
rect 13590 12010 13830 12250
rect 13920 12010 14160 12250
rect 14250 12010 14490 12250
rect 14580 12010 14820 12250
rect 14910 12010 15150 12250
rect 15240 12010 15480 12250
rect 15570 12010 15810 12250
rect 15900 12010 16140 12250
rect 16230 12010 16470 12250
rect 16560 12010 16800 12250
rect 16890 12010 17130 12250
rect 17220 12010 17460 12250
rect 17550 12010 17790 12250
rect 17880 12010 18120 12250
rect 18210 12010 18450 12250
rect 18540 12010 18780 12250
rect 18870 12010 19110 12250
rect 19200 12010 19440 12250
rect 19530 12010 19770 12250
rect 19860 12010 20100 12250
rect 8310 11680 8550 11920
rect 8640 11680 8880 11920
rect 8970 11680 9210 11920
rect 9300 11680 9540 11920
rect 9630 11680 9870 11920
rect 9960 11680 10200 11920
rect 10290 11680 10530 11920
rect 10620 11680 10860 11920
rect 10950 11680 11190 11920
rect 11280 11680 11520 11920
rect 11610 11680 11850 11920
rect 11940 11680 12180 11920
rect 12270 11680 12510 11920
rect 12600 11680 12840 11920
rect 12930 11680 13170 11920
rect 13260 11680 13500 11920
rect 13590 11680 13830 11920
rect 13920 11680 14160 11920
rect 14250 11680 14490 11920
rect 14580 11680 14820 11920
rect 14910 11680 15150 11920
rect 15240 11680 15480 11920
rect 15570 11680 15810 11920
rect 15900 11680 16140 11920
rect 16230 11680 16470 11920
rect 16560 11680 16800 11920
rect 16890 11680 17130 11920
rect 17220 11680 17460 11920
rect 17550 11680 17790 11920
rect 17880 11680 18120 11920
rect 18210 11680 18450 11920
rect 18540 11680 18780 11920
rect 18870 11680 19110 11920
rect 19200 11680 19440 11920
rect 19530 11680 19770 11920
rect 19860 11680 20100 11920
rect 8310 11350 8550 11590
rect 8640 11350 8880 11590
rect 8970 11350 9210 11590
rect 9300 11350 9540 11590
rect 9630 11350 9870 11590
rect 9960 11350 10200 11590
rect 10290 11350 10530 11590
rect 10620 11350 10860 11590
rect 10950 11350 11190 11590
rect 11280 11350 11520 11590
rect 11610 11350 11850 11590
rect 11940 11350 12180 11590
rect 12270 11350 12510 11590
rect 12600 11350 12840 11590
rect 12930 11350 13170 11590
rect 13260 11350 13500 11590
rect 13590 11350 13830 11590
rect 13920 11350 14160 11590
rect 14250 11350 14490 11590
rect 14580 11350 14820 11590
rect 14910 11350 15150 11590
rect 15240 11350 15480 11590
rect 15570 11350 15810 11590
rect 15900 11350 16140 11590
rect 16230 11350 16470 11590
rect 16560 11350 16800 11590
rect 16890 11350 17130 11590
rect 17220 11350 17460 11590
rect 17550 11350 17790 11590
rect 17880 11350 18120 11590
rect 18210 11350 18450 11590
rect 18540 11350 18780 11590
rect 18870 11350 19110 11590
rect 19200 11350 19440 11590
rect 19530 11350 19770 11590
rect 19860 11350 20100 11590
rect 8310 11020 8550 11260
rect 8640 11020 8880 11260
rect 8970 11020 9210 11260
rect 9300 11020 9540 11260
rect 9630 11020 9870 11260
rect 9960 11020 10200 11260
rect 10290 11020 10530 11260
rect 10620 11020 10860 11260
rect 10950 11020 11190 11260
rect 11280 11020 11520 11260
rect 11610 11020 11850 11260
rect 11940 11020 12180 11260
rect 12270 11020 12510 11260
rect 12600 11020 12840 11260
rect 12930 11020 13170 11260
rect 13260 11020 13500 11260
rect 13590 11020 13830 11260
rect 13920 11020 14160 11260
rect 14250 11020 14490 11260
rect 14580 11020 14820 11260
rect 14910 11020 15150 11260
rect 15240 11020 15480 11260
rect 15570 11020 15810 11260
rect 15900 11020 16140 11260
rect 16230 11020 16470 11260
rect 16560 11020 16800 11260
rect 16890 11020 17130 11260
rect 17220 11020 17460 11260
rect 17550 11020 17790 11260
rect 17880 11020 18120 11260
rect 18210 11020 18450 11260
rect 18540 11020 18780 11260
rect 18870 11020 19110 11260
rect 19200 11020 19440 11260
rect 19530 11020 19770 11260
rect 19860 11020 20100 11260
rect 8310 10690 8550 10930
rect 8640 10690 8880 10930
rect 8970 10690 9210 10930
rect 9300 10690 9540 10930
rect 9630 10690 9870 10930
rect 9960 10690 10200 10930
rect 10290 10690 10530 10930
rect 10620 10690 10860 10930
rect 10950 10690 11190 10930
rect 11280 10690 11520 10930
rect 11610 10690 11850 10930
rect 11940 10690 12180 10930
rect 12270 10690 12510 10930
rect 12600 10690 12840 10930
rect 12930 10690 13170 10930
rect 13260 10690 13500 10930
rect 13590 10690 13830 10930
rect 13920 10690 14160 10930
rect 14250 10690 14490 10930
rect 14580 10690 14820 10930
rect 14910 10690 15150 10930
rect 15240 10690 15480 10930
rect 15570 10690 15810 10930
rect 15900 10690 16140 10930
rect 16230 10690 16470 10930
rect 16560 10690 16800 10930
rect 16890 10690 17130 10930
rect 17220 10690 17460 10930
rect 17550 10690 17790 10930
rect 17880 10690 18120 10930
rect 18210 10690 18450 10930
rect 18540 10690 18780 10930
rect 18870 10690 19110 10930
rect 19200 10690 19440 10930
rect 19530 10690 19770 10930
rect 19860 10690 20100 10930
rect 8310 10360 8550 10600
rect 8640 10360 8880 10600
rect 8970 10360 9210 10600
rect 9300 10360 9540 10600
rect 9630 10360 9870 10600
rect 9960 10360 10200 10600
rect 10290 10360 10530 10600
rect 10620 10360 10860 10600
rect 10950 10360 11190 10600
rect 11280 10360 11520 10600
rect 11610 10360 11850 10600
rect 11940 10360 12180 10600
rect 12270 10360 12510 10600
rect 12600 10360 12840 10600
rect 12930 10360 13170 10600
rect 13260 10360 13500 10600
rect 13590 10360 13830 10600
rect 13920 10360 14160 10600
rect 14250 10360 14490 10600
rect 14580 10360 14820 10600
rect 14910 10360 15150 10600
rect 15240 10360 15480 10600
rect 15570 10360 15810 10600
rect 15900 10360 16140 10600
rect 16230 10360 16470 10600
rect 16560 10360 16800 10600
rect 16890 10360 17130 10600
rect 17220 10360 17460 10600
rect 17550 10360 17790 10600
rect 17880 10360 18120 10600
rect 18210 10360 18450 10600
rect 18540 10360 18780 10600
rect 18870 10360 19110 10600
rect 19200 10360 19440 10600
rect 19530 10360 19770 10600
rect 19860 10360 20100 10600
rect 8310 10030 8550 10270
rect 8640 10030 8880 10270
rect 8970 10030 9210 10270
rect 9300 10030 9540 10270
rect 9630 10030 9870 10270
rect 9960 10030 10200 10270
rect 10290 10030 10530 10270
rect 10620 10030 10860 10270
rect 10950 10030 11190 10270
rect 11280 10030 11520 10270
rect 11610 10030 11850 10270
rect 11940 10030 12180 10270
rect 12270 10030 12510 10270
rect 12600 10030 12840 10270
rect 12930 10030 13170 10270
rect 13260 10030 13500 10270
rect 13590 10030 13830 10270
rect 13920 10030 14160 10270
rect 14250 10030 14490 10270
rect 14580 10030 14820 10270
rect 14910 10030 15150 10270
rect 15240 10030 15480 10270
rect 15570 10030 15810 10270
rect 15900 10030 16140 10270
rect 16230 10030 16470 10270
rect 16560 10030 16800 10270
rect 16890 10030 17130 10270
rect 17220 10030 17460 10270
rect 17550 10030 17790 10270
rect 17880 10030 18120 10270
rect 18210 10030 18450 10270
rect 18540 10030 18780 10270
rect 18870 10030 19110 10270
rect 19200 10030 19440 10270
rect 19530 10030 19770 10270
rect 19860 10030 20100 10270
rect 8310 9700 8550 9940
rect 8640 9700 8880 9940
rect 8970 9700 9210 9940
rect 9300 9700 9540 9940
rect 9630 9700 9870 9940
rect 9960 9700 10200 9940
rect 10290 9700 10530 9940
rect 10620 9700 10860 9940
rect 10950 9700 11190 9940
rect 11280 9700 11520 9940
rect 11610 9700 11850 9940
rect 11940 9700 12180 9940
rect 12270 9700 12510 9940
rect 12600 9700 12840 9940
rect 12930 9700 13170 9940
rect 13260 9700 13500 9940
rect 13590 9700 13830 9940
rect 13920 9700 14160 9940
rect 14250 9700 14490 9940
rect 14580 9700 14820 9940
rect 14910 9700 15150 9940
rect 15240 9700 15480 9940
rect 15570 9700 15810 9940
rect 15900 9700 16140 9940
rect 16230 9700 16470 9940
rect 16560 9700 16800 9940
rect 16890 9700 17130 9940
rect 17220 9700 17460 9940
rect 17550 9700 17790 9940
rect 17880 9700 18120 9940
rect 18210 9700 18450 9940
rect 18540 9700 18780 9940
rect 18870 9700 19110 9940
rect 19200 9700 19440 9940
rect 19530 9700 19770 9940
rect 19860 9700 20100 9940
rect 8310 9370 8550 9610
rect 8640 9370 8880 9610
rect 8970 9370 9210 9610
rect 9300 9370 9540 9610
rect 9630 9370 9870 9610
rect 9960 9370 10200 9610
rect 10290 9370 10530 9610
rect 10620 9370 10860 9610
rect 10950 9370 11190 9610
rect 11280 9370 11520 9610
rect 11610 9370 11850 9610
rect 11940 9370 12180 9610
rect 12270 9370 12510 9610
rect 12600 9370 12840 9610
rect 12930 9370 13170 9610
rect 13260 9370 13500 9610
rect 13590 9370 13830 9610
rect 13920 9370 14160 9610
rect 14250 9370 14490 9610
rect 14580 9370 14820 9610
rect 14910 9370 15150 9610
rect 15240 9370 15480 9610
rect 15570 9370 15810 9610
rect 15900 9370 16140 9610
rect 16230 9370 16470 9610
rect 16560 9370 16800 9610
rect 16890 9370 17130 9610
rect 17220 9370 17460 9610
rect 17550 9370 17790 9610
rect 17880 9370 18120 9610
rect 18210 9370 18450 9610
rect 18540 9370 18780 9610
rect 18870 9370 19110 9610
rect 19200 9370 19440 9610
rect 19530 9370 19770 9610
rect 19860 9370 20100 9610
rect 8310 9040 8550 9280
rect 8640 9040 8880 9280
rect 8970 9040 9210 9280
rect 9300 9040 9540 9280
rect 9630 9040 9870 9280
rect 9960 9040 10200 9280
rect 10290 9040 10530 9280
rect 10620 9040 10860 9280
rect 10950 9040 11190 9280
rect 11280 9040 11520 9280
rect 11610 9040 11850 9280
rect 11940 9040 12180 9280
rect 12270 9040 12510 9280
rect 12600 9040 12840 9280
rect 12930 9040 13170 9280
rect 13260 9040 13500 9280
rect 13590 9040 13830 9280
rect 13920 9040 14160 9280
rect 14250 9040 14490 9280
rect 14580 9040 14820 9280
rect 14910 9040 15150 9280
rect 15240 9040 15480 9280
rect 15570 9040 15810 9280
rect 15900 9040 16140 9280
rect 16230 9040 16470 9280
rect 16560 9040 16800 9280
rect 16890 9040 17130 9280
rect 17220 9040 17460 9280
rect 17550 9040 17790 9280
rect 17880 9040 18120 9280
rect 18210 9040 18450 9280
rect 18540 9040 18780 9280
rect 18870 9040 19110 9280
rect 19200 9040 19440 9280
rect 19530 9040 19770 9280
rect 19860 9040 20100 9280
rect 31180 7590 31420 7830
rect 31510 7590 31750 7830
rect 31840 7590 32080 7830
rect 32170 7590 32410 7830
rect 32500 7590 32740 7830
rect 32830 7590 33070 7830
rect 33160 7590 33400 7830
rect 33490 7590 33730 7830
rect 33820 7590 34060 7830
rect 34150 7590 34390 7830
rect 34480 7590 34720 7830
rect 34810 7590 35050 7830
rect 35140 7590 35380 7830
rect 35470 7590 35710 7830
rect 35800 7590 36040 7830
rect 36130 7590 36370 7830
rect 36460 7590 36700 7830
rect 36790 7590 37030 7830
rect 37120 7590 37360 7830
rect 37450 7590 37690 7830
rect 31180 7260 31420 7500
rect 31510 7260 31750 7500
rect 31840 7260 32080 7500
rect 32170 7260 32410 7500
rect 32500 7260 32740 7500
rect 32830 7260 33070 7500
rect 33160 7260 33400 7500
rect 33490 7260 33730 7500
rect 33820 7260 34060 7500
rect 34150 7260 34390 7500
rect 34480 7260 34720 7500
rect 34810 7260 35050 7500
rect 35140 7260 35380 7500
rect 35470 7260 35710 7500
rect 35800 7260 36040 7500
rect 36130 7260 36370 7500
rect 36460 7260 36700 7500
rect 36790 7260 37030 7500
rect 37120 7260 37360 7500
rect 37450 7260 37690 7500
rect 31180 6930 31420 7170
rect 31510 6930 31750 7170
rect 31840 6930 32080 7170
rect 32170 6930 32410 7170
rect 32500 6930 32740 7170
rect 32830 6930 33070 7170
rect 33160 6930 33400 7170
rect 33490 6930 33730 7170
rect 33820 6930 34060 7170
rect 34150 6930 34390 7170
rect 34480 6930 34720 7170
rect 34810 6930 35050 7170
rect 35140 6930 35380 7170
rect 35470 6930 35710 7170
rect 35800 6930 36040 7170
rect 36130 6930 36370 7170
rect 36460 6930 36700 7170
rect 36790 6930 37030 7170
rect 37120 6930 37360 7170
rect 37450 6930 37690 7170
rect 31180 6600 31420 6840
rect 31510 6600 31750 6840
rect 31840 6600 32080 6840
rect 32170 6600 32410 6840
rect 32500 6600 32740 6840
rect 32830 6600 33070 6840
rect 33160 6600 33400 6840
rect 33490 6600 33730 6840
rect 33820 6600 34060 6840
rect 34150 6600 34390 6840
rect 34480 6600 34720 6840
rect 34810 6600 35050 6840
rect 35140 6600 35380 6840
rect 35470 6600 35710 6840
rect 35800 6600 36040 6840
rect 36130 6600 36370 6840
rect 36460 6600 36700 6840
rect 36790 6600 37030 6840
rect 37120 6600 37360 6840
rect 37450 6600 37690 6840
rect 31180 6270 31420 6510
rect 31510 6270 31750 6510
rect 31840 6270 32080 6510
rect 32170 6270 32410 6510
rect 32500 6270 32740 6510
rect 32830 6270 33070 6510
rect 33160 6270 33400 6510
rect 33490 6270 33730 6510
rect 33820 6270 34060 6510
rect 34150 6270 34390 6510
rect 34480 6270 34720 6510
rect 34810 6270 35050 6510
rect 35140 6270 35380 6510
rect 35470 6270 35710 6510
rect 35800 6270 36040 6510
rect 36130 6270 36370 6510
rect 36460 6270 36700 6510
rect 36790 6270 37030 6510
rect 37120 6270 37360 6510
rect 37450 6270 37690 6510
rect 31180 5940 31420 6180
rect 31510 5940 31750 6180
rect 31840 5940 32080 6180
rect 32170 5940 32410 6180
rect 32500 5940 32740 6180
rect 32830 5940 33070 6180
rect 33160 5940 33400 6180
rect 33490 5940 33730 6180
rect 33820 5940 34060 6180
rect 34150 5940 34390 6180
rect 34480 5940 34720 6180
rect 34810 5940 35050 6180
rect 35140 5940 35380 6180
rect 35470 5940 35710 6180
rect 35800 5940 36040 6180
rect 36130 5940 36370 6180
rect 36460 5940 36700 6180
rect 36790 5940 37030 6180
rect 37120 5940 37360 6180
rect 37450 5940 37690 6180
rect 31180 5610 31420 5850
rect 31510 5610 31750 5850
rect 31840 5610 32080 5850
rect 32170 5610 32410 5850
rect 32500 5610 32740 5850
rect 32830 5610 33070 5850
rect 33160 5610 33400 5850
rect 33490 5610 33730 5850
rect 33820 5610 34060 5850
rect 34150 5610 34390 5850
rect 34480 5610 34720 5850
rect 34810 5610 35050 5850
rect 35140 5610 35380 5850
rect 35470 5610 35710 5850
rect 35800 5610 36040 5850
rect 36130 5610 36370 5850
rect 36460 5610 36700 5850
rect 36790 5610 37030 5850
rect 37120 5610 37360 5850
rect 37450 5610 37690 5850
rect 31180 5280 31420 5520
rect 31510 5280 31750 5520
rect 31840 5280 32080 5520
rect 32170 5280 32410 5520
rect 32500 5280 32740 5520
rect 32830 5280 33070 5520
rect 33160 5280 33400 5520
rect 33490 5280 33730 5520
rect 33820 5280 34060 5520
rect 34150 5280 34390 5520
rect 34480 5280 34720 5520
rect 34810 5280 35050 5520
rect 35140 5280 35380 5520
rect 35470 5280 35710 5520
rect 35800 5280 36040 5520
rect 36130 5280 36370 5520
rect 36460 5280 36700 5520
rect 36790 5280 37030 5520
rect 37120 5280 37360 5520
rect 37450 5280 37690 5520
rect 31180 4950 31420 5190
rect 31510 4950 31750 5190
rect 31840 4950 32080 5190
rect 32170 4950 32410 5190
rect 32500 4950 32740 5190
rect 32830 4950 33070 5190
rect 33160 4950 33400 5190
rect 33490 4950 33730 5190
rect 33820 4950 34060 5190
rect 34150 4950 34390 5190
rect 34480 4950 34720 5190
rect 34810 4950 35050 5190
rect 35140 4950 35380 5190
rect 35470 4950 35710 5190
rect 35800 4950 36040 5190
rect 36130 4950 36370 5190
rect 36460 4950 36700 5190
rect 36790 4950 37030 5190
rect 37120 4950 37360 5190
rect 37450 4950 37690 5190
rect 31180 4620 31420 4860
rect 31510 4620 31750 4860
rect 31840 4620 32080 4860
rect 32170 4620 32410 4860
rect 32500 4620 32740 4860
rect 32830 4620 33070 4860
rect 33160 4620 33400 4860
rect 33490 4620 33730 4860
rect 33820 4620 34060 4860
rect 34150 4620 34390 4860
rect 34480 4620 34720 4860
rect 34810 4620 35050 4860
rect 35140 4620 35380 4860
rect 35470 4620 35710 4860
rect 35800 4620 36040 4860
rect 36130 4620 36370 4860
rect 36460 4620 36700 4860
rect 36790 4620 37030 4860
rect 37120 4620 37360 4860
rect 37450 4620 37690 4860
rect 31180 4290 31420 4530
rect 31510 4290 31750 4530
rect 31840 4290 32080 4530
rect 32170 4290 32410 4530
rect 32500 4290 32740 4530
rect 32830 4290 33070 4530
rect 33160 4290 33400 4530
rect 33490 4290 33730 4530
rect 33820 4290 34060 4530
rect 34150 4290 34390 4530
rect 34480 4290 34720 4530
rect 34810 4290 35050 4530
rect 35140 4290 35380 4530
rect 35470 4290 35710 4530
rect 35800 4290 36040 4530
rect 36130 4290 36370 4530
rect 36460 4290 36700 4530
rect 36790 4290 37030 4530
rect 37120 4290 37360 4530
rect 37450 4290 37690 4530
rect 31180 3960 31420 4200
rect 31510 3960 31750 4200
rect 31840 3960 32080 4200
rect 32170 3960 32410 4200
rect 32500 3960 32740 4200
rect 32830 3960 33070 4200
rect 33160 3960 33400 4200
rect 33490 3960 33730 4200
rect 33820 3960 34060 4200
rect 34150 3960 34390 4200
rect 34480 3960 34720 4200
rect 34810 3960 35050 4200
rect 35140 3960 35380 4200
rect 35470 3960 35710 4200
rect 35800 3960 36040 4200
rect 36130 3960 36370 4200
rect 36460 3960 36700 4200
rect 36790 3960 37030 4200
rect 37120 3960 37360 4200
rect 37450 3960 37690 4200
rect 31180 3630 31420 3870
rect 31510 3630 31750 3870
rect 31840 3630 32080 3870
rect 32170 3630 32410 3870
rect 32500 3630 32740 3870
rect 32830 3630 33070 3870
rect 33160 3630 33400 3870
rect 33490 3630 33730 3870
rect 33820 3630 34060 3870
rect 34150 3630 34390 3870
rect 34480 3630 34720 3870
rect 34810 3630 35050 3870
rect 35140 3630 35380 3870
rect 35470 3630 35710 3870
rect 35800 3630 36040 3870
rect 36130 3630 36370 3870
rect 36460 3630 36700 3870
rect 36790 3630 37030 3870
rect 37120 3630 37360 3870
rect 37450 3630 37690 3870
rect 31180 3300 31420 3540
rect 31510 3300 31750 3540
rect 31840 3300 32080 3540
rect 32170 3300 32410 3540
rect 32500 3300 32740 3540
rect 32830 3300 33070 3540
rect 33160 3300 33400 3540
rect 33490 3300 33730 3540
rect 33820 3300 34060 3540
rect 34150 3300 34390 3540
rect 34480 3300 34720 3540
rect 34810 3300 35050 3540
rect 35140 3300 35380 3540
rect 35470 3300 35710 3540
rect 35800 3300 36040 3540
rect 36130 3300 36370 3540
rect 36460 3300 36700 3540
rect 36790 3300 37030 3540
rect 37120 3300 37360 3540
rect 37450 3300 37690 3540
rect 31180 2970 31420 3210
rect 31510 2970 31750 3210
rect 31840 2970 32080 3210
rect 32170 2970 32410 3210
rect 32500 2970 32740 3210
rect 32830 2970 33070 3210
rect 33160 2970 33400 3210
rect 33490 2970 33730 3210
rect 33820 2970 34060 3210
rect 34150 2970 34390 3210
rect 34480 2970 34720 3210
rect 34810 2970 35050 3210
rect 35140 2970 35380 3210
rect 35470 2970 35710 3210
rect 35800 2970 36040 3210
rect 36130 2970 36370 3210
rect 36460 2970 36700 3210
rect 36790 2970 37030 3210
rect 37120 2970 37360 3210
rect 37450 2970 37690 3210
rect 31180 2640 31420 2880
rect 31510 2640 31750 2880
rect 31840 2640 32080 2880
rect 32170 2640 32410 2880
rect 32500 2640 32740 2880
rect 32830 2640 33070 2880
rect 33160 2640 33400 2880
rect 33490 2640 33730 2880
rect 33820 2640 34060 2880
rect 34150 2640 34390 2880
rect 34480 2640 34720 2880
rect 34810 2640 35050 2880
rect 35140 2640 35380 2880
rect 35470 2640 35710 2880
rect 35800 2640 36040 2880
rect 36130 2640 36370 2880
rect 36460 2640 36700 2880
rect 36790 2640 37030 2880
rect 37120 2640 37360 2880
rect 37450 2640 37690 2880
rect 31180 2310 31420 2550
rect 31510 2310 31750 2550
rect 31840 2310 32080 2550
rect 32170 2310 32410 2550
rect 32500 2310 32740 2550
rect 32830 2310 33070 2550
rect 33160 2310 33400 2550
rect 33490 2310 33730 2550
rect 33820 2310 34060 2550
rect 34150 2310 34390 2550
rect 34480 2310 34720 2550
rect 34810 2310 35050 2550
rect 35140 2310 35380 2550
rect 35470 2310 35710 2550
rect 35800 2310 36040 2550
rect 36130 2310 36370 2550
rect 36460 2310 36700 2550
rect 36790 2310 37030 2550
rect 37120 2310 37360 2550
rect 37450 2310 37690 2550
rect 31180 1980 31420 2220
rect 31510 1980 31750 2220
rect 31840 1980 32080 2220
rect 32170 1980 32410 2220
rect 32500 1980 32740 2220
rect 32830 1980 33070 2220
rect 33160 1980 33400 2220
rect 33490 1980 33730 2220
rect 33820 1980 34060 2220
rect 34150 1980 34390 2220
rect 34480 1980 34720 2220
rect 34810 1980 35050 2220
rect 35140 1980 35380 2220
rect 35470 1980 35710 2220
rect 35800 1980 36040 2220
rect 36130 1980 36370 2220
rect 36460 1980 36700 2220
rect 36790 1980 37030 2220
rect 37120 1980 37360 2220
rect 37450 1980 37690 2220
rect 31180 1650 31420 1890
rect 31510 1650 31750 1890
rect 31840 1650 32080 1890
rect 32170 1650 32410 1890
rect 32500 1650 32740 1890
rect 32830 1650 33070 1890
rect 33160 1650 33400 1890
rect 33490 1650 33730 1890
rect 33820 1650 34060 1890
rect 34150 1650 34390 1890
rect 34480 1650 34720 1890
rect 34810 1650 35050 1890
rect 35140 1650 35380 1890
rect 35470 1650 35710 1890
rect 35800 1650 36040 1890
rect 36130 1650 36370 1890
rect 36460 1650 36700 1890
rect 36790 1650 37030 1890
rect 37120 1650 37360 1890
rect 37450 1650 37690 1890
rect 31180 1320 31420 1560
rect 31510 1320 31750 1560
rect 31840 1320 32080 1560
rect 32170 1320 32410 1560
rect 32500 1320 32740 1560
rect 32830 1320 33070 1560
rect 33160 1320 33400 1560
rect 33490 1320 33730 1560
rect 33820 1320 34060 1560
rect 34150 1320 34390 1560
rect 34480 1320 34720 1560
rect 34810 1320 35050 1560
rect 35140 1320 35380 1560
rect 35470 1320 35710 1560
rect 35800 1320 36040 1560
rect 36130 1320 36370 1560
rect 36460 1320 36700 1560
rect 36790 1320 37030 1560
rect 37120 1320 37360 1560
rect 37450 1320 37690 1560
rect 31180 -10 31420 230
rect 31510 -10 31750 230
rect 31840 -10 32080 230
rect 32170 -10 32410 230
rect 32500 -10 32740 230
rect 32830 -10 33070 230
rect 33160 -10 33400 230
rect 33490 -10 33730 230
rect 33820 -10 34060 230
rect 34150 -10 34390 230
rect 34480 -10 34720 230
rect 34810 -10 35050 230
rect 35140 -10 35380 230
rect 35470 -10 35710 230
rect 35800 -10 36040 230
rect 36130 -10 36370 230
rect 36460 -10 36700 230
rect 36790 -10 37030 230
rect 37120 -10 37360 230
rect 37450 -10 37690 230
rect 31180 -340 31420 -100
rect 31510 -340 31750 -100
rect 31840 -340 32080 -100
rect 32170 -340 32410 -100
rect 32500 -340 32740 -100
rect 32830 -340 33070 -100
rect 33160 -340 33400 -100
rect 33490 -340 33730 -100
rect 33820 -340 34060 -100
rect 34150 -340 34390 -100
rect 34480 -340 34720 -100
rect 34810 -340 35050 -100
rect 35140 -340 35380 -100
rect 35470 -340 35710 -100
rect 35800 -340 36040 -100
rect 36130 -340 36370 -100
rect 36460 -340 36700 -100
rect 36790 -340 37030 -100
rect 37120 -340 37360 -100
rect 37450 -340 37690 -100
rect 31180 -670 31420 -430
rect 31510 -670 31750 -430
rect 31840 -670 32080 -430
rect 32170 -670 32410 -430
rect 32500 -670 32740 -430
rect 32830 -670 33070 -430
rect 33160 -670 33400 -430
rect 33490 -670 33730 -430
rect 33820 -670 34060 -430
rect 34150 -670 34390 -430
rect 34480 -670 34720 -430
rect 34810 -670 35050 -430
rect 35140 -670 35380 -430
rect 35470 -670 35710 -430
rect 35800 -670 36040 -430
rect 36130 -670 36370 -430
rect 36460 -670 36700 -430
rect 36790 -670 37030 -430
rect 37120 -670 37360 -430
rect 37450 -670 37690 -430
rect 31180 -1000 31420 -760
rect 31510 -1000 31750 -760
rect 31840 -1000 32080 -760
rect 32170 -1000 32410 -760
rect 32500 -1000 32740 -760
rect 32830 -1000 33070 -760
rect 33160 -1000 33400 -760
rect 33490 -1000 33730 -760
rect 33820 -1000 34060 -760
rect 34150 -1000 34390 -760
rect 34480 -1000 34720 -760
rect 34810 -1000 35050 -760
rect 35140 -1000 35380 -760
rect 35470 -1000 35710 -760
rect 35800 -1000 36040 -760
rect 36130 -1000 36370 -760
rect 36460 -1000 36700 -760
rect 36790 -1000 37030 -760
rect 37120 -1000 37360 -760
rect 37450 -1000 37690 -760
rect 31180 -1330 31420 -1090
rect 31510 -1330 31750 -1090
rect 31840 -1330 32080 -1090
rect 32170 -1330 32410 -1090
rect 32500 -1330 32740 -1090
rect 32830 -1330 33070 -1090
rect 33160 -1330 33400 -1090
rect 33490 -1330 33730 -1090
rect 33820 -1330 34060 -1090
rect 34150 -1330 34390 -1090
rect 34480 -1330 34720 -1090
rect 34810 -1330 35050 -1090
rect 35140 -1330 35380 -1090
rect 35470 -1330 35710 -1090
rect 35800 -1330 36040 -1090
rect 36130 -1330 36370 -1090
rect 36460 -1330 36700 -1090
rect 36790 -1330 37030 -1090
rect 37120 -1330 37360 -1090
rect 37450 -1330 37690 -1090
rect 31180 -1660 31420 -1420
rect 31510 -1660 31750 -1420
rect 31840 -1660 32080 -1420
rect 32170 -1660 32410 -1420
rect 32500 -1660 32740 -1420
rect 32830 -1660 33070 -1420
rect 33160 -1660 33400 -1420
rect 33490 -1660 33730 -1420
rect 33820 -1660 34060 -1420
rect 34150 -1660 34390 -1420
rect 34480 -1660 34720 -1420
rect 34810 -1660 35050 -1420
rect 35140 -1660 35380 -1420
rect 35470 -1660 35710 -1420
rect 35800 -1660 36040 -1420
rect 36130 -1660 36370 -1420
rect 36460 -1660 36700 -1420
rect 36790 -1660 37030 -1420
rect 37120 -1660 37360 -1420
rect 37450 -1660 37690 -1420
rect 31180 -1990 31420 -1750
rect 31510 -1990 31750 -1750
rect 31840 -1990 32080 -1750
rect 32170 -1990 32410 -1750
rect 32500 -1990 32740 -1750
rect 32830 -1990 33070 -1750
rect 33160 -1990 33400 -1750
rect 33490 -1990 33730 -1750
rect 33820 -1990 34060 -1750
rect 34150 -1990 34390 -1750
rect 34480 -1990 34720 -1750
rect 34810 -1990 35050 -1750
rect 35140 -1990 35380 -1750
rect 35470 -1990 35710 -1750
rect 35800 -1990 36040 -1750
rect 36130 -1990 36370 -1750
rect 36460 -1990 36700 -1750
rect 36790 -1990 37030 -1750
rect 37120 -1990 37360 -1750
rect 37450 -1990 37690 -1750
rect 31180 -2320 31420 -2080
rect 31510 -2320 31750 -2080
rect 31840 -2320 32080 -2080
rect 32170 -2320 32410 -2080
rect 32500 -2320 32740 -2080
rect 32830 -2320 33070 -2080
rect 33160 -2320 33400 -2080
rect 33490 -2320 33730 -2080
rect 33820 -2320 34060 -2080
rect 34150 -2320 34390 -2080
rect 34480 -2320 34720 -2080
rect 34810 -2320 35050 -2080
rect 35140 -2320 35380 -2080
rect 35470 -2320 35710 -2080
rect 35800 -2320 36040 -2080
rect 36130 -2320 36370 -2080
rect 36460 -2320 36700 -2080
rect 36790 -2320 37030 -2080
rect 37120 -2320 37360 -2080
rect 37450 -2320 37690 -2080
rect 31180 -2650 31420 -2410
rect 31510 -2650 31750 -2410
rect 31840 -2650 32080 -2410
rect 32170 -2650 32410 -2410
rect 32500 -2650 32740 -2410
rect 32830 -2650 33070 -2410
rect 33160 -2650 33400 -2410
rect 33490 -2650 33730 -2410
rect 33820 -2650 34060 -2410
rect 34150 -2650 34390 -2410
rect 34480 -2650 34720 -2410
rect 34810 -2650 35050 -2410
rect 35140 -2650 35380 -2410
rect 35470 -2650 35710 -2410
rect 35800 -2650 36040 -2410
rect 36130 -2650 36370 -2410
rect 36460 -2650 36700 -2410
rect 36790 -2650 37030 -2410
rect 37120 -2650 37360 -2410
rect 37450 -2650 37690 -2410
rect 31180 -2980 31420 -2740
rect 31510 -2980 31750 -2740
rect 31840 -2980 32080 -2740
rect 32170 -2980 32410 -2740
rect 32500 -2980 32740 -2740
rect 32830 -2980 33070 -2740
rect 33160 -2980 33400 -2740
rect 33490 -2980 33730 -2740
rect 33820 -2980 34060 -2740
rect 34150 -2980 34390 -2740
rect 34480 -2980 34720 -2740
rect 34810 -2980 35050 -2740
rect 35140 -2980 35380 -2740
rect 35470 -2980 35710 -2740
rect 35800 -2980 36040 -2740
rect 36130 -2980 36370 -2740
rect 36460 -2980 36700 -2740
rect 36790 -2980 37030 -2740
rect 37120 -2980 37360 -2740
rect 37450 -2980 37690 -2740
rect 31180 -3310 31420 -3070
rect 31510 -3310 31750 -3070
rect 31840 -3310 32080 -3070
rect 32170 -3310 32410 -3070
rect 32500 -3310 32740 -3070
rect 32830 -3310 33070 -3070
rect 33160 -3310 33400 -3070
rect 33490 -3310 33730 -3070
rect 33820 -3310 34060 -3070
rect 34150 -3310 34390 -3070
rect 34480 -3310 34720 -3070
rect 34810 -3310 35050 -3070
rect 35140 -3310 35380 -3070
rect 35470 -3310 35710 -3070
rect 35800 -3310 36040 -3070
rect 36130 -3310 36370 -3070
rect 36460 -3310 36700 -3070
rect 36790 -3310 37030 -3070
rect 37120 -3310 37360 -3070
rect 37450 -3310 37690 -3070
rect 31180 -3640 31420 -3400
rect 31510 -3640 31750 -3400
rect 31840 -3640 32080 -3400
rect 32170 -3640 32410 -3400
rect 32500 -3640 32740 -3400
rect 32830 -3640 33070 -3400
rect 33160 -3640 33400 -3400
rect 33490 -3640 33730 -3400
rect 33820 -3640 34060 -3400
rect 34150 -3640 34390 -3400
rect 34480 -3640 34720 -3400
rect 34810 -3640 35050 -3400
rect 35140 -3640 35380 -3400
rect 35470 -3640 35710 -3400
rect 35800 -3640 36040 -3400
rect 36130 -3640 36370 -3400
rect 36460 -3640 36700 -3400
rect 36790 -3640 37030 -3400
rect 37120 -3640 37360 -3400
rect 37450 -3640 37690 -3400
rect 31180 -3970 31420 -3730
rect 31510 -3970 31750 -3730
rect 31840 -3970 32080 -3730
rect 32170 -3970 32410 -3730
rect 32500 -3970 32740 -3730
rect 32830 -3970 33070 -3730
rect 33160 -3970 33400 -3730
rect 33490 -3970 33730 -3730
rect 33820 -3970 34060 -3730
rect 34150 -3970 34390 -3730
rect 34480 -3970 34720 -3730
rect 34810 -3970 35050 -3730
rect 35140 -3970 35380 -3730
rect 35470 -3970 35710 -3730
rect 35800 -3970 36040 -3730
rect 36130 -3970 36370 -3730
rect 36460 -3970 36700 -3730
rect 36790 -3970 37030 -3730
rect 37120 -3970 37360 -3730
rect 37450 -3970 37690 -3730
rect 31180 -4300 31420 -4060
rect 31510 -4300 31750 -4060
rect 31840 -4300 32080 -4060
rect 32170 -4300 32410 -4060
rect 32500 -4300 32740 -4060
rect 32830 -4300 33070 -4060
rect 33160 -4300 33400 -4060
rect 33490 -4300 33730 -4060
rect 33820 -4300 34060 -4060
rect 34150 -4300 34390 -4060
rect 34480 -4300 34720 -4060
rect 34810 -4300 35050 -4060
rect 35140 -4300 35380 -4060
rect 35470 -4300 35710 -4060
rect 35800 -4300 36040 -4060
rect 36130 -4300 36370 -4060
rect 36460 -4300 36700 -4060
rect 36790 -4300 37030 -4060
rect 37120 -4300 37360 -4060
rect 37450 -4300 37690 -4060
rect 31180 -4630 31420 -4390
rect 31510 -4630 31750 -4390
rect 31840 -4630 32080 -4390
rect 32170 -4630 32410 -4390
rect 32500 -4630 32740 -4390
rect 32830 -4630 33070 -4390
rect 33160 -4630 33400 -4390
rect 33490 -4630 33730 -4390
rect 33820 -4630 34060 -4390
rect 34150 -4630 34390 -4390
rect 34480 -4630 34720 -4390
rect 34810 -4630 35050 -4390
rect 35140 -4630 35380 -4390
rect 35470 -4630 35710 -4390
rect 35800 -4630 36040 -4390
rect 36130 -4630 36370 -4390
rect 36460 -4630 36700 -4390
rect 36790 -4630 37030 -4390
rect 37120 -4630 37360 -4390
rect 37450 -4630 37690 -4390
rect -1180 -5080 -940 -4840
rect -850 -5080 -610 -4840
rect -520 -5080 -280 -4840
rect -190 -5080 50 -4840
rect -1180 -5410 -940 -5170
rect -850 -5410 -610 -5170
rect -520 -5410 -280 -5170
rect -190 -5410 50 -5170
rect -1180 -5740 -940 -5500
rect -850 -5740 -610 -5500
rect -520 -5740 -280 -5500
rect -190 -5740 50 -5500
rect -1180 -6070 -940 -5830
rect -850 -6070 -610 -5830
rect -520 -6070 -280 -5830
rect -190 -6070 50 -5830
rect 14730 -5080 14970 -4840
rect 15060 -5080 15300 -4840
rect 15390 -5080 15630 -4840
rect 15720 -5080 15960 -4840
rect 14730 -5410 14970 -5170
rect 15060 -5410 15300 -5170
rect 15390 -5410 15630 -5170
rect 15720 -5410 15960 -5170
rect 14730 -5740 14970 -5500
rect 15060 -5740 15300 -5500
rect 15390 -5740 15630 -5500
rect 15720 -5740 15960 -5500
rect 14730 -6070 14970 -5830
rect 15060 -6070 15300 -5830
rect 15390 -6070 15630 -5830
rect 15720 -6070 15960 -5830
rect 31180 -4960 31420 -4720
rect 31510 -4960 31750 -4720
rect 31840 -4960 32080 -4720
rect 32170 -4960 32410 -4720
rect 32500 -4960 32740 -4720
rect 32830 -4960 33070 -4720
rect 33160 -4960 33400 -4720
rect 33490 -4960 33730 -4720
rect 33820 -4960 34060 -4720
rect 34150 -4960 34390 -4720
rect 34480 -4960 34720 -4720
rect 34810 -4960 35050 -4720
rect 35140 -4960 35380 -4720
rect 35470 -4960 35710 -4720
rect 35800 -4960 36040 -4720
rect 36130 -4960 36370 -4720
rect 36460 -4960 36700 -4720
rect 36790 -4960 37030 -4720
rect 37120 -4960 37360 -4720
rect 37450 -4960 37690 -4720
rect 31180 -5290 31420 -5050
rect 31510 -5290 31750 -5050
rect 31840 -5290 32080 -5050
rect 32170 -5290 32410 -5050
rect 32500 -5290 32740 -5050
rect 32830 -5290 33070 -5050
rect 33160 -5290 33400 -5050
rect 33490 -5290 33730 -5050
rect 33820 -5290 34060 -5050
rect 34150 -5290 34390 -5050
rect 34480 -5290 34720 -5050
rect 34810 -5290 35050 -5050
rect 35140 -5290 35380 -5050
rect 35470 -5290 35710 -5050
rect 35800 -5290 36040 -5050
rect 36130 -5290 36370 -5050
rect 36460 -5290 36700 -5050
rect 36790 -5290 37030 -5050
rect 37120 -5290 37360 -5050
rect 37450 -5290 37690 -5050
rect 31180 -5620 31420 -5380
rect 31510 -5620 31750 -5380
rect 31840 -5620 32080 -5380
rect 32170 -5620 32410 -5380
rect 32500 -5620 32740 -5380
rect 32830 -5620 33070 -5380
rect 33160 -5620 33400 -5380
rect 33490 -5620 33730 -5380
rect 33820 -5620 34060 -5380
rect 34150 -5620 34390 -5380
rect 34480 -5620 34720 -5380
rect 34810 -5620 35050 -5380
rect 35140 -5620 35380 -5380
rect 35470 -5620 35710 -5380
rect 35800 -5620 36040 -5380
rect 36130 -5620 36370 -5380
rect 36460 -5620 36700 -5380
rect 36790 -5620 37030 -5380
rect 37120 -5620 37360 -5380
rect 37450 -5620 37690 -5380
rect 31180 -5950 31420 -5710
rect 31510 -5950 31750 -5710
rect 31840 -5950 32080 -5710
rect 32170 -5950 32410 -5710
rect 32500 -5950 32740 -5710
rect 32830 -5950 33070 -5710
rect 33160 -5950 33400 -5710
rect 33490 -5950 33730 -5710
rect 33820 -5950 34060 -5710
rect 34150 -5950 34390 -5710
rect 34480 -5950 34720 -5710
rect 34810 -5950 35050 -5710
rect 35140 -5950 35380 -5710
rect 35470 -5950 35710 -5710
rect 35800 -5950 36040 -5710
rect 36130 -5950 36370 -5710
rect 36460 -5950 36700 -5710
rect 36790 -5950 37030 -5710
rect 37120 -5950 37360 -5710
rect 37450 -5950 37690 -5710
rect 31180 -6280 31420 -6040
rect 31510 -6280 31750 -6040
rect 31840 -6280 32080 -6040
rect 32170 -6280 32410 -6040
rect 32500 -6280 32740 -6040
rect 32830 -6280 33070 -6040
rect 33160 -6280 33400 -6040
rect 33490 -6280 33730 -6040
rect 33820 -6280 34060 -6040
rect 34150 -6280 34390 -6040
rect 34480 -6280 34720 -6040
rect 34810 -6280 35050 -6040
rect 35140 -6280 35380 -6040
rect 35470 -6280 35710 -6040
rect 35800 -6280 36040 -6040
rect 36130 -6280 36370 -6040
rect 36460 -6280 36700 -6040
rect 36790 -6280 37030 -6040
rect 37120 -6280 37360 -6040
rect 37450 -6280 37690 -6040
<< metal5 >>
rect -5550 21610 6760 21640
rect -5550 21370 -5180 21610
rect -4940 21370 -4850 21610
rect -4610 21370 -4520 21610
rect -4280 21370 -4190 21610
rect -3950 21370 -3860 21610
rect -3620 21370 -3530 21610
rect -3290 21370 -3200 21610
rect -2960 21370 -2870 21610
rect -2630 21370 -2540 21610
rect -2300 21370 -2170 21610
rect -1930 21370 -1840 21610
rect -1600 21370 -1510 21610
rect -1270 21370 -1180 21610
rect -940 21370 -850 21610
rect -610 21370 -520 21610
rect -280 21370 -190 21610
rect 50 21370 140 21610
rect 380 21370 470 21610
rect 710 21370 840 21610
rect 1080 21370 1170 21610
rect 1410 21370 1500 21610
rect 1740 21370 1830 21610
rect 2070 21370 2160 21610
rect 2400 21370 2490 21610
rect 2730 21370 2820 21610
rect 3060 21370 3150 21610
rect 3390 21370 3480 21610
rect 3720 21370 3850 21610
rect 4090 21370 4180 21610
rect 4420 21370 4510 21610
rect 4750 21370 4840 21610
rect 5080 21370 5170 21610
rect 5410 21370 5500 21610
rect 5740 21370 5830 21610
rect 6070 21370 6160 21610
rect 6400 21370 6490 21610
rect 6730 21370 6760 21610
rect -5550 20830 6760 21370
rect -5550 20590 -5200 20830
rect -4960 20590 -4870 20830
rect -4630 20590 -4540 20830
rect -4300 20590 -4210 20830
rect -3970 20590 -3880 20830
rect -3640 20590 -3550 20830
rect -3310 20590 -3220 20830
rect -2980 20590 -2890 20830
rect -2650 20590 -2560 20830
rect -2320 20590 -2230 20830
rect -1990 20590 -1900 20830
rect -1660 20590 -1570 20830
rect -1330 20590 -1240 20830
rect -1000 20590 -910 20830
rect -670 20590 -580 20830
rect -340 20590 -250 20830
rect -10 20590 80 20830
rect 320 20590 410 20830
rect 650 20590 740 20830
rect 980 20590 1070 20830
rect 1310 20590 1400 20830
rect 1640 20590 1730 20830
rect 1970 20590 2060 20830
rect 2300 20590 2390 20830
rect 2630 20590 2720 20830
rect 2960 20590 3050 20830
rect 3290 20590 3380 20830
rect 3620 20590 3710 20830
rect 3950 20590 4040 20830
rect 4280 20590 4370 20830
rect 4610 20590 4700 20830
rect 4940 20590 5030 20830
rect 5270 20590 5360 20830
rect 5600 20590 5690 20830
rect 5930 20590 6020 20830
rect 6260 20590 6350 20830
rect 6590 20590 6760 20830
rect -5550 20500 6760 20590
rect -5550 20260 -5200 20500
rect -4960 20260 -4870 20500
rect -4630 20260 -4540 20500
rect -4300 20260 -4210 20500
rect -3970 20260 -3880 20500
rect -3640 20260 -3550 20500
rect -3310 20260 -3220 20500
rect -2980 20260 -2890 20500
rect -2650 20260 -2560 20500
rect -2320 20260 -2230 20500
rect -1990 20260 -1900 20500
rect -1660 20260 -1570 20500
rect -1330 20260 -1240 20500
rect -1000 20260 -910 20500
rect -670 20260 -580 20500
rect -340 20260 -250 20500
rect -10 20260 80 20500
rect 320 20260 410 20500
rect 650 20260 740 20500
rect 980 20260 1070 20500
rect 1310 20260 1400 20500
rect 1640 20260 1730 20500
rect 1970 20260 2060 20500
rect 2300 20260 2390 20500
rect 2630 20260 2720 20500
rect 2960 20260 3050 20500
rect 3290 20260 3380 20500
rect 3620 20260 3710 20500
rect 3950 20260 4040 20500
rect 4280 20260 4370 20500
rect 4610 20260 4700 20500
rect 4940 20260 5030 20500
rect 5270 20260 5360 20500
rect 5600 20260 5690 20500
rect 5930 20260 6020 20500
rect 6260 20260 6350 20500
rect 6590 20260 6760 20500
rect -5550 20170 6760 20260
rect -5550 19930 -5200 20170
rect -4960 19930 -4870 20170
rect -4630 19930 -4540 20170
rect -4300 19930 -4210 20170
rect -3970 19930 -3880 20170
rect -3640 19930 -3550 20170
rect -3310 19930 -3220 20170
rect -2980 19930 -2890 20170
rect -2650 19930 -2560 20170
rect -2320 19930 -2230 20170
rect -1990 19930 -1900 20170
rect -1660 19930 -1570 20170
rect -1330 19930 -1240 20170
rect -1000 19930 -910 20170
rect -670 19930 -580 20170
rect -340 19930 -250 20170
rect -10 19930 80 20170
rect 320 19930 410 20170
rect 650 19930 740 20170
rect 980 19930 1070 20170
rect 1310 19930 1400 20170
rect 1640 19930 1730 20170
rect 1970 19930 2060 20170
rect 2300 19930 2390 20170
rect 2630 19930 2720 20170
rect 2960 19930 3050 20170
rect 3290 19930 3380 20170
rect 3620 19930 3710 20170
rect 3950 19930 4040 20170
rect 4280 19930 4370 20170
rect 4610 19930 4700 20170
rect 4940 19930 5030 20170
rect 5270 19930 5360 20170
rect 5600 19930 5690 20170
rect 5930 19930 6020 20170
rect 6260 19930 6350 20170
rect 6590 19930 6760 20170
rect -5550 19840 6760 19930
rect -5550 19600 -5200 19840
rect -4960 19600 -4870 19840
rect -4630 19600 -4540 19840
rect -4300 19600 -4210 19840
rect -3970 19600 -3880 19840
rect -3640 19600 -3550 19840
rect -3310 19600 -3220 19840
rect -2980 19600 -2890 19840
rect -2650 19600 -2560 19840
rect -2320 19600 -2230 19840
rect -1990 19600 -1900 19840
rect -1660 19600 -1570 19840
rect -1330 19600 -1240 19840
rect -1000 19600 -910 19840
rect -670 19600 -580 19840
rect -340 19600 -250 19840
rect -10 19600 80 19840
rect 320 19600 410 19840
rect 650 19600 740 19840
rect 980 19600 1070 19840
rect 1310 19600 1400 19840
rect 1640 19600 1730 19840
rect 1970 19600 2060 19840
rect 2300 19600 2390 19840
rect 2630 19600 2720 19840
rect 2960 19600 3050 19840
rect 3290 19600 3380 19840
rect 3620 19600 3710 19840
rect 3950 19600 4040 19840
rect 4280 19600 4370 19840
rect 4610 19600 4700 19840
rect 4940 19600 5030 19840
rect 5270 19600 5360 19840
rect 5600 19600 5690 19840
rect 5930 19600 6020 19840
rect 6260 19600 6350 19840
rect 6590 19600 6760 19840
rect -5550 19510 6760 19600
rect -5550 19270 -5200 19510
rect -4960 19270 -4870 19510
rect -4630 19270 -4540 19510
rect -4300 19270 -4210 19510
rect -3970 19270 -3880 19510
rect -3640 19270 -3550 19510
rect -3310 19270 -3220 19510
rect -2980 19270 -2890 19510
rect -2650 19270 -2560 19510
rect -2320 19270 -2230 19510
rect -1990 19270 -1900 19510
rect -1660 19270 -1570 19510
rect -1330 19270 -1240 19510
rect -1000 19270 -910 19510
rect -670 19270 -580 19510
rect -340 19270 -250 19510
rect -10 19270 80 19510
rect 320 19270 410 19510
rect 650 19270 740 19510
rect 980 19270 1070 19510
rect 1310 19270 1400 19510
rect 1640 19270 1730 19510
rect 1970 19270 2060 19510
rect 2300 19270 2390 19510
rect 2630 19270 2720 19510
rect 2960 19270 3050 19510
rect 3290 19270 3380 19510
rect 3620 19270 3710 19510
rect 3950 19270 4040 19510
rect 4280 19270 4370 19510
rect 4610 19270 4700 19510
rect 4940 19270 5030 19510
rect 5270 19270 5360 19510
rect 5600 19270 5690 19510
rect 5930 19270 6020 19510
rect 6260 19270 6350 19510
rect 6590 19270 6760 19510
rect -5550 19180 6760 19270
rect -5550 18940 -5200 19180
rect -4960 18940 -4870 19180
rect -4630 18940 -4540 19180
rect -4300 18940 -4210 19180
rect -3970 18940 -3880 19180
rect -3640 18940 -3550 19180
rect -3310 18940 -3220 19180
rect -2980 18940 -2890 19180
rect -2650 18940 -2560 19180
rect -2320 18940 -2230 19180
rect -1990 18940 -1900 19180
rect -1660 18940 -1570 19180
rect -1330 18940 -1240 19180
rect -1000 18940 -910 19180
rect -670 18940 -580 19180
rect -340 18940 -250 19180
rect -10 18940 80 19180
rect 320 18940 410 19180
rect 650 18940 740 19180
rect 980 18940 1070 19180
rect 1310 18940 1400 19180
rect 1640 18940 1730 19180
rect 1970 18940 2060 19180
rect 2300 18940 2390 19180
rect 2630 18940 2720 19180
rect 2960 18940 3050 19180
rect 3290 18940 3380 19180
rect 3620 18940 3710 19180
rect 3950 18940 4040 19180
rect 4280 18940 4370 19180
rect 4610 18940 4700 19180
rect 4940 18940 5030 19180
rect 5270 18940 5360 19180
rect 5600 18940 5690 19180
rect 5930 18940 6020 19180
rect 6260 18940 6350 19180
rect 6590 18940 6760 19180
rect -5550 18850 6760 18940
rect -5550 18610 -5200 18850
rect -4960 18610 -4870 18850
rect -4630 18610 -4540 18850
rect -4300 18610 -4210 18850
rect -3970 18610 -3880 18850
rect -3640 18610 -3550 18850
rect -3310 18610 -3220 18850
rect -2980 18610 -2890 18850
rect -2650 18610 -2560 18850
rect -2320 18610 -2230 18850
rect -1990 18610 -1900 18850
rect -1660 18610 -1570 18850
rect -1330 18610 -1240 18850
rect -1000 18610 -910 18850
rect -670 18610 -580 18850
rect -340 18610 -250 18850
rect -10 18610 80 18850
rect 320 18610 410 18850
rect 650 18610 740 18850
rect 980 18610 1070 18850
rect 1310 18610 1400 18850
rect 1640 18610 1730 18850
rect 1970 18610 2060 18850
rect 2300 18610 2390 18850
rect 2630 18610 2720 18850
rect 2960 18610 3050 18850
rect 3290 18610 3380 18850
rect 3620 18610 3710 18850
rect 3950 18610 4040 18850
rect 4280 18610 4370 18850
rect 4610 18610 4700 18850
rect 4940 18610 5030 18850
rect 5270 18610 5360 18850
rect 5600 18610 5690 18850
rect 5930 18610 6020 18850
rect 6260 18610 6350 18850
rect 6590 18610 6760 18850
rect -5550 18520 6760 18610
rect -5550 18280 -5200 18520
rect -4960 18280 -4870 18520
rect -4630 18280 -4540 18520
rect -4300 18280 -4210 18520
rect -3970 18280 -3880 18520
rect -3640 18280 -3550 18520
rect -3310 18280 -3220 18520
rect -2980 18280 -2890 18520
rect -2650 18280 -2560 18520
rect -2320 18280 -2230 18520
rect -1990 18280 -1900 18520
rect -1660 18280 -1570 18520
rect -1330 18280 -1240 18520
rect -1000 18280 -910 18520
rect -670 18280 -580 18520
rect -340 18280 -250 18520
rect -10 18280 80 18520
rect 320 18280 410 18520
rect 650 18280 740 18520
rect 980 18280 1070 18520
rect 1310 18280 1400 18520
rect 1640 18280 1730 18520
rect 1970 18280 2060 18520
rect 2300 18280 2390 18520
rect 2630 18280 2720 18520
rect 2960 18280 3050 18520
rect 3290 18280 3380 18520
rect 3620 18280 3710 18520
rect 3950 18280 4040 18520
rect 4280 18280 4370 18520
rect 4610 18280 4700 18520
rect 4940 18280 5030 18520
rect 5270 18280 5360 18520
rect 5600 18280 5690 18520
rect 5930 18280 6020 18520
rect 6260 18280 6350 18520
rect 6590 18280 6760 18520
rect -5550 18190 6760 18280
rect -5550 17950 -5200 18190
rect -4960 17950 -4870 18190
rect -4630 17950 -4540 18190
rect -4300 17950 -4210 18190
rect -3970 17950 -3880 18190
rect -3640 17950 -3550 18190
rect -3310 17950 -3220 18190
rect -2980 17950 -2890 18190
rect -2650 17950 -2560 18190
rect -2320 17950 -2230 18190
rect -1990 17950 -1900 18190
rect -1660 17950 -1570 18190
rect -1330 17950 -1240 18190
rect -1000 17950 -910 18190
rect -670 17950 -580 18190
rect -340 17950 -250 18190
rect -10 17950 80 18190
rect 320 17950 410 18190
rect 650 17950 740 18190
rect 980 17950 1070 18190
rect 1310 17950 1400 18190
rect 1640 17950 1730 18190
rect 1970 17950 2060 18190
rect 2300 17950 2390 18190
rect 2630 17950 2720 18190
rect 2960 17950 3050 18190
rect 3290 17950 3380 18190
rect 3620 17950 3710 18190
rect 3950 17950 4040 18190
rect 4280 17950 4370 18190
rect 4610 17950 4700 18190
rect 4940 17950 5030 18190
rect 5270 17950 5360 18190
rect 5600 17950 5690 18190
rect 5930 17950 6020 18190
rect 6260 17950 6350 18190
rect 6590 17950 6760 18190
rect -5550 17860 6760 17950
rect -5550 17620 -5200 17860
rect -4960 17620 -4870 17860
rect -4630 17620 -4540 17860
rect -4300 17620 -4210 17860
rect -3970 17620 -3880 17860
rect -3640 17620 -3550 17860
rect -3310 17620 -3220 17860
rect -2980 17620 -2890 17860
rect -2650 17620 -2560 17860
rect -2320 17620 -2230 17860
rect -1990 17620 -1900 17860
rect -1660 17620 -1570 17860
rect -1330 17620 -1240 17860
rect -1000 17620 -910 17860
rect -670 17620 -580 17860
rect -340 17620 -250 17860
rect -10 17620 80 17860
rect 320 17620 410 17860
rect 650 17620 740 17860
rect 980 17620 1070 17860
rect 1310 17620 1400 17860
rect 1640 17620 1730 17860
rect 1970 17620 2060 17860
rect 2300 17620 2390 17860
rect 2630 17620 2720 17860
rect 2960 17620 3050 17860
rect 3290 17620 3380 17860
rect 3620 17620 3710 17860
rect 3950 17620 4040 17860
rect 4280 17620 4370 17860
rect 4610 17620 4700 17860
rect 4940 17620 5030 17860
rect 5270 17620 5360 17860
rect 5600 17620 5690 17860
rect 5930 17620 6020 17860
rect 6260 17620 6350 17860
rect 6590 17620 6760 17860
rect -5550 17530 6760 17620
rect -5550 17290 -5200 17530
rect -4960 17290 -4870 17530
rect -4630 17290 -4540 17530
rect -4300 17290 -4210 17530
rect -3970 17290 -3880 17530
rect -3640 17290 -3550 17530
rect -3310 17290 -3220 17530
rect -2980 17290 -2890 17530
rect -2650 17290 -2560 17530
rect -2320 17290 -2230 17530
rect -1990 17290 -1900 17530
rect -1660 17290 -1570 17530
rect -1330 17290 -1240 17530
rect -1000 17290 -910 17530
rect -670 17290 -580 17530
rect -340 17290 -250 17530
rect -10 17290 80 17530
rect 320 17290 410 17530
rect 650 17290 740 17530
rect 980 17290 1070 17530
rect 1310 17290 1400 17530
rect 1640 17290 1730 17530
rect 1970 17290 2060 17530
rect 2300 17290 2390 17530
rect 2630 17290 2720 17530
rect 2960 17290 3050 17530
rect 3290 17290 3380 17530
rect 3620 17290 3710 17530
rect 3950 17290 4040 17530
rect 4280 17290 4370 17530
rect 4610 17290 4700 17530
rect 4940 17290 5030 17530
rect 5270 17290 5360 17530
rect 5600 17290 5690 17530
rect 5930 17290 6020 17530
rect 6260 17290 6350 17530
rect 6590 17290 6760 17530
rect -5550 17200 6760 17290
rect -5550 16960 -5200 17200
rect -4960 16960 -4870 17200
rect -4630 16960 -4540 17200
rect -4300 16960 -4210 17200
rect -3970 16960 -3880 17200
rect -3640 16960 -3550 17200
rect -3310 16960 -3220 17200
rect -2980 16960 -2890 17200
rect -2650 16960 -2560 17200
rect -2320 16960 -2230 17200
rect -1990 16960 -1900 17200
rect -1660 16960 -1570 17200
rect -1330 16960 -1240 17200
rect -1000 16960 -910 17200
rect -670 16960 -580 17200
rect -340 16960 -250 17200
rect -10 16960 80 17200
rect 320 16960 410 17200
rect 650 16960 740 17200
rect 980 16960 1070 17200
rect 1310 16960 1400 17200
rect 1640 16960 1730 17200
rect 1970 16960 2060 17200
rect 2300 16960 2390 17200
rect 2630 16960 2720 17200
rect 2960 16960 3050 17200
rect 3290 16960 3380 17200
rect 3620 16960 3710 17200
rect 3950 16960 4040 17200
rect 4280 16960 4370 17200
rect 4610 16960 4700 17200
rect 4940 16960 5030 17200
rect 5270 16960 5360 17200
rect 5600 16960 5690 17200
rect 5930 16960 6020 17200
rect 6260 16960 6350 17200
rect 6590 16960 6760 17200
rect -5550 16870 6760 16960
rect -5550 16630 -5200 16870
rect -4960 16630 -4870 16870
rect -4630 16630 -4540 16870
rect -4300 16630 -4210 16870
rect -3970 16630 -3880 16870
rect -3640 16630 -3550 16870
rect -3310 16630 -3220 16870
rect -2980 16630 -2890 16870
rect -2650 16630 -2560 16870
rect -2320 16630 -2230 16870
rect -1990 16630 -1900 16870
rect -1660 16630 -1570 16870
rect -1330 16630 -1240 16870
rect -1000 16630 -910 16870
rect -670 16630 -580 16870
rect -340 16630 -250 16870
rect -10 16630 80 16870
rect 320 16630 410 16870
rect 650 16630 740 16870
rect 980 16630 1070 16870
rect 1310 16630 1400 16870
rect 1640 16630 1730 16870
rect 1970 16630 2060 16870
rect 2300 16630 2390 16870
rect 2630 16630 2720 16870
rect 2960 16630 3050 16870
rect 3290 16630 3380 16870
rect 3620 16630 3710 16870
rect 3950 16630 4040 16870
rect 4280 16630 4370 16870
rect 4610 16630 4700 16870
rect 4940 16630 5030 16870
rect 5270 16630 5360 16870
rect 5600 16630 5690 16870
rect 5930 16630 6020 16870
rect 6260 16630 6350 16870
rect 6590 16630 6760 16870
rect -5550 16540 6760 16630
rect -5550 16300 -5200 16540
rect -4960 16300 -4870 16540
rect -4630 16300 -4540 16540
rect -4300 16300 -4210 16540
rect -3970 16300 -3880 16540
rect -3640 16300 -3550 16540
rect -3310 16300 -3220 16540
rect -2980 16300 -2890 16540
rect -2650 16300 -2560 16540
rect -2320 16300 -2230 16540
rect -1990 16300 -1900 16540
rect -1660 16300 -1570 16540
rect -1330 16300 -1240 16540
rect -1000 16300 -910 16540
rect -670 16300 -580 16540
rect -340 16300 -250 16540
rect -10 16300 80 16540
rect 320 16300 410 16540
rect 650 16300 740 16540
rect 980 16300 1070 16540
rect 1310 16300 1400 16540
rect 1640 16300 1730 16540
rect 1970 16300 2060 16540
rect 2300 16300 2390 16540
rect 2630 16300 2720 16540
rect 2960 16300 3050 16540
rect 3290 16300 3380 16540
rect 3620 16300 3710 16540
rect 3950 16300 4040 16540
rect 4280 16300 4370 16540
rect 4610 16300 4700 16540
rect 4940 16300 5030 16540
rect 5270 16300 5360 16540
rect 5600 16300 5690 16540
rect 5930 16300 6020 16540
rect 6260 16300 6350 16540
rect 6590 16300 6760 16540
rect -5550 16210 6760 16300
rect -5550 15970 -5200 16210
rect -4960 15970 -4870 16210
rect -4630 15970 -4540 16210
rect -4300 15970 -4210 16210
rect -3970 15970 -3880 16210
rect -3640 15970 -3550 16210
rect -3310 15970 -3220 16210
rect -2980 15970 -2890 16210
rect -2650 15970 -2560 16210
rect -2320 15970 -2230 16210
rect -1990 15970 -1900 16210
rect -1660 15970 -1570 16210
rect -1330 15970 -1240 16210
rect -1000 15970 -910 16210
rect -670 15970 -580 16210
rect -340 15970 -250 16210
rect -10 15970 80 16210
rect 320 15970 410 16210
rect 650 15970 740 16210
rect 980 15970 1070 16210
rect 1310 15970 1400 16210
rect 1640 15970 1730 16210
rect 1970 15970 2060 16210
rect 2300 15970 2390 16210
rect 2630 15970 2720 16210
rect 2960 15970 3050 16210
rect 3290 15970 3380 16210
rect 3620 15970 3710 16210
rect 3950 15970 4040 16210
rect 4280 15970 4370 16210
rect 4610 15970 4700 16210
rect 4940 15970 5030 16210
rect 5270 15970 5360 16210
rect 5600 15970 5690 16210
rect 5930 15970 6020 16210
rect 6260 15970 6350 16210
rect 6590 15970 6760 16210
rect -5550 15880 6760 15970
rect -5550 15640 -5200 15880
rect -4960 15640 -4870 15880
rect -4630 15640 -4540 15880
rect -4300 15640 -4210 15880
rect -3970 15640 -3880 15880
rect -3640 15640 -3550 15880
rect -3310 15640 -3220 15880
rect -2980 15640 -2890 15880
rect -2650 15640 -2560 15880
rect -2320 15640 -2230 15880
rect -1990 15640 -1900 15880
rect -1660 15640 -1570 15880
rect -1330 15640 -1240 15880
rect -1000 15640 -910 15880
rect -670 15640 -580 15880
rect -340 15640 -250 15880
rect -10 15640 80 15880
rect 320 15640 410 15880
rect 650 15640 740 15880
rect 980 15640 1070 15880
rect 1310 15640 1400 15880
rect 1640 15640 1730 15880
rect 1970 15640 2060 15880
rect 2300 15640 2390 15880
rect 2630 15640 2720 15880
rect 2960 15640 3050 15880
rect 3290 15640 3380 15880
rect 3620 15640 3710 15880
rect 3950 15640 4040 15880
rect 4280 15640 4370 15880
rect 4610 15640 4700 15880
rect 4940 15640 5030 15880
rect 5270 15640 5360 15880
rect 5600 15640 5690 15880
rect 5930 15640 6020 15880
rect 6260 15640 6350 15880
rect 6590 15640 6760 15880
rect -5550 15550 6760 15640
rect -5550 15310 -5200 15550
rect -4960 15310 -4870 15550
rect -4630 15310 -4540 15550
rect -4300 15310 -4210 15550
rect -3970 15310 -3880 15550
rect -3640 15310 -3550 15550
rect -3310 15310 -3220 15550
rect -2980 15310 -2890 15550
rect -2650 15310 -2560 15550
rect -2320 15310 -2230 15550
rect -1990 15310 -1900 15550
rect -1660 15310 -1570 15550
rect -1330 15310 -1240 15550
rect -1000 15310 -910 15550
rect -670 15310 -580 15550
rect -340 15310 -250 15550
rect -10 15310 80 15550
rect 320 15310 410 15550
rect 650 15310 740 15550
rect 980 15310 1070 15550
rect 1310 15310 1400 15550
rect 1640 15310 1730 15550
rect 1970 15310 2060 15550
rect 2300 15310 2390 15550
rect 2630 15310 2720 15550
rect 2960 15310 3050 15550
rect 3290 15310 3380 15550
rect 3620 15310 3710 15550
rect 3950 15310 4040 15550
rect 4280 15310 4370 15550
rect 4610 15310 4700 15550
rect 4940 15310 5030 15550
rect 5270 15310 5360 15550
rect 5600 15310 5690 15550
rect 5930 15310 6020 15550
rect 6260 15310 6350 15550
rect 6590 15310 6760 15550
rect -5550 15220 6760 15310
rect -5550 14980 -5200 15220
rect -4960 14980 -4870 15220
rect -4630 14980 -4540 15220
rect -4300 14980 -4210 15220
rect -3970 14980 -3880 15220
rect -3640 14980 -3550 15220
rect -3310 14980 -3220 15220
rect -2980 14980 -2890 15220
rect -2650 14980 -2560 15220
rect -2320 14980 -2230 15220
rect -1990 14980 -1900 15220
rect -1660 14980 -1570 15220
rect -1330 14980 -1240 15220
rect -1000 14980 -910 15220
rect -670 14980 -580 15220
rect -340 14980 -250 15220
rect -10 14980 80 15220
rect 320 14980 410 15220
rect 650 14980 740 15220
rect 980 14980 1070 15220
rect 1310 14980 1400 15220
rect 1640 14980 1730 15220
rect 1970 14980 2060 15220
rect 2300 14980 2390 15220
rect 2630 14980 2720 15220
rect 2960 14980 3050 15220
rect 3290 14980 3380 15220
rect 3620 14980 3710 15220
rect 3950 14980 4040 15220
rect 4280 14980 4370 15220
rect 4610 14980 4700 15220
rect 4940 14980 5030 15220
rect 5270 14980 5360 15220
rect 5600 14980 5690 15220
rect 5930 14980 6020 15220
rect 6260 14980 6350 15220
rect 6590 14980 6760 15220
rect -5550 14890 6760 14980
rect -5550 14650 -5200 14890
rect -4960 14650 -4870 14890
rect -4630 14650 -4540 14890
rect -4300 14650 -4210 14890
rect -3970 14650 -3880 14890
rect -3640 14650 -3550 14890
rect -3310 14650 -3220 14890
rect -2980 14650 -2890 14890
rect -2650 14650 -2560 14890
rect -2320 14650 -2230 14890
rect -1990 14650 -1900 14890
rect -1660 14650 -1570 14890
rect -1330 14650 -1240 14890
rect -1000 14650 -910 14890
rect -670 14650 -580 14890
rect -340 14650 -250 14890
rect -10 14650 80 14890
rect 320 14650 410 14890
rect 650 14650 740 14890
rect 980 14650 1070 14890
rect 1310 14650 1400 14890
rect 1640 14650 1730 14890
rect 1970 14650 2060 14890
rect 2300 14650 2390 14890
rect 2630 14650 2720 14890
rect 2960 14650 3050 14890
rect 3290 14650 3380 14890
rect 3620 14650 3710 14890
rect 3950 14650 4040 14890
rect 4280 14650 4370 14890
rect 4610 14650 4700 14890
rect 4940 14650 5030 14890
rect 5270 14650 5360 14890
rect 5600 14650 5690 14890
rect 5930 14650 6020 14890
rect 6260 14650 6350 14890
rect 6590 14650 6760 14890
rect -5550 14560 6760 14650
rect -5550 14320 -5200 14560
rect -4960 14320 -4870 14560
rect -4630 14320 -4540 14560
rect -4300 14320 -4210 14560
rect -3970 14320 -3880 14560
rect -3640 14320 -3550 14560
rect -3310 14320 -3220 14560
rect -2980 14320 -2890 14560
rect -2650 14320 -2560 14560
rect -2320 14320 -2230 14560
rect -1990 14320 -1900 14560
rect -1660 14320 -1570 14560
rect -1330 14320 -1240 14560
rect -1000 14320 -910 14560
rect -670 14320 -580 14560
rect -340 14320 -250 14560
rect -10 14320 80 14560
rect 320 14320 410 14560
rect 650 14320 740 14560
rect 980 14320 1070 14560
rect 1310 14320 1400 14560
rect 1640 14320 1730 14560
rect 1970 14320 2060 14560
rect 2300 14320 2390 14560
rect 2630 14320 2720 14560
rect 2960 14320 3050 14560
rect 3290 14320 3380 14560
rect 3620 14320 3710 14560
rect 3950 14320 4040 14560
rect 4280 14320 4370 14560
rect 4610 14320 4700 14560
rect 4940 14320 5030 14560
rect 5270 14320 5360 14560
rect 5600 14320 5690 14560
rect 5930 14320 6020 14560
rect 6260 14320 6350 14560
rect 6590 14320 6760 14560
rect -5550 14230 6760 14320
rect -5550 13990 -5200 14230
rect -4960 13990 -4870 14230
rect -4630 13990 -4540 14230
rect -4300 13990 -4210 14230
rect -3970 13990 -3880 14230
rect -3640 13990 -3550 14230
rect -3310 13990 -3220 14230
rect -2980 13990 -2890 14230
rect -2650 13990 -2560 14230
rect -2320 13990 -2230 14230
rect -1990 13990 -1900 14230
rect -1660 13990 -1570 14230
rect -1330 13990 -1240 14230
rect -1000 13990 -910 14230
rect -670 13990 -580 14230
rect -340 13990 -250 14230
rect -10 13990 80 14230
rect 320 13990 410 14230
rect 650 13990 740 14230
rect 980 13990 1070 14230
rect 1310 13990 1400 14230
rect 1640 13990 1730 14230
rect 1970 13990 2060 14230
rect 2300 13990 2390 14230
rect 2630 13990 2720 14230
rect 2960 13990 3050 14230
rect 3290 13990 3380 14230
rect 3620 13990 3710 14230
rect 3950 13990 4040 14230
rect 4280 13990 4370 14230
rect 4610 13990 4700 14230
rect 4940 13990 5030 14230
rect 5270 13990 5360 14230
rect 5600 13990 5690 14230
rect 5930 13990 6020 14230
rect 6260 13990 6350 14230
rect 6590 13990 6760 14230
rect -5550 13900 6760 13990
rect -5550 13660 -5200 13900
rect -4960 13660 -4870 13900
rect -4630 13660 -4540 13900
rect -4300 13660 -4210 13900
rect -3970 13660 -3880 13900
rect -3640 13660 -3550 13900
rect -3310 13660 -3220 13900
rect -2980 13660 -2890 13900
rect -2650 13660 -2560 13900
rect -2320 13660 -2230 13900
rect -1990 13660 -1900 13900
rect -1660 13660 -1570 13900
rect -1330 13660 -1240 13900
rect -1000 13660 -910 13900
rect -670 13660 -580 13900
rect -340 13660 -250 13900
rect -10 13660 80 13900
rect 320 13660 410 13900
rect 650 13660 740 13900
rect 980 13660 1070 13900
rect 1310 13660 1400 13900
rect 1640 13660 1730 13900
rect 1970 13660 2060 13900
rect 2300 13660 2390 13900
rect 2630 13660 2720 13900
rect 2960 13660 3050 13900
rect 3290 13660 3380 13900
rect 3620 13660 3710 13900
rect 3950 13660 4040 13900
rect 4280 13660 4370 13900
rect 4610 13660 4700 13900
rect 4940 13660 5030 13900
rect 5270 13660 5360 13900
rect 5600 13660 5690 13900
rect 5930 13660 6020 13900
rect 6260 13660 6350 13900
rect 6590 13660 6760 13900
rect -5550 13570 6760 13660
rect -5550 13330 -5200 13570
rect -4960 13330 -4870 13570
rect -4630 13330 -4540 13570
rect -4300 13330 -4210 13570
rect -3970 13330 -3880 13570
rect -3640 13330 -3550 13570
rect -3310 13330 -3220 13570
rect -2980 13330 -2890 13570
rect -2650 13330 -2560 13570
rect -2320 13330 -2230 13570
rect -1990 13330 -1900 13570
rect -1660 13330 -1570 13570
rect -1330 13330 -1240 13570
rect -1000 13330 -910 13570
rect -670 13330 -580 13570
rect -340 13330 -250 13570
rect -10 13330 80 13570
rect 320 13330 410 13570
rect 650 13330 740 13570
rect 980 13330 1070 13570
rect 1310 13330 1400 13570
rect 1640 13330 1730 13570
rect 1970 13330 2060 13570
rect 2300 13330 2390 13570
rect 2630 13330 2720 13570
rect 2960 13330 3050 13570
rect 3290 13330 3380 13570
rect 3620 13330 3710 13570
rect 3950 13330 4040 13570
rect 4280 13330 4370 13570
rect 4610 13330 4700 13570
rect 4940 13330 5030 13570
rect 5270 13330 5360 13570
rect 5600 13330 5690 13570
rect 5930 13330 6020 13570
rect 6260 13330 6350 13570
rect 6590 13330 6760 13570
rect -5550 13240 6760 13330
rect -5550 13000 -5200 13240
rect -4960 13000 -4870 13240
rect -4630 13000 -4540 13240
rect -4300 13000 -4210 13240
rect -3970 13000 -3880 13240
rect -3640 13000 -3550 13240
rect -3310 13000 -3220 13240
rect -2980 13000 -2890 13240
rect -2650 13000 -2560 13240
rect -2320 13000 -2230 13240
rect -1990 13000 -1900 13240
rect -1660 13000 -1570 13240
rect -1330 13000 -1240 13240
rect -1000 13000 -910 13240
rect -670 13000 -580 13240
rect -340 13000 -250 13240
rect -10 13000 80 13240
rect 320 13000 410 13240
rect 650 13000 740 13240
rect 980 13000 1070 13240
rect 1310 13000 1400 13240
rect 1640 13000 1730 13240
rect 1970 13000 2060 13240
rect 2300 13000 2390 13240
rect 2630 13000 2720 13240
rect 2960 13000 3050 13240
rect 3290 13000 3380 13240
rect 3620 13000 3710 13240
rect 3950 13000 4040 13240
rect 4280 13000 4370 13240
rect 4610 13000 4700 13240
rect 4940 13000 5030 13240
rect 5270 13000 5360 13240
rect 5600 13000 5690 13240
rect 5930 13000 6020 13240
rect 6260 13000 6350 13240
rect 6590 13000 6760 13240
rect -5550 12910 6760 13000
rect -5550 12670 -5200 12910
rect -4960 12670 -4870 12910
rect -4630 12670 -4540 12910
rect -4300 12670 -4210 12910
rect -3970 12670 -3880 12910
rect -3640 12670 -3550 12910
rect -3310 12670 -3220 12910
rect -2980 12670 -2890 12910
rect -2650 12670 -2560 12910
rect -2320 12670 -2230 12910
rect -1990 12670 -1900 12910
rect -1660 12670 -1570 12910
rect -1330 12670 -1240 12910
rect -1000 12670 -910 12910
rect -670 12670 -580 12910
rect -340 12670 -250 12910
rect -10 12670 80 12910
rect 320 12670 410 12910
rect 650 12670 740 12910
rect 980 12670 1070 12910
rect 1310 12670 1400 12910
rect 1640 12670 1730 12910
rect 1970 12670 2060 12910
rect 2300 12670 2390 12910
rect 2630 12670 2720 12910
rect 2960 12670 3050 12910
rect 3290 12670 3380 12910
rect 3620 12670 3710 12910
rect 3950 12670 4040 12910
rect 4280 12670 4370 12910
rect 4610 12670 4700 12910
rect 4940 12670 5030 12910
rect 5270 12670 5360 12910
rect 5600 12670 5690 12910
rect 5930 12670 6020 12910
rect 6260 12670 6350 12910
rect 6590 12670 6760 12910
rect -5550 12580 6760 12670
rect -5550 12340 -5200 12580
rect -4960 12340 -4870 12580
rect -4630 12340 -4540 12580
rect -4300 12340 -4210 12580
rect -3970 12340 -3880 12580
rect -3640 12340 -3550 12580
rect -3310 12340 -3220 12580
rect -2980 12340 -2890 12580
rect -2650 12340 -2560 12580
rect -2320 12340 -2230 12580
rect -1990 12340 -1900 12580
rect -1660 12340 -1570 12580
rect -1330 12340 -1240 12580
rect -1000 12340 -910 12580
rect -670 12340 -580 12580
rect -340 12340 -250 12580
rect -10 12340 80 12580
rect 320 12340 410 12580
rect 650 12340 740 12580
rect 980 12340 1070 12580
rect 1310 12340 1400 12580
rect 1640 12340 1730 12580
rect 1970 12340 2060 12580
rect 2300 12340 2390 12580
rect 2630 12340 2720 12580
rect 2960 12340 3050 12580
rect 3290 12340 3380 12580
rect 3620 12340 3710 12580
rect 3950 12340 4040 12580
rect 4280 12340 4370 12580
rect 4610 12340 4700 12580
rect 4940 12340 5030 12580
rect 5270 12340 5360 12580
rect 5600 12340 5690 12580
rect 5930 12340 6020 12580
rect 6260 12340 6350 12580
rect 6590 12340 6760 12580
rect -5550 12250 6760 12340
rect -5550 12010 -5200 12250
rect -4960 12010 -4870 12250
rect -4630 12010 -4540 12250
rect -4300 12010 -4210 12250
rect -3970 12010 -3880 12250
rect -3640 12010 -3550 12250
rect -3310 12010 -3220 12250
rect -2980 12010 -2890 12250
rect -2650 12010 -2560 12250
rect -2320 12010 -2230 12250
rect -1990 12010 -1900 12250
rect -1660 12010 -1570 12250
rect -1330 12010 -1240 12250
rect -1000 12010 -910 12250
rect -670 12010 -580 12250
rect -340 12010 -250 12250
rect -10 12010 80 12250
rect 320 12010 410 12250
rect 650 12010 740 12250
rect 980 12010 1070 12250
rect 1310 12010 1400 12250
rect 1640 12010 1730 12250
rect 1970 12010 2060 12250
rect 2300 12010 2390 12250
rect 2630 12010 2720 12250
rect 2960 12010 3050 12250
rect 3290 12010 3380 12250
rect 3620 12010 3710 12250
rect 3950 12010 4040 12250
rect 4280 12010 4370 12250
rect 4610 12010 4700 12250
rect 4940 12010 5030 12250
rect 5270 12010 5360 12250
rect 5600 12010 5690 12250
rect 5930 12010 6020 12250
rect 6260 12010 6350 12250
rect 6590 12010 6760 12250
rect -5550 11920 6760 12010
rect -5550 11680 -5200 11920
rect -4960 11680 -4870 11920
rect -4630 11680 -4540 11920
rect -4300 11680 -4210 11920
rect -3970 11680 -3880 11920
rect -3640 11680 -3550 11920
rect -3310 11680 -3220 11920
rect -2980 11680 -2890 11920
rect -2650 11680 -2560 11920
rect -2320 11680 -2230 11920
rect -1990 11680 -1900 11920
rect -1660 11680 -1570 11920
rect -1330 11680 -1240 11920
rect -1000 11680 -910 11920
rect -670 11680 -580 11920
rect -340 11680 -250 11920
rect -10 11680 80 11920
rect 320 11680 410 11920
rect 650 11680 740 11920
rect 980 11680 1070 11920
rect 1310 11680 1400 11920
rect 1640 11680 1730 11920
rect 1970 11680 2060 11920
rect 2300 11680 2390 11920
rect 2630 11680 2720 11920
rect 2960 11680 3050 11920
rect 3290 11680 3380 11920
rect 3620 11680 3710 11920
rect 3950 11680 4040 11920
rect 4280 11680 4370 11920
rect 4610 11680 4700 11920
rect 4940 11680 5030 11920
rect 5270 11680 5360 11920
rect 5600 11680 5690 11920
rect 5930 11680 6020 11920
rect 6260 11680 6350 11920
rect 6590 11680 6760 11920
rect -5550 11590 6760 11680
rect -5550 11350 -5200 11590
rect -4960 11350 -4870 11590
rect -4630 11350 -4540 11590
rect -4300 11350 -4210 11590
rect -3970 11350 -3880 11590
rect -3640 11350 -3550 11590
rect -3310 11350 -3220 11590
rect -2980 11350 -2890 11590
rect -2650 11350 -2560 11590
rect -2320 11350 -2230 11590
rect -1990 11350 -1900 11590
rect -1660 11350 -1570 11590
rect -1330 11350 -1240 11590
rect -1000 11350 -910 11590
rect -670 11350 -580 11590
rect -340 11350 -250 11590
rect -10 11350 80 11590
rect 320 11350 410 11590
rect 650 11350 740 11590
rect 980 11350 1070 11590
rect 1310 11350 1400 11590
rect 1640 11350 1730 11590
rect 1970 11350 2060 11590
rect 2300 11350 2390 11590
rect 2630 11350 2720 11590
rect 2960 11350 3050 11590
rect 3290 11350 3380 11590
rect 3620 11350 3710 11590
rect 3950 11350 4040 11590
rect 4280 11350 4370 11590
rect 4610 11350 4700 11590
rect 4940 11350 5030 11590
rect 5270 11350 5360 11590
rect 5600 11350 5690 11590
rect 5930 11350 6020 11590
rect 6260 11350 6350 11590
rect 6590 11350 6760 11590
rect -5550 11260 6760 11350
rect -5550 11020 -5200 11260
rect -4960 11020 -4870 11260
rect -4630 11020 -4540 11260
rect -4300 11020 -4210 11260
rect -3970 11020 -3880 11260
rect -3640 11020 -3550 11260
rect -3310 11020 -3220 11260
rect -2980 11020 -2890 11260
rect -2650 11020 -2560 11260
rect -2320 11020 -2230 11260
rect -1990 11020 -1900 11260
rect -1660 11020 -1570 11260
rect -1330 11020 -1240 11260
rect -1000 11020 -910 11260
rect -670 11020 -580 11260
rect -340 11020 -250 11260
rect -10 11020 80 11260
rect 320 11020 410 11260
rect 650 11020 740 11260
rect 980 11020 1070 11260
rect 1310 11020 1400 11260
rect 1640 11020 1730 11260
rect 1970 11020 2060 11260
rect 2300 11020 2390 11260
rect 2630 11020 2720 11260
rect 2960 11020 3050 11260
rect 3290 11020 3380 11260
rect 3620 11020 3710 11260
rect 3950 11020 4040 11260
rect 4280 11020 4370 11260
rect 4610 11020 4700 11260
rect 4940 11020 5030 11260
rect 5270 11020 5360 11260
rect 5600 11020 5690 11260
rect 5930 11020 6020 11260
rect 6260 11020 6350 11260
rect 6590 11020 6760 11260
rect -5550 10930 6760 11020
rect -5550 10690 -5200 10930
rect -4960 10690 -4870 10930
rect -4630 10690 -4540 10930
rect -4300 10690 -4210 10930
rect -3970 10690 -3880 10930
rect -3640 10690 -3550 10930
rect -3310 10690 -3220 10930
rect -2980 10690 -2890 10930
rect -2650 10690 -2560 10930
rect -2320 10690 -2230 10930
rect -1990 10690 -1900 10930
rect -1660 10690 -1570 10930
rect -1330 10690 -1240 10930
rect -1000 10690 -910 10930
rect -670 10690 -580 10930
rect -340 10690 -250 10930
rect -10 10690 80 10930
rect 320 10690 410 10930
rect 650 10690 740 10930
rect 980 10690 1070 10930
rect 1310 10690 1400 10930
rect 1640 10690 1730 10930
rect 1970 10690 2060 10930
rect 2300 10690 2390 10930
rect 2630 10690 2720 10930
rect 2960 10690 3050 10930
rect 3290 10690 3380 10930
rect 3620 10690 3710 10930
rect 3950 10690 4040 10930
rect 4280 10690 4370 10930
rect 4610 10690 4700 10930
rect 4940 10690 5030 10930
rect 5270 10690 5360 10930
rect 5600 10690 5690 10930
rect 5930 10690 6020 10930
rect 6260 10690 6350 10930
rect 6590 10690 6760 10930
rect -5550 10600 6760 10690
rect -5550 10360 -5200 10600
rect -4960 10360 -4870 10600
rect -4630 10360 -4540 10600
rect -4300 10360 -4210 10600
rect -3970 10360 -3880 10600
rect -3640 10360 -3550 10600
rect -3310 10360 -3220 10600
rect -2980 10360 -2890 10600
rect -2650 10360 -2560 10600
rect -2320 10360 -2230 10600
rect -1990 10360 -1900 10600
rect -1660 10360 -1570 10600
rect -1330 10360 -1240 10600
rect -1000 10360 -910 10600
rect -670 10360 -580 10600
rect -340 10360 -250 10600
rect -10 10360 80 10600
rect 320 10360 410 10600
rect 650 10360 740 10600
rect 980 10360 1070 10600
rect 1310 10360 1400 10600
rect 1640 10360 1730 10600
rect 1970 10360 2060 10600
rect 2300 10360 2390 10600
rect 2630 10360 2720 10600
rect 2960 10360 3050 10600
rect 3290 10360 3380 10600
rect 3620 10360 3710 10600
rect 3950 10360 4040 10600
rect 4280 10360 4370 10600
rect 4610 10360 4700 10600
rect 4940 10360 5030 10600
rect 5270 10360 5360 10600
rect 5600 10360 5690 10600
rect 5930 10360 6020 10600
rect 6260 10360 6350 10600
rect 6590 10360 6760 10600
rect -5550 10270 6760 10360
rect -5550 10030 -5200 10270
rect -4960 10030 -4870 10270
rect -4630 10030 -4540 10270
rect -4300 10030 -4210 10270
rect -3970 10030 -3880 10270
rect -3640 10030 -3550 10270
rect -3310 10030 -3220 10270
rect -2980 10030 -2890 10270
rect -2650 10030 -2560 10270
rect -2320 10030 -2230 10270
rect -1990 10030 -1900 10270
rect -1660 10030 -1570 10270
rect -1330 10030 -1240 10270
rect -1000 10030 -910 10270
rect -670 10030 -580 10270
rect -340 10030 -250 10270
rect -10 10030 80 10270
rect 320 10030 410 10270
rect 650 10030 740 10270
rect 980 10030 1070 10270
rect 1310 10030 1400 10270
rect 1640 10030 1730 10270
rect 1970 10030 2060 10270
rect 2300 10030 2390 10270
rect 2630 10030 2720 10270
rect 2960 10030 3050 10270
rect 3290 10030 3380 10270
rect 3620 10030 3710 10270
rect 3950 10030 4040 10270
rect 4280 10030 4370 10270
rect 4610 10030 4700 10270
rect 4940 10030 5030 10270
rect 5270 10030 5360 10270
rect 5600 10030 5690 10270
rect 5930 10030 6020 10270
rect 6260 10030 6350 10270
rect 6590 10030 6760 10270
rect -5550 9940 6760 10030
rect -5550 9700 -5200 9940
rect -4960 9700 -4870 9940
rect -4630 9700 -4540 9940
rect -4300 9700 -4210 9940
rect -3970 9700 -3880 9940
rect -3640 9700 -3550 9940
rect -3310 9700 -3220 9940
rect -2980 9700 -2890 9940
rect -2650 9700 -2560 9940
rect -2320 9700 -2230 9940
rect -1990 9700 -1900 9940
rect -1660 9700 -1570 9940
rect -1330 9700 -1240 9940
rect -1000 9700 -910 9940
rect -670 9700 -580 9940
rect -340 9700 -250 9940
rect -10 9700 80 9940
rect 320 9700 410 9940
rect 650 9700 740 9940
rect 980 9700 1070 9940
rect 1310 9700 1400 9940
rect 1640 9700 1730 9940
rect 1970 9700 2060 9940
rect 2300 9700 2390 9940
rect 2630 9700 2720 9940
rect 2960 9700 3050 9940
rect 3290 9700 3380 9940
rect 3620 9700 3710 9940
rect 3950 9700 4040 9940
rect 4280 9700 4370 9940
rect 4610 9700 4700 9940
rect 4940 9700 5030 9940
rect 5270 9700 5360 9940
rect 5600 9700 5690 9940
rect 5930 9700 6020 9940
rect 6260 9700 6350 9940
rect 6590 9700 6760 9940
rect -5550 9610 6760 9700
rect -5550 9370 -5200 9610
rect -4960 9370 -4870 9610
rect -4630 9370 -4540 9610
rect -4300 9370 -4210 9610
rect -3970 9370 -3880 9610
rect -3640 9370 -3550 9610
rect -3310 9370 -3220 9610
rect -2980 9370 -2890 9610
rect -2650 9370 -2560 9610
rect -2320 9370 -2230 9610
rect -1990 9370 -1900 9610
rect -1660 9370 -1570 9610
rect -1330 9370 -1240 9610
rect -1000 9370 -910 9610
rect -670 9370 -580 9610
rect -340 9370 -250 9610
rect -10 9370 80 9610
rect 320 9370 410 9610
rect 650 9370 740 9610
rect 980 9370 1070 9610
rect 1310 9370 1400 9610
rect 1640 9370 1730 9610
rect 1970 9370 2060 9610
rect 2300 9370 2390 9610
rect 2630 9370 2720 9610
rect 2960 9370 3050 9610
rect 3290 9370 3380 9610
rect 3620 9370 3710 9610
rect 3950 9370 4040 9610
rect 4280 9370 4370 9610
rect 4610 9370 4700 9610
rect 4940 9370 5030 9610
rect 5270 9370 5360 9610
rect 5600 9370 5690 9610
rect 5930 9370 6020 9610
rect 6260 9370 6350 9610
rect 6590 9370 6760 9610
rect -5550 9280 6760 9370
rect -5550 9040 -5200 9280
rect -4960 9040 -4870 9280
rect -4630 9040 -4540 9280
rect -4300 9040 -4210 9280
rect -3970 9040 -3880 9280
rect -3640 9040 -3550 9280
rect -3310 9040 -3220 9280
rect -2980 9040 -2890 9280
rect -2650 9040 -2560 9280
rect -2320 9040 -2230 9280
rect -1990 9040 -1900 9280
rect -1660 9040 -1570 9280
rect -1330 9040 -1240 9280
rect -1000 9040 -910 9280
rect -670 9040 -580 9280
rect -340 9040 -250 9280
rect -10 9040 80 9280
rect 320 9040 410 9280
rect 650 9040 740 9280
rect 980 9040 1070 9280
rect 1310 9040 1400 9280
rect 1640 9040 1730 9280
rect 1970 9040 2060 9280
rect 2300 9040 2390 9280
rect 2630 9040 2720 9280
rect 2960 9040 3050 9280
rect 3290 9040 3380 9280
rect 3620 9040 3710 9280
rect 3950 9040 4040 9280
rect 4280 9040 4370 9280
rect 4610 9040 4700 9280
rect 4940 9040 5030 9280
rect 5270 9040 5360 9280
rect 5600 9040 5690 9280
rect 5930 9040 6020 9280
rect 6260 9040 6350 9280
rect 6590 9040 6760 9280
rect -5550 8690 6760 9040
rect 8140 21610 20450 21640
rect 8140 21370 8170 21610
rect 8410 21370 8500 21610
rect 8740 21370 8830 21610
rect 9070 21370 9160 21610
rect 9400 21370 9490 21610
rect 9730 21370 9820 21610
rect 10060 21370 10150 21610
rect 10390 21370 10480 21610
rect 10720 21370 10810 21610
rect 11050 21370 11180 21610
rect 11420 21370 11510 21610
rect 11750 21370 11840 21610
rect 12080 21370 12170 21610
rect 12410 21370 12500 21610
rect 12740 21370 12830 21610
rect 13070 21370 13160 21610
rect 13400 21370 13490 21610
rect 13730 21370 13820 21610
rect 14060 21370 14190 21610
rect 14430 21370 14520 21610
rect 14760 21370 14850 21610
rect 15090 21370 15180 21610
rect 15420 21370 15510 21610
rect 15750 21370 15840 21610
rect 16080 21370 16170 21610
rect 16410 21370 16500 21610
rect 16740 21370 16830 21610
rect 17070 21370 17200 21610
rect 17440 21370 17530 21610
rect 17770 21370 17860 21610
rect 18100 21370 18190 21610
rect 18430 21370 18520 21610
rect 18760 21370 18850 21610
rect 19090 21370 19180 21610
rect 19420 21370 19510 21610
rect 19750 21370 19840 21610
rect 20080 21370 20450 21610
rect 8140 20830 20450 21370
rect 8140 20590 8310 20830
rect 8550 20590 8640 20830
rect 8880 20590 8970 20830
rect 9210 20590 9300 20830
rect 9540 20590 9630 20830
rect 9870 20590 9960 20830
rect 10200 20590 10290 20830
rect 10530 20590 10620 20830
rect 10860 20590 10950 20830
rect 11190 20590 11280 20830
rect 11520 20590 11610 20830
rect 11850 20590 11940 20830
rect 12180 20590 12270 20830
rect 12510 20590 12600 20830
rect 12840 20590 12930 20830
rect 13170 20590 13260 20830
rect 13500 20590 13590 20830
rect 13830 20590 13920 20830
rect 14160 20590 14250 20830
rect 14490 20590 14580 20830
rect 14820 20590 14910 20830
rect 15150 20590 15240 20830
rect 15480 20590 15570 20830
rect 15810 20590 15900 20830
rect 16140 20590 16230 20830
rect 16470 20590 16560 20830
rect 16800 20590 16890 20830
rect 17130 20590 17220 20830
rect 17460 20590 17550 20830
rect 17790 20590 17880 20830
rect 18120 20590 18210 20830
rect 18450 20590 18540 20830
rect 18780 20590 18870 20830
rect 19110 20590 19200 20830
rect 19440 20590 19530 20830
rect 19770 20590 19860 20830
rect 20100 20590 20450 20830
rect 8140 20500 20450 20590
rect 8140 20260 8310 20500
rect 8550 20260 8640 20500
rect 8880 20260 8970 20500
rect 9210 20260 9300 20500
rect 9540 20260 9630 20500
rect 9870 20260 9960 20500
rect 10200 20260 10290 20500
rect 10530 20260 10620 20500
rect 10860 20260 10950 20500
rect 11190 20260 11280 20500
rect 11520 20260 11610 20500
rect 11850 20260 11940 20500
rect 12180 20260 12270 20500
rect 12510 20260 12600 20500
rect 12840 20260 12930 20500
rect 13170 20260 13260 20500
rect 13500 20260 13590 20500
rect 13830 20260 13920 20500
rect 14160 20260 14250 20500
rect 14490 20260 14580 20500
rect 14820 20260 14910 20500
rect 15150 20260 15240 20500
rect 15480 20260 15570 20500
rect 15810 20260 15900 20500
rect 16140 20260 16230 20500
rect 16470 20260 16560 20500
rect 16800 20260 16890 20500
rect 17130 20260 17220 20500
rect 17460 20260 17550 20500
rect 17790 20260 17880 20500
rect 18120 20260 18210 20500
rect 18450 20260 18540 20500
rect 18780 20260 18870 20500
rect 19110 20260 19200 20500
rect 19440 20260 19530 20500
rect 19770 20260 19860 20500
rect 20100 20260 20450 20500
rect 8140 20170 20450 20260
rect 8140 19930 8310 20170
rect 8550 19930 8640 20170
rect 8880 19930 8970 20170
rect 9210 19930 9300 20170
rect 9540 19930 9630 20170
rect 9870 19930 9960 20170
rect 10200 19930 10290 20170
rect 10530 19930 10620 20170
rect 10860 19930 10950 20170
rect 11190 19930 11280 20170
rect 11520 19930 11610 20170
rect 11850 19930 11940 20170
rect 12180 19930 12270 20170
rect 12510 19930 12600 20170
rect 12840 19930 12930 20170
rect 13170 19930 13260 20170
rect 13500 19930 13590 20170
rect 13830 19930 13920 20170
rect 14160 19930 14250 20170
rect 14490 19930 14580 20170
rect 14820 19930 14910 20170
rect 15150 19930 15240 20170
rect 15480 19930 15570 20170
rect 15810 19930 15900 20170
rect 16140 19930 16230 20170
rect 16470 19930 16560 20170
rect 16800 19930 16890 20170
rect 17130 19930 17220 20170
rect 17460 19930 17550 20170
rect 17790 19930 17880 20170
rect 18120 19930 18210 20170
rect 18450 19930 18540 20170
rect 18780 19930 18870 20170
rect 19110 19930 19200 20170
rect 19440 19930 19530 20170
rect 19770 19930 19860 20170
rect 20100 19930 20450 20170
rect 8140 19840 20450 19930
rect 8140 19600 8310 19840
rect 8550 19600 8640 19840
rect 8880 19600 8970 19840
rect 9210 19600 9300 19840
rect 9540 19600 9630 19840
rect 9870 19600 9960 19840
rect 10200 19600 10290 19840
rect 10530 19600 10620 19840
rect 10860 19600 10950 19840
rect 11190 19600 11280 19840
rect 11520 19600 11610 19840
rect 11850 19600 11940 19840
rect 12180 19600 12270 19840
rect 12510 19600 12600 19840
rect 12840 19600 12930 19840
rect 13170 19600 13260 19840
rect 13500 19600 13590 19840
rect 13830 19600 13920 19840
rect 14160 19600 14250 19840
rect 14490 19600 14580 19840
rect 14820 19600 14910 19840
rect 15150 19600 15240 19840
rect 15480 19600 15570 19840
rect 15810 19600 15900 19840
rect 16140 19600 16230 19840
rect 16470 19600 16560 19840
rect 16800 19600 16890 19840
rect 17130 19600 17220 19840
rect 17460 19600 17550 19840
rect 17790 19600 17880 19840
rect 18120 19600 18210 19840
rect 18450 19600 18540 19840
rect 18780 19600 18870 19840
rect 19110 19600 19200 19840
rect 19440 19600 19530 19840
rect 19770 19600 19860 19840
rect 20100 19600 20450 19840
rect 8140 19510 20450 19600
rect 8140 19270 8310 19510
rect 8550 19270 8640 19510
rect 8880 19270 8970 19510
rect 9210 19270 9300 19510
rect 9540 19270 9630 19510
rect 9870 19270 9960 19510
rect 10200 19270 10290 19510
rect 10530 19270 10620 19510
rect 10860 19270 10950 19510
rect 11190 19270 11280 19510
rect 11520 19270 11610 19510
rect 11850 19270 11940 19510
rect 12180 19270 12270 19510
rect 12510 19270 12600 19510
rect 12840 19270 12930 19510
rect 13170 19270 13260 19510
rect 13500 19270 13590 19510
rect 13830 19270 13920 19510
rect 14160 19270 14250 19510
rect 14490 19270 14580 19510
rect 14820 19270 14910 19510
rect 15150 19270 15240 19510
rect 15480 19270 15570 19510
rect 15810 19270 15900 19510
rect 16140 19270 16230 19510
rect 16470 19270 16560 19510
rect 16800 19270 16890 19510
rect 17130 19270 17220 19510
rect 17460 19270 17550 19510
rect 17790 19270 17880 19510
rect 18120 19270 18210 19510
rect 18450 19270 18540 19510
rect 18780 19270 18870 19510
rect 19110 19270 19200 19510
rect 19440 19270 19530 19510
rect 19770 19270 19860 19510
rect 20100 19270 20450 19510
rect 8140 19180 20450 19270
rect 8140 18940 8310 19180
rect 8550 18940 8640 19180
rect 8880 18940 8970 19180
rect 9210 18940 9300 19180
rect 9540 18940 9630 19180
rect 9870 18940 9960 19180
rect 10200 18940 10290 19180
rect 10530 18940 10620 19180
rect 10860 18940 10950 19180
rect 11190 18940 11280 19180
rect 11520 18940 11610 19180
rect 11850 18940 11940 19180
rect 12180 18940 12270 19180
rect 12510 18940 12600 19180
rect 12840 18940 12930 19180
rect 13170 18940 13260 19180
rect 13500 18940 13590 19180
rect 13830 18940 13920 19180
rect 14160 18940 14250 19180
rect 14490 18940 14580 19180
rect 14820 18940 14910 19180
rect 15150 18940 15240 19180
rect 15480 18940 15570 19180
rect 15810 18940 15900 19180
rect 16140 18940 16230 19180
rect 16470 18940 16560 19180
rect 16800 18940 16890 19180
rect 17130 18940 17220 19180
rect 17460 18940 17550 19180
rect 17790 18940 17880 19180
rect 18120 18940 18210 19180
rect 18450 18940 18540 19180
rect 18780 18940 18870 19180
rect 19110 18940 19200 19180
rect 19440 18940 19530 19180
rect 19770 18940 19860 19180
rect 20100 18940 20450 19180
rect 8140 18850 20450 18940
rect 8140 18610 8310 18850
rect 8550 18610 8640 18850
rect 8880 18610 8970 18850
rect 9210 18610 9300 18850
rect 9540 18610 9630 18850
rect 9870 18610 9960 18850
rect 10200 18610 10290 18850
rect 10530 18610 10620 18850
rect 10860 18610 10950 18850
rect 11190 18610 11280 18850
rect 11520 18610 11610 18850
rect 11850 18610 11940 18850
rect 12180 18610 12270 18850
rect 12510 18610 12600 18850
rect 12840 18610 12930 18850
rect 13170 18610 13260 18850
rect 13500 18610 13590 18850
rect 13830 18610 13920 18850
rect 14160 18610 14250 18850
rect 14490 18610 14580 18850
rect 14820 18610 14910 18850
rect 15150 18610 15240 18850
rect 15480 18610 15570 18850
rect 15810 18610 15900 18850
rect 16140 18610 16230 18850
rect 16470 18610 16560 18850
rect 16800 18610 16890 18850
rect 17130 18610 17220 18850
rect 17460 18610 17550 18850
rect 17790 18610 17880 18850
rect 18120 18610 18210 18850
rect 18450 18610 18540 18850
rect 18780 18610 18870 18850
rect 19110 18610 19200 18850
rect 19440 18610 19530 18850
rect 19770 18610 19860 18850
rect 20100 18610 20450 18850
rect 8140 18520 20450 18610
rect 8140 18280 8310 18520
rect 8550 18280 8640 18520
rect 8880 18280 8970 18520
rect 9210 18280 9300 18520
rect 9540 18280 9630 18520
rect 9870 18280 9960 18520
rect 10200 18280 10290 18520
rect 10530 18280 10620 18520
rect 10860 18280 10950 18520
rect 11190 18280 11280 18520
rect 11520 18280 11610 18520
rect 11850 18280 11940 18520
rect 12180 18280 12270 18520
rect 12510 18280 12600 18520
rect 12840 18280 12930 18520
rect 13170 18280 13260 18520
rect 13500 18280 13590 18520
rect 13830 18280 13920 18520
rect 14160 18280 14250 18520
rect 14490 18280 14580 18520
rect 14820 18280 14910 18520
rect 15150 18280 15240 18520
rect 15480 18280 15570 18520
rect 15810 18280 15900 18520
rect 16140 18280 16230 18520
rect 16470 18280 16560 18520
rect 16800 18280 16890 18520
rect 17130 18280 17220 18520
rect 17460 18280 17550 18520
rect 17790 18280 17880 18520
rect 18120 18280 18210 18520
rect 18450 18280 18540 18520
rect 18780 18280 18870 18520
rect 19110 18280 19200 18520
rect 19440 18280 19530 18520
rect 19770 18280 19860 18520
rect 20100 18280 20450 18520
rect 8140 18190 20450 18280
rect 8140 17950 8310 18190
rect 8550 17950 8640 18190
rect 8880 17950 8970 18190
rect 9210 17950 9300 18190
rect 9540 17950 9630 18190
rect 9870 17950 9960 18190
rect 10200 17950 10290 18190
rect 10530 17950 10620 18190
rect 10860 17950 10950 18190
rect 11190 17950 11280 18190
rect 11520 17950 11610 18190
rect 11850 17950 11940 18190
rect 12180 17950 12270 18190
rect 12510 17950 12600 18190
rect 12840 17950 12930 18190
rect 13170 17950 13260 18190
rect 13500 17950 13590 18190
rect 13830 17950 13920 18190
rect 14160 17950 14250 18190
rect 14490 17950 14580 18190
rect 14820 17950 14910 18190
rect 15150 17950 15240 18190
rect 15480 17950 15570 18190
rect 15810 17950 15900 18190
rect 16140 17950 16230 18190
rect 16470 17950 16560 18190
rect 16800 17950 16890 18190
rect 17130 17950 17220 18190
rect 17460 17950 17550 18190
rect 17790 17950 17880 18190
rect 18120 17950 18210 18190
rect 18450 17950 18540 18190
rect 18780 17950 18870 18190
rect 19110 17950 19200 18190
rect 19440 17950 19530 18190
rect 19770 17950 19860 18190
rect 20100 17950 20450 18190
rect 8140 17860 20450 17950
rect 8140 17620 8310 17860
rect 8550 17620 8640 17860
rect 8880 17620 8970 17860
rect 9210 17620 9300 17860
rect 9540 17620 9630 17860
rect 9870 17620 9960 17860
rect 10200 17620 10290 17860
rect 10530 17620 10620 17860
rect 10860 17620 10950 17860
rect 11190 17620 11280 17860
rect 11520 17620 11610 17860
rect 11850 17620 11940 17860
rect 12180 17620 12270 17860
rect 12510 17620 12600 17860
rect 12840 17620 12930 17860
rect 13170 17620 13260 17860
rect 13500 17620 13590 17860
rect 13830 17620 13920 17860
rect 14160 17620 14250 17860
rect 14490 17620 14580 17860
rect 14820 17620 14910 17860
rect 15150 17620 15240 17860
rect 15480 17620 15570 17860
rect 15810 17620 15900 17860
rect 16140 17620 16230 17860
rect 16470 17620 16560 17860
rect 16800 17620 16890 17860
rect 17130 17620 17220 17860
rect 17460 17620 17550 17860
rect 17790 17620 17880 17860
rect 18120 17620 18210 17860
rect 18450 17620 18540 17860
rect 18780 17620 18870 17860
rect 19110 17620 19200 17860
rect 19440 17620 19530 17860
rect 19770 17620 19860 17860
rect 20100 17620 20450 17860
rect 8140 17530 20450 17620
rect 8140 17290 8310 17530
rect 8550 17290 8640 17530
rect 8880 17290 8970 17530
rect 9210 17290 9300 17530
rect 9540 17290 9630 17530
rect 9870 17290 9960 17530
rect 10200 17290 10290 17530
rect 10530 17290 10620 17530
rect 10860 17290 10950 17530
rect 11190 17290 11280 17530
rect 11520 17290 11610 17530
rect 11850 17290 11940 17530
rect 12180 17290 12270 17530
rect 12510 17290 12600 17530
rect 12840 17290 12930 17530
rect 13170 17290 13260 17530
rect 13500 17290 13590 17530
rect 13830 17290 13920 17530
rect 14160 17290 14250 17530
rect 14490 17290 14580 17530
rect 14820 17290 14910 17530
rect 15150 17290 15240 17530
rect 15480 17290 15570 17530
rect 15810 17290 15900 17530
rect 16140 17290 16230 17530
rect 16470 17290 16560 17530
rect 16800 17290 16890 17530
rect 17130 17290 17220 17530
rect 17460 17290 17550 17530
rect 17790 17290 17880 17530
rect 18120 17290 18210 17530
rect 18450 17290 18540 17530
rect 18780 17290 18870 17530
rect 19110 17290 19200 17530
rect 19440 17290 19530 17530
rect 19770 17290 19860 17530
rect 20100 17290 20450 17530
rect 8140 17200 20450 17290
rect 8140 16960 8310 17200
rect 8550 16960 8640 17200
rect 8880 16960 8970 17200
rect 9210 16960 9300 17200
rect 9540 16960 9630 17200
rect 9870 16960 9960 17200
rect 10200 16960 10290 17200
rect 10530 16960 10620 17200
rect 10860 16960 10950 17200
rect 11190 16960 11280 17200
rect 11520 16960 11610 17200
rect 11850 16960 11940 17200
rect 12180 16960 12270 17200
rect 12510 16960 12600 17200
rect 12840 16960 12930 17200
rect 13170 16960 13260 17200
rect 13500 16960 13590 17200
rect 13830 16960 13920 17200
rect 14160 16960 14250 17200
rect 14490 16960 14580 17200
rect 14820 16960 14910 17200
rect 15150 16960 15240 17200
rect 15480 16960 15570 17200
rect 15810 16960 15900 17200
rect 16140 16960 16230 17200
rect 16470 16960 16560 17200
rect 16800 16960 16890 17200
rect 17130 16960 17220 17200
rect 17460 16960 17550 17200
rect 17790 16960 17880 17200
rect 18120 16960 18210 17200
rect 18450 16960 18540 17200
rect 18780 16960 18870 17200
rect 19110 16960 19200 17200
rect 19440 16960 19530 17200
rect 19770 16960 19860 17200
rect 20100 16960 20450 17200
rect 8140 16870 20450 16960
rect 8140 16630 8310 16870
rect 8550 16630 8640 16870
rect 8880 16630 8970 16870
rect 9210 16630 9300 16870
rect 9540 16630 9630 16870
rect 9870 16630 9960 16870
rect 10200 16630 10290 16870
rect 10530 16630 10620 16870
rect 10860 16630 10950 16870
rect 11190 16630 11280 16870
rect 11520 16630 11610 16870
rect 11850 16630 11940 16870
rect 12180 16630 12270 16870
rect 12510 16630 12600 16870
rect 12840 16630 12930 16870
rect 13170 16630 13260 16870
rect 13500 16630 13590 16870
rect 13830 16630 13920 16870
rect 14160 16630 14250 16870
rect 14490 16630 14580 16870
rect 14820 16630 14910 16870
rect 15150 16630 15240 16870
rect 15480 16630 15570 16870
rect 15810 16630 15900 16870
rect 16140 16630 16230 16870
rect 16470 16630 16560 16870
rect 16800 16630 16890 16870
rect 17130 16630 17220 16870
rect 17460 16630 17550 16870
rect 17790 16630 17880 16870
rect 18120 16630 18210 16870
rect 18450 16630 18540 16870
rect 18780 16630 18870 16870
rect 19110 16630 19200 16870
rect 19440 16630 19530 16870
rect 19770 16630 19860 16870
rect 20100 16630 20450 16870
rect 8140 16540 20450 16630
rect 8140 16300 8310 16540
rect 8550 16300 8640 16540
rect 8880 16300 8970 16540
rect 9210 16300 9300 16540
rect 9540 16300 9630 16540
rect 9870 16300 9960 16540
rect 10200 16300 10290 16540
rect 10530 16300 10620 16540
rect 10860 16300 10950 16540
rect 11190 16300 11280 16540
rect 11520 16300 11610 16540
rect 11850 16300 11940 16540
rect 12180 16300 12270 16540
rect 12510 16300 12600 16540
rect 12840 16300 12930 16540
rect 13170 16300 13260 16540
rect 13500 16300 13590 16540
rect 13830 16300 13920 16540
rect 14160 16300 14250 16540
rect 14490 16300 14580 16540
rect 14820 16300 14910 16540
rect 15150 16300 15240 16540
rect 15480 16300 15570 16540
rect 15810 16300 15900 16540
rect 16140 16300 16230 16540
rect 16470 16300 16560 16540
rect 16800 16300 16890 16540
rect 17130 16300 17220 16540
rect 17460 16300 17550 16540
rect 17790 16300 17880 16540
rect 18120 16300 18210 16540
rect 18450 16300 18540 16540
rect 18780 16300 18870 16540
rect 19110 16300 19200 16540
rect 19440 16300 19530 16540
rect 19770 16300 19860 16540
rect 20100 16300 20450 16540
rect 8140 16210 20450 16300
rect 8140 15970 8310 16210
rect 8550 15970 8640 16210
rect 8880 15970 8970 16210
rect 9210 15970 9300 16210
rect 9540 15970 9630 16210
rect 9870 15970 9960 16210
rect 10200 15970 10290 16210
rect 10530 15970 10620 16210
rect 10860 15970 10950 16210
rect 11190 15970 11280 16210
rect 11520 15970 11610 16210
rect 11850 15970 11940 16210
rect 12180 15970 12270 16210
rect 12510 15970 12600 16210
rect 12840 15970 12930 16210
rect 13170 15970 13260 16210
rect 13500 15970 13590 16210
rect 13830 15970 13920 16210
rect 14160 15970 14250 16210
rect 14490 15970 14580 16210
rect 14820 15970 14910 16210
rect 15150 15970 15240 16210
rect 15480 15970 15570 16210
rect 15810 15970 15900 16210
rect 16140 15970 16230 16210
rect 16470 15970 16560 16210
rect 16800 15970 16890 16210
rect 17130 15970 17220 16210
rect 17460 15970 17550 16210
rect 17790 15970 17880 16210
rect 18120 15970 18210 16210
rect 18450 15970 18540 16210
rect 18780 15970 18870 16210
rect 19110 15970 19200 16210
rect 19440 15970 19530 16210
rect 19770 15970 19860 16210
rect 20100 15970 20450 16210
rect 8140 15880 20450 15970
rect 8140 15640 8310 15880
rect 8550 15640 8640 15880
rect 8880 15640 8970 15880
rect 9210 15640 9300 15880
rect 9540 15640 9630 15880
rect 9870 15640 9960 15880
rect 10200 15640 10290 15880
rect 10530 15640 10620 15880
rect 10860 15640 10950 15880
rect 11190 15640 11280 15880
rect 11520 15640 11610 15880
rect 11850 15640 11940 15880
rect 12180 15640 12270 15880
rect 12510 15640 12600 15880
rect 12840 15640 12930 15880
rect 13170 15640 13260 15880
rect 13500 15640 13590 15880
rect 13830 15640 13920 15880
rect 14160 15640 14250 15880
rect 14490 15640 14580 15880
rect 14820 15640 14910 15880
rect 15150 15640 15240 15880
rect 15480 15640 15570 15880
rect 15810 15640 15900 15880
rect 16140 15640 16230 15880
rect 16470 15640 16560 15880
rect 16800 15640 16890 15880
rect 17130 15640 17220 15880
rect 17460 15640 17550 15880
rect 17790 15640 17880 15880
rect 18120 15640 18210 15880
rect 18450 15640 18540 15880
rect 18780 15640 18870 15880
rect 19110 15640 19200 15880
rect 19440 15640 19530 15880
rect 19770 15640 19860 15880
rect 20100 15640 20450 15880
rect 8140 15550 20450 15640
rect 8140 15310 8310 15550
rect 8550 15310 8640 15550
rect 8880 15310 8970 15550
rect 9210 15310 9300 15550
rect 9540 15310 9630 15550
rect 9870 15310 9960 15550
rect 10200 15310 10290 15550
rect 10530 15310 10620 15550
rect 10860 15310 10950 15550
rect 11190 15310 11280 15550
rect 11520 15310 11610 15550
rect 11850 15310 11940 15550
rect 12180 15310 12270 15550
rect 12510 15310 12600 15550
rect 12840 15310 12930 15550
rect 13170 15310 13260 15550
rect 13500 15310 13590 15550
rect 13830 15310 13920 15550
rect 14160 15310 14250 15550
rect 14490 15310 14580 15550
rect 14820 15310 14910 15550
rect 15150 15310 15240 15550
rect 15480 15310 15570 15550
rect 15810 15310 15900 15550
rect 16140 15310 16230 15550
rect 16470 15310 16560 15550
rect 16800 15310 16890 15550
rect 17130 15310 17220 15550
rect 17460 15310 17550 15550
rect 17790 15310 17880 15550
rect 18120 15310 18210 15550
rect 18450 15310 18540 15550
rect 18780 15310 18870 15550
rect 19110 15310 19200 15550
rect 19440 15310 19530 15550
rect 19770 15310 19860 15550
rect 20100 15310 20450 15550
rect 8140 15220 20450 15310
rect 8140 14980 8310 15220
rect 8550 14980 8640 15220
rect 8880 14980 8970 15220
rect 9210 14980 9300 15220
rect 9540 14980 9630 15220
rect 9870 14980 9960 15220
rect 10200 14980 10290 15220
rect 10530 14980 10620 15220
rect 10860 14980 10950 15220
rect 11190 14980 11280 15220
rect 11520 14980 11610 15220
rect 11850 14980 11940 15220
rect 12180 14980 12270 15220
rect 12510 14980 12600 15220
rect 12840 14980 12930 15220
rect 13170 14980 13260 15220
rect 13500 14980 13590 15220
rect 13830 14980 13920 15220
rect 14160 14980 14250 15220
rect 14490 14980 14580 15220
rect 14820 14980 14910 15220
rect 15150 14980 15240 15220
rect 15480 14980 15570 15220
rect 15810 14980 15900 15220
rect 16140 14980 16230 15220
rect 16470 14980 16560 15220
rect 16800 14980 16890 15220
rect 17130 14980 17220 15220
rect 17460 14980 17550 15220
rect 17790 14980 17880 15220
rect 18120 14980 18210 15220
rect 18450 14980 18540 15220
rect 18780 14980 18870 15220
rect 19110 14980 19200 15220
rect 19440 14980 19530 15220
rect 19770 14980 19860 15220
rect 20100 14980 20450 15220
rect 8140 14890 20450 14980
rect 8140 14650 8310 14890
rect 8550 14650 8640 14890
rect 8880 14650 8970 14890
rect 9210 14650 9300 14890
rect 9540 14650 9630 14890
rect 9870 14650 9960 14890
rect 10200 14650 10290 14890
rect 10530 14650 10620 14890
rect 10860 14650 10950 14890
rect 11190 14650 11280 14890
rect 11520 14650 11610 14890
rect 11850 14650 11940 14890
rect 12180 14650 12270 14890
rect 12510 14650 12600 14890
rect 12840 14650 12930 14890
rect 13170 14650 13260 14890
rect 13500 14650 13590 14890
rect 13830 14650 13920 14890
rect 14160 14650 14250 14890
rect 14490 14650 14580 14890
rect 14820 14650 14910 14890
rect 15150 14650 15240 14890
rect 15480 14650 15570 14890
rect 15810 14650 15900 14890
rect 16140 14650 16230 14890
rect 16470 14650 16560 14890
rect 16800 14650 16890 14890
rect 17130 14650 17220 14890
rect 17460 14650 17550 14890
rect 17790 14650 17880 14890
rect 18120 14650 18210 14890
rect 18450 14650 18540 14890
rect 18780 14650 18870 14890
rect 19110 14650 19200 14890
rect 19440 14650 19530 14890
rect 19770 14650 19860 14890
rect 20100 14650 20450 14890
rect 8140 14560 20450 14650
rect 8140 14320 8310 14560
rect 8550 14320 8640 14560
rect 8880 14320 8970 14560
rect 9210 14320 9300 14560
rect 9540 14320 9630 14560
rect 9870 14320 9960 14560
rect 10200 14320 10290 14560
rect 10530 14320 10620 14560
rect 10860 14320 10950 14560
rect 11190 14320 11280 14560
rect 11520 14320 11610 14560
rect 11850 14320 11940 14560
rect 12180 14320 12270 14560
rect 12510 14320 12600 14560
rect 12840 14320 12930 14560
rect 13170 14320 13260 14560
rect 13500 14320 13590 14560
rect 13830 14320 13920 14560
rect 14160 14320 14250 14560
rect 14490 14320 14580 14560
rect 14820 14320 14910 14560
rect 15150 14320 15240 14560
rect 15480 14320 15570 14560
rect 15810 14320 15900 14560
rect 16140 14320 16230 14560
rect 16470 14320 16560 14560
rect 16800 14320 16890 14560
rect 17130 14320 17220 14560
rect 17460 14320 17550 14560
rect 17790 14320 17880 14560
rect 18120 14320 18210 14560
rect 18450 14320 18540 14560
rect 18780 14320 18870 14560
rect 19110 14320 19200 14560
rect 19440 14320 19530 14560
rect 19770 14320 19860 14560
rect 20100 14320 20450 14560
rect 8140 14230 20450 14320
rect 8140 13990 8310 14230
rect 8550 13990 8640 14230
rect 8880 13990 8970 14230
rect 9210 13990 9300 14230
rect 9540 13990 9630 14230
rect 9870 13990 9960 14230
rect 10200 13990 10290 14230
rect 10530 13990 10620 14230
rect 10860 13990 10950 14230
rect 11190 13990 11280 14230
rect 11520 13990 11610 14230
rect 11850 13990 11940 14230
rect 12180 13990 12270 14230
rect 12510 13990 12600 14230
rect 12840 13990 12930 14230
rect 13170 13990 13260 14230
rect 13500 13990 13590 14230
rect 13830 13990 13920 14230
rect 14160 13990 14250 14230
rect 14490 13990 14580 14230
rect 14820 13990 14910 14230
rect 15150 13990 15240 14230
rect 15480 13990 15570 14230
rect 15810 13990 15900 14230
rect 16140 13990 16230 14230
rect 16470 13990 16560 14230
rect 16800 13990 16890 14230
rect 17130 13990 17220 14230
rect 17460 13990 17550 14230
rect 17790 13990 17880 14230
rect 18120 13990 18210 14230
rect 18450 13990 18540 14230
rect 18780 13990 18870 14230
rect 19110 13990 19200 14230
rect 19440 13990 19530 14230
rect 19770 13990 19860 14230
rect 20100 13990 20450 14230
rect 8140 13900 20450 13990
rect 8140 13660 8310 13900
rect 8550 13660 8640 13900
rect 8880 13660 8970 13900
rect 9210 13660 9300 13900
rect 9540 13660 9630 13900
rect 9870 13660 9960 13900
rect 10200 13660 10290 13900
rect 10530 13660 10620 13900
rect 10860 13660 10950 13900
rect 11190 13660 11280 13900
rect 11520 13660 11610 13900
rect 11850 13660 11940 13900
rect 12180 13660 12270 13900
rect 12510 13660 12600 13900
rect 12840 13660 12930 13900
rect 13170 13660 13260 13900
rect 13500 13660 13590 13900
rect 13830 13660 13920 13900
rect 14160 13660 14250 13900
rect 14490 13660 14580 13900
rect 14820 13660 14910 13900
rect 15150 13660 15240 13900
rect 15480 13660 15570 13900
rect 15810 13660 15900 13900
rect 16140 13660 16230 13900
rect 16470 13660 16560 13900
rect 16800 13660 16890 13900
rect 17130 13660 17220 13900
rect 17460 13660 17550 13900
rect 17790 13660 17880 13900
rect 18120 13660 18210 13900
rect 18450 13660 18540 13900
rect 18780 13660 18870 13900
rect 19110 13660 19200 13900
rect 19440 13660 19530 13900
rect 19770 13660 19860 13900
rect 20100 13660 20450 13900
rect 8140 13570 20450 13660
rect 8140 13330 8310 13570
rect 8550 13330 8640 13570
rect 8880 13330 8970 13570
rect 9210 13330 9300 13570
rect 9540 13330 9630 13570
rect 9870 13330 9960 13570
rect 10200 13330 10290 13570
rect 10530 13330 10620 13570
rect 10860 13330 10950 13570
rect 11190 13330 11280 13570
rect 11520 13330 11610 13570
rect 11850 13330 11940 13570
rect 12180 13330 12270 13570
rect 12510 13330 12600 13570
rect 12840 13330 12930 13570
rect 13170 13330 13260 13570
rect 13500 13330 13590 13570
rect 13830 13330 13920 13570
rect 14160 13330 14250 13570
rect 14490 13330 14580 13570
rect 14820 13330 14910 13570
rect 15150 13330 15240 13570
rect 15480 13330 15570 13570
rect 15810 13330 15900 13570
rect 16140 13330 16230 13570
rect 16470 13330 16560 13570
rect 16800 13330 16890 13570
rect 17130 13330 17220 13570
rect 17460 13330 17550 13570
rect 17790 13330 17880 13570
rect 18120 13330 18210 13570
rect 18450 13330 18540 13570
rect 18780 13330 18870 13570
rect 19110 13330 19200 13570
rect 19440 13330 19530 13570
rect 19770 13330 19860 13570
rect 20100 13330 20450 13570
rect 8140 13240 20450 13330
rect 8140 13000 8310 13240
rect 8550 13000 8640 13240
rect 8880 13000 8970 13240
rect 9210 13000 9300 13240
rect 9540 13000 9630 13240
rect 9870 13000 9960 13240
rect 10200 13000 10290 13240
rect 10530 13000 10620 13240
rect 10860 13000 10950 13240
rect 11190 13000 11280 13240
rect 11520 13000 11610 13240
rect 11850 13000 11940 13240
rect 12180 13000 12270 13240
rect 12510 13000 12600 13240
rect 12840 13000 12930 13240
rect 13170 13000 13260 13240
rect 13500 13000 13590 13240
rect 13830 13000 13920 13240
rect 14160 13000 14250 13240
rect 14490 13000 14580 13240
rect 14820 13000 14910 13240
rect 15150 13000 15240 13240
rect 15480 13000 15570 13240
rect 15810 13000 15900 13240
rect 16140 13000 16230 13240
rect 16470 13000 16560 13240
rect 16800 13000 16890 13240
rect 17130 13000 17220 13240
rect 17460 13000 17550 13240
rect 17790 13000 17880 13240
rect 18120 13000 18210 13240
rect 18450 13000 18540 13240
rect 18780 13000 18870 13240
rect 19110 13000 19200 13240
rect 19440 13000 19530 13240
rect 19770 13000 19860 13240
rect 20100 13000 20450 13240
rect 8140 12910 20450 13000
rect 8140 12670 8310 12910
rect 8550 12670 8640 12910
rect 8880 12670 8970 12910
rect 9210 12670 9300 12910
rect 9540 12670 9630 12910
rect 9870 12670 9960 12910
rect 10200 12670 10290 12910
rect 10530 12670 10620 12910
rect 10860 12670 10950 12910
rect 11190 12670 11280 12910
rect 11520 12670 11610 12910
rect 11850 12670 11940 12910
rect 12180 12670 12270 12910
rect 12510 12670 12600 12910
rect 12840 12670 12930 12910
rect 13170 12670 13260 12910
rect 13500 12670 13590 12910
rect 13830 12670 13920 12910
rect 14160 12670 14250 12910
rect 14490 12670 14580 12910
rect 14820 12670 14910 12910
rect 15150 12670 15240 12910
rect 15480 12670 15570 12910
rect 15810 12670 15900 12910
rect 16140 12670 16230 12910
rect 16470 12670 16560 12910
rect 16800 12670 16890 12910
rect 17130 12670 17220 12910
rect 17460 12670 17550 12910
rect 17790 12670 17880 12910
rect 18120 12670 18210 12910
rect 18450 12670 18540 12910
rect 18780 12670 18870 12910
rect 19110 12670 19200 12910
rect 19440 12670 19530 12910
rect 19770 12670 19860 12910
rect 20100 12670 20450 12910
rect 8140 12580 20450 12670
rect 8140 12340 8310 12580
rect 8550 12340 8640 12580
rect 8880 12340 8970 12580
rect 9210 12340 9300 12580
rect 9540 12340 9630 12580
rect 9870 12340 9960 12580
rect 10200 12340 10290 12580
rect 10530 12340 10620 12580
rect 10860 12340 10950 12580
rect 11190 12340 11280 12580
rect 11520 12340 11610 12580
rect 11850 12340 11940 12580
rect 12180 12340 12270 12580
rect 12510 12340 12600 12580
rect 12840 12340 12930 12580
rect 13170 12340 13260 12580
rect 13500 12340 13590 12580
rect 13830 12340 13920 12580
rect 14160 12340 14250 12580
rect 14490 12340 14580 12580
rect 14820 12340 14910 12580
rect 15150 12340 15240 12580
rect 15480 12340 15570 12580
rect 15810 12340 15900 12580
rect 16140 12340 16230 12580
rect 16470 12340 16560 12580
rect 16800 12340 16890 12580
rect 17130 12340 17220 12580
rect 17460 12340 17550 12580
rect 17790 12340 17880 12580
rect 18120 12340 18210 12580
rect 18450 12340 18540 12580
rect 18780 12340 18870 12580
rect 19110 12340 19200 12580
rect 19440 12340 19530 12580
rect 19770 12340 19860 12580
rect 20100 12340 20450 12580
rect 8140 12250 20450 12340
rect 8140 12010 8310 12250
rect 8550 12010 8640 12250
rect 8880 12010 8970 12250
rect 9210 12010 9300 12250
rect 9540 12010 9630 12250
rect 9870 12010 9960 12250
rect 10200 12010 10290 12250
rect 10530 12010 10620 12250
rect 10860 12010 10950 12250
rect 11190 12010 11280 12250
rect 11520 12010 11610 12250
rect 11850 12010 11940 12250
rect 12180 12010 12270 12250
rect 12510 12010 12600 12250
rect 12840 12010 12930 12250
rect 13170 12010 13260 12250
rect 13500 12010 13590 12250
rect 13830 12010 13920 12250
rect 14160 12010 14250 12250
rect 14490 12010 14580 12250
rect 14820 12010 14910 12250
rect 15150 12010 15240 12250
rect 15480 12010 15570 12250
rect 15810 12010 15900 12250
rect 16140 12010 16230 12250
rect 16470 12010 16560 12250
rect 16800 12010 16890 12250
rect 17130 12010 17220 12250
rect 17460 12010 17550 12250
rect 17790 12010 17880 12250
rect 18120 12010 18210 12250
rect 18450 12010 18540 12250
rect 18780 12010 18870 12250
rect 19110 12010 19200 12250
rect 19440 12010 19530 12250
rect 19770 12010 19860 12250
rect 20100 12010 20450 12250
rect 8140 11920 20450 12010
rect 8140 11680 8310 11920
rect 8550 11680 8640 11920
rect 8880 11680 8970 11920
rect 9210 11680 9300 11920
rect 9540 11680 9630 11920
rect 9870 11680 9960 11920
rect 10200 11680 10290 11920
rect 10530 11680 10620 11920
rect 10860 11680 10950 11920
rect 11190 11680 11280 11920
rect 11520 11680 11610 11920
rect 11850 11680 11940 11920
rect 12180 11680 12270 11920
rect 12510 11680 12600 11920
rect 12840 11680 12930 11920
rect 13170 11680 13260 11920
rect 13500 11680 13590 11920
rect 13830 11680 13920 11920
rect 14160 11680 14250 11920
rect 14490 11680 14580 11920
rect 14820 11680 14910 11920
rect 15150 11680 15240 11920
rect 15480 11680 15570 11920
rect 15810 11680 15900 11920
rect 16140 11680 16230 11920
rect 16470 11680 16560 11920
rect 16800 11680 16890 11920
rect 17130 11680 17220 11920
rect 17460 11680 17550 11920
rect 17790 11680 17880 11920
rect 18120 11680 18210 11920
rect 18450 11680 18540 11920
rect 18780 11680 18870 11920
rect 19110 11680 19200 11920
rect 19440 11680 19530 11920
rect 19770 11680 19860 11920
rect 20100 11680 20450 11920
rect 8140 11590 20450 11680
rect 8140 11350 8310 11590
rect 8550 11350 8640 11590
rect 8880 11350 8970 11590
rect 9210 11350 9300 11590
rect 9540 11350 9630 11590
rect 9870 11350 9960 11590
rect 10200 11350 10290 11590
rect 10530 11350 10620 11590
rect 10860 11350 10950 11590
rect 11190 11350 11280 11590
rect 11520 11350 11610 11590
rect 11850 11350 11940 11590
rect 12180 11350 12270 11590
rect 12510 11350 12600 11590
rect 12840 11350 12930 11590
rect 13170 11350 13260 11590
rect 13500 11350 13590 11590
rect 13830 11350 13920 11590
rect 14160 11350 14250 11590
rect 14490 11350 14580 11590
rect 14820 11350 14910 11590
rect 15150 11350 15240 11590
rect 15480 11350 15570 11590
rect 15810 11350 15900 11590
rect 16140 11350 16230 11590
rect 16470 11350 16560 11590
rect 16800 11350 16890 11590
rect 17130 11350 17220 11590
rect 17460 11350 17550 11590
rect 17790 11350 17880 11590
rect 18120 11350 18210 11590
rect 18450 11350 18540 11590
rect 18780 11350 18870 11590
rect 19110 11350 19200 11590
rect 19440 11350 19530 11590
rect 19770 11350 19860 11590
rect 20100 11350 20450 11590
rect 8140 11260 20450 11350
rect 8140 11020 8310 11260
rect 8550 11020 8640 11260
rect 8880 11020 8970 11260
rect 9210 11020 9300 11260
rect 9540 11020 9630 11260
rect 9870 11020 9960 11260
rect 10200 11020 10290 11260
rect 10530 11020 10620 11260
rect 10860 11020 10950 11260
rect 11190 11020 11280 11260
rect 11520 11020 11610 11260
rect 11850 11020 11940 11260
rect 12180 11020 12270 11260
rect 12510 11020 12600 11260
rect 12840 11020 12930 11260
rect 13170 11020 13260 11260
rect 13500 11020 13590 11260
rect 13830 11020 13920 11260
rect 14160 11020 14250 11260
rect 14490 11020 14580 11260
rect 14820 11020 14910 11260
rect 15150 11020 15240 11260
rect 15480 11020 15570 11260
rect 15810 11020 15900 11260
rect 16140 11020 16230 11260
rect 16470 11020 16560 11260
rect 16800 11020 16890 11260
rect 17130 11020 17220 11260
rect 17460 11020 17550 11260
rect 17790 11020 17880 11260
rect 18120 11020 18210 11260
rect 18450 11020 18540 11260
rect 18780 11020 18870 11260
rect 19110 11020 19200 11260
rect 19440 11020 19530 11260
rect 19770 11020 19860 11260
rect 20100 11020 20450 11260
rect 8140 10930 20450 11020
rect 8140 10690 8310 10930
rect 8550 10690 8640 10930
rect 8880 10690 8970 10930
rect 9210 10690 9300 10930
rect 9540 10690 9630 10930
rect 9870 10690 9960 10930
rect 10200 10690 10290 10930
rect 10530 10690 10620 10930
rect 10860 10690 10950 10930
rect 11190 10690 11280 10930
rect 11520 10690 11610 10930
rect 11850 10690 11940 10930
rect 12180 10690 12270 10930
rect 12510 10690 12600 10930
rect 12840 10690 12930 10930
rect 13170 10690 13260 10930
rect 13500 10690 13590 10930
rect 13830 10690 13920 10930
rect 14160 10690 14250 10930
rect 14490 10690 14580 10930
rect 14820 10690 14910 10930
rect 15150 10690 15240 10930
rect 15480 10690 15570 10930
rect 15810 10690 15900 10930
rect 16140 10690 16230 10930
rect 16470 10690 16560 10930
rect 16800 10690 16890 10930
rect 17130 10690 17220 10930
rect 17460 10690 17550 10930
rect 17790 10690 17880 10930
rect 18120 10690 18210 10930
rect 18450 10690 18540 10930
rect 18780 10690 18870 10930
rect 19110 10690 19200 10930
rect 19440 10690 19530 10930
rect 19770 10690 19860 10930
rect 20100 10690 20450 10930
rect 8140 10600 20450 10690
rect 8140 10360 8310 10600
rect 8550 10360 8640 10600
rect 8880 10360 8970 10600
rect 9210 10360 9300 10600
rect 9540 10360 9630 10600
rect 9870 10360 9960 10600
rect 10200 10360 10290 10600
rect 10530 10360 10620 10600
rect 10860 10360 10950 10600
rect 11190 10360 11280 10600
rect 11520 10360 11610 10600
rect 11850 10360 11940 10600
rect 12180 10360 12270 10600
rect 12510 10360 12600 10600
rect 12840 10360 12930 10600
rect 13170 10360 13260 10600
rect 13500 10360 13590 10600
rect 13830 10360 13920 10600
rect 14160 10360 14250 10600
rect 14490 10360 14580 10600
rect 14820 10360 14910 10600
rect 15150 10360 15240 10600
rect 15480 10360 15570 10600
rect 15810 10360 15900 10600
rect 16140 10360 16230 10600
rect 16470 10360 16560 10600
rect 16800 10360 16890 10600
rect 17130 10360 17220 10600
rect 17460 10360 17550 10600
rect 17790 10360 17880 10600
rect 18120 10360 18210 10600
rect 18450 10360 18540 10600
rect 18780 10360 18870 10600
rect 19110 10360 19200 10600
rect 19440 10360 19530 10600
rect 19770 10360 19860 10600
rect 20100 10360 20450 10600
rect 8140 10270 20450 10360
rect 8140 10030 8310 10270
rect 8550 10030 8640 10270
rect 8880 10030 8970 10270
rect 9210 10030 9300 10270
rect 9540 10030 9630 10270
rect 9870 10030 9960 10270
rect 10200 10030 10290 10270
rect 10530 10030 10620 10270
rect 10860 10030 10950 10270
rect 11190 10030 11280 10270
rect 11520 10030 11610 10270
rect 11850 10030 11940 10270
rect 12180 10030 12270 10270
rect 12510 10030 12600 10270
rect 12840 10030 12930 10270
rect 13170 10030 13260 10270
rect 13500 10030 13590 10270
rect 13830 10030 13920 10270
rect 14160 10030 14250 10270
rect 14490 10030 14580 10270
rect 14820 10030 14910 10270
rect 15150 10030 15240 10270
rect 15480 10030 15570 10270
rect 15810 10030 15900 10270
rect 16140 10030 16230 10270
rect 16470 10030 16560 10270
rect 16800 10030 16890 10270
rect 17130 10030 17220 10270
rect 17460 10030 17550 10270
rect 17790 10030 17880 10270
rect 18120 10030 18210 10270
rect 18450 10030 18540 10270
rect 18780 10030 18870 10270
rect 19110 10030 19200 10270
rect 19440 10030 19530 10270
rect 19770 10030 19860 10270
rect 20100 10030 20450 10270
rect 8140 9940 20450 10030
rect 8140 9700 8310 9940
rect 8550 9700 8640 9940
rect 8880 9700 8970 9940
rect 9210 9700 9300 9940
rect 9540 9700 9630 9940
rect 9870 9700 9960 9940
rect 10200 9700 10290 9940
rect 10530 9700 10620 9940
rect 10860 9700 10950 9940
rect 11190 9700 11280 9940
rect 11520 9700 11610 9940
rect 11850 9700 11940 9940
rect 12180 9700 12270 9940
rect 12510 9700 12600 9940
rect 12840 9700 12930 9940
rect 13170 9700 13260 9940
rect 13500 9700 13590 9940
rect 13830 9700 13920 9940
rect 14160 9700 14250 9940
rect 14490 9700 14580 9940
rect 14820 9700 14910 9940
rect 15150 9700 15240 9940
rect 15480 9700 15570 9940
rect 15810 9700 15900 9940
rect 16140 9700 16230 9940
rect 16470 9700 16560 9940
rect 16800 9700 16890 9940
rect 17130 9700 17220 9940
rect 17460 9700 17550 9940
rect 17790 9700 17880 9940
rect 18120 9700 18210 9940
rect 18450 9700 18540 9940
rect 18780 9700 18870 9940
rect 19110 9700 19200 9940
rect 19440 9700 19530 9940
rect 19770 9700 19860 9940
rect 20100 9700 20450 9940
rect 8140 9610 20450 9700
rect 8140 9370 8310 9610
rect 8550 9370 8640 9610
rect 8880 9370 8970 9610
rect 9210 9370 9300 9610
rect 9540 9370 9630 9610
rect 9870 9370 9960 9610
rect 10200 9370 10290 9610
rect 10530 9370 10620 9610
rect 10860 9370 10950 9610
rect 11190 9370 11280 9610
rect 11520 9370 11610 9610
rect 11850 9370 11940 9610
rect 12180 9370 12270 9610
rect 12510 9370 12600 9610
rect 12840 9370 12930 9610
rect 13170 9370 13260 9610
rect 13500 9370 13590 9610
rect 13830 9370 13920 9610
rect 14160 9370 14250 9610
rect 14490 9370 14580 9610
rect 14820 9370 14910 9610
rect 15150 9370 15240 9610
rect 15480 9370 15570 9610
rect 15810 9370 15900 9610
rect 16140 9370 16230 9610
rect 16470 9370 16560 9610
rect 16800 9370 16890 9610
rect 17130 9370 17220 9610
rect 17460 9370 17550 9610
rect 17790 9370 17880 9610
rect 18120 9370 18210 9610
rect 18450 9370 18540 9610
rect 18780 9370 18870 9610
rect 19110 9370 19200 9610
rect 19440 9370 19530 9610
rect 19770 9370 19860 9610
rect 20100 9370 20450 9610
rect 8140 9280 20450 9370
rect 8140 9040 8310 9280
rect 8550 9040 8640 9280
rect 8880 9040 8970 9280
rect 9210 9040 9300 9280
rect 9540 9040 9630 9280
rect 9870 9040 9960 9280
rect 10200 9040 10290 9280
rect 10530 9040 10620 9280
rect 10860 9040 10950 9280
rect 11190 9040 11280 9280
rect 11520 9040 11610 9280
rect 11850 9040 11940 9280
rect 12180 9040 12270 9280
rect 12510 9040 12600 9280
rect 12840 9040 12930 9280
rect 13170 9040 13260 9280
rect 13500 9040 13590 9280
rect 13830 9040 13920 9280
rect 14160 9040 14250 9280
rect 14490 9040 14580 9280
rect 14820 9040 14910 9280
rect 15150 9040 15240 9280
rect 15480 9040 15570 9280
rect 15810 9040 15900 9280
rect 16140 9040 16230 9280
rect 16470 9040 16560 9280
rect 16800 9040 16890 9280
rect 17130 9040 17220 9280
rect 17460 9040 17550 9280
rect 17790 9040 17880 9280
rect 18120 9040 18210 9280
rect 18450 9040 18540 9280
rect 18780 9040 18870 9280
rect 19110 9040 19200 9280
rect 19440 9040 19530 9280
rect 19770 9040 19860 9280
rect 20100 9040 20450 9280
rect 8140 8690 20450 9040
rect -6530 7270 29270 8130
rect -6530 7100 23510 7270
rect -6530 -2160 -2830 7100
rect 1540 6910 3140 7100
rect 1540 6670 1720 6910
rect 1960 6670 2050 6910
rect 2290 6670 2390 6910
rect 2630 6670 2720 6910
rect 2960 6670 3140 6910
rect 11760 6940 13360 7100
rect 23460 7030 23510 7100
rect 23880 7100 25910 7270
rect 23880 7030 23940 7100
rect 23460 7000 23940 7030
rect 25860 7030 25910 7100
rect 26280 7100 29270 7270
rect 26280 7030 26340 7100
rect 25860 7000 26340 7030
rect 11760 6700 11940 6940
rect 12180 6700 12270 6940
rect 12510 6700 12610 6940
rect 12850 6700 12940 6940
rect 13180 6700 13360 6940
rect 11760 6670 13360 6700
rect 1540 6640 3140 6670
rect 17610 2500 21610 6760
rect 22420 2600 22900 2630
rect 22420 2500 22480 2600
rect 17610 2360 22480 2500
rect 22850 2500 22900 2600
rect 26900 2600 27380 2630
rect 26900 2500 26960 2600
rect 22850 2360 26960 2500
rect 27330 2360 27380 2600
rect 17610 2100 27380 2360
rect 1080 -790 2680 -760
rect 1080 -1030 1260 -790
rect 1500 -1030 1590 -790
rect 1830 -1030 1930 -790
rect 2170 -1030 2260 -790
rect 2500 -1030 2680 -790
rect 1080 -1040 2680 -1030
rect 12220 -790 13820 -760
rect 12220 -1030 12400 -790
rect 12640 -1030 12730 -790
rect 12970 -1030 13070 -790
rect 13310 -1030 13400 -790
rect 13640 -1030 13820 -790
rect 12220 -1040 13820 -1030
rect 17610 -1040 21610 2100
rect 28580 1440 29270 7100
rect 22080 1040 29270 1440
rect 31100 7830 38500 7910
rect 31100 7590 31180 7830
rect 31420 7590 31510 7830
rect 31750 7590 31840 7830
rect 32080 7590 32170 7830
rect 32410 7590 32500 7830
rect 32740 7590 32830 7830
rect 33070 7590 33160 7830
rect 33400 7590 33490 7830
rect 33730 7590 33820 7830
rect 34060 7590 34150 7830
rect 34390 7590 34480 7830
rect 34720 7590 34810 7830
rect 35050 7590 35140 7830
rect 35380 7590 35470 7830
rect 35710 7590 35800 7830
rect 36040 7590 36130 7830
rect 36370 7590 36460 7830
rect 36700 7590 36790 7830
rect 37030 7590 37120 7830
rect 37360 7590 37450 7830
rect 37690 7770 38500 7830
rect 37690 7590 38230 7770
rect 31100 7530 38230 7590
rect 38470 7530 38500 7770
rect 31100 7500 38500 7530
rect 31100 7260 31180 7500
rect 31420 7260 31510 7500
rect 31750 7260 31840 7500
rect 32080 7260 32170 7500
rect 32410 7260 32500 7500
rect 32740 7260 32830 7500
rect 33070 7260 33160 7500
rect 33400 7260 33490 7500
rect 33730 7260 33820 7500
rect 34060 7260 34150 7500
rect 34390 7260 34480 7500
rect 34720 7260 34810 7500
rect 35050 7260 35140 7500
rect 35380 7260 35470 7500
rect 35710 7260 35800 7500
rect 36040 7260 36130 7500
rect 36370 7260 36460 7500
rect 36700 7260 36790 7500
rect 37030 7260 37120 7500
rect 37360 7260 37450 7500
rect 37690 7440 38500 7500
rect 37690 7260 38230 7440
rect 31100 7200 38230 7260
rect 38470 7200 38500 7440
rect 31100 7170 38500 7200
rect 31100 6930 31180 7170
rect 31420 6930 31510 7170
rect 31750 6930 31840 7170
rect 32080 6930 32170 7170
rect 32410 6930 32500 7170
rect 32740 6930 32830 7170
rect 33070 6930 33160 7170
rect 33400 6930 33490 7170
rect 33730 6930 33820 7170
rect 34060 6930 34150 7170
rect 34390 6930 34480 7170
rect 34720 6930 34810 7170
rect 35050 6930 35140 7170
rect 35380 6930 35470 7170
rect 35710 6930 35800 7170
rect 36040 6930 36130 7170
rect 36370 6930 36460 7170
rect 36700 6930 36790 7170
rect 37030 6930 37120 7170
rect 37360 6930 37450 7170
rect 37690 7070 38500 7170
rect 37690 6930 38230 7070
rect 31100 6840 38230 6930
rect 31100 6600 31180 6840
rect 31420 6600 31510 6840
rect 31750 6600 31840 6840
rect 32080 6600 32170 6840
rect 32410 6600 32500 6840
rect 32740 6600 32830 6840
rect 33070 6600 33160 6840
rect 33400 6600 33490 6840
rect 33730 6600 33820 6840
rect 34060 6600 34150 6840
rect 34390 6600 34480 6840
rect 34720 6600 34810 6840
rect 35050 6600 35140 6840
rect 35380 6600 35470 6840
rect 35710 6600 35800 6840
rect 36040 6600 36130 6840
rect 36370 6600 36460 6840
rect 36700 6600 36790 6840
rect 37030 6600 37120 6840
rect 37360 6600 37450 6840
rect 37690 6830 38230 6840
rect 38470 6830 38500 7070
rect 37690 6740 38500 6830
rect 37690 6600 38230 6740
rect 31100 6510 38230 6600
rect 31100 6270 31180 6510
rect 31420 6270 31510 6510
rect 31750 6270 31840 6510
rect 32080 6270 32170 6510
rect 32410 6270 32500 6510
rect 32740 6270 32830 6510
rect 33070 6270 33160 6510
rect 33400 6270 33490 6510
rect 33730 6270 33820 6510
rect 34060 6270 34150 6510
rect 34390 6270 34480 6510
rect 34720 6270 34810 6510
rect 35050 6270 35140 6510
rect 35380 6270 35470 6510
rect 35710 6270 35800 6510
rect 36040 6270 36130 6510
rect 36370 6270 36460 6510
rect 36700 6270 36790 6510
rect 37030 6270 37120 6510
rect 37360 6270 37450 6510
rect 37690 6500 38230 6510
rect 38470 6500 38500 6740
rect 37690 6410 38500 6500
rect 37690 6270 38230 6410
rect 31100 6180 38230 6270
rect 31100 5940 31180 6180
rect 31420 5940 31510 6180
rect 31750 5940 31840 6180
rect 32080 5940 32170 6180
rect 32410 5940 32500 6180
rect 32740 5940 32830 6180
rect 33070 5940 33160 6180
rect 33400 5940 33490 6180
rect 33730 5940 33820 6180
rect 34060 5940 34150 6180
rect 34390 5940 34480 6180
rect 34720 5940 34810 6180
rect 35050 5940 35140 6180
rect 35380 5940 35470 6180
rect 35710 5940 35800 6180
rect 36040 5940 36130 6180
rect 36370 5940 36460 6180
rect 36700 5940 36790 6180
rect 37030 5940 37120 6180
rect 37360 5940 37450 6180
rect 37690 6170 38230 6180
rect 38470 6170 38500 6410
rect 37690 6080 38500 6170
rect 37690 5940 38230 6080
rect 31100 5850 38230 5940
rect 31100 5610 31180 5850
rect 31420 5610 31510 5850
rect 31750 5610 31840 5850
rect 32080 5610 32170 5850
rect 32410 5610 32500 5850
rect 32740 5610 32830 5850
rect 33070 5610 33160 5850
rect 33400 5610 33490 5850
rect 33730 5610 33820 5850
rect 34060 5610 34150 5850
rect 34390 5610 34480 5850
rect 34720 5610 34810 5850
rect 35050 5610 35140 5850
rect 35380 5610 35470 5850
rect 35710 5610 35800 5850
rect 36040 5610 36130 5850
rect 36370 5610 36460 5850
rect 36700 5610 36790 5850
rect 37030 5610 37120 5850
rect 37360 5610 37450 5850
rect 37690 5840 38230 5850
rect 38470 5840 38500 6080
rect 37690 5750 38500 5840
rect 37690 5610 38230 5750
rect 31100 5520 38230 5610
rect 31100 5280 31180 5520
rect 31420 5280 31510 5520
rect 31750 5280 31840 5520
rect 32080 5280 32170 5520
rect 32410 5280 32500 5520
rect 32740 5280 32830 5520
rect 33070 5280 33160 5520
rect 33400 5280 33490 5520
rect 33730 5280 33820 5520
rect 34060 5280 34150 5520
rect 34390 5280 34480 5520
rect 34720 5280 34810 5520
rect 35050 5280 35140 5520
rect 35380 5280 35470 5520
rect 35710 5280 35800 5520
rect 36040 5280 36130 5520
rect 36370 5280 36460 5520
rect 36700 5280 36790 5520
rect 37030 5280 37120 5520
rect 37360 5280 37450 5520
rect 37690 5510 38230 5520
rect 38470 5510 38500 5750
rect 37690 5420 38500 5510
rect 37690 5280 38230 5420
rect 31100 5190 38230 5280
rect 31100 4950 31180 5190
rect 31420 4950 31510 5190
rect 31750 4950 31840 5190
rect 32080 4950 32170 5190
rect 32410 4950 32500 5190
rect 32740 4950 32830 5190
rect 33070 4950 33160 5190
rect 33400 4950 33490 5190
rect 33730 4950 33820 5190
rect 34060 4950 34150 5190
rect 34390 4950 34480 5190
rect 34720 4950 34810 5190
rect 35050 4950 35140 5190
rect 35380 4950 35470 5190
rect 35710 4950 35800 5190
rect 36040 4950 36130 5190
rect 36370 4950 36460 5190
rect 36700 4950 36790 5190
rect 37030 4950 37120 5190
rect 37360 4950 37450 5190
rect 37690 5180 38230 5190
rect 38470 5180 38500 5420
rect 37690 5090 38500 5180
rect 37690 4950 38230 5090
rect 31100 4860 38230 4950
rect 31100 4620 31180 4860
rect 31420 4620 31510 4860
rect 31750 4620 31840 4860
rect 32080 4620 32170 4860
rect 32410 4620 32500 4860
rect 32740 4620 32830 4860
rect 33070 4620 33160 4860
rect 33400 4620 33490 4860
rect 33730 4620 33820 4860
rect 34060 4620 34150 4860
rect 34390 4620 34480 4860
rect 34720 4620 34810 4860
rect 35050 4620 35140 4860
rect 35380 4620 35470 4860
rect 35710 4620 35800 4860
rect 36040 4620 36130 4860
rect 36370 4620 36460 4860
rect 36700 4620 36790 4860
rect 37030 4620 37120 4860
rect 37360 4620 37450 4860
rect 37690 4850 38230 4860
rect 38470 4850 38500 5090
rect 37690 4760 38500 4850
rect 37690 4620 38230 4760
rect 31100 4530 38230 4620
rect 31100 4290 31180 4530
rect 31420 4290 31510 4530
rect 31750 4290 31840 4530
rect 32080 4290 32170 4530
rect 32410 4290 32500 4530
rect 32740 4290 32830 4530
rect 33070 4290 33160 4530
rect 33400 4290 33490 4530
rect 33730 4290 33820 4530
rect 34060 4290 34150 4530
rect 34390 4290 34480 4530
rect 34720 4290 34810 4530
rect 35050 4290 35140 4530
rect 35380 4290 35470 4530
rect 35710 4290 35800 4530
rect 36040 4290 36130 4530
rect 36370 4290 36460 4530
rect 36700 4290 36790 4530
rect 37030 4290 37120 4530
rect 37360 4290 37450 4530
rect 37690 4520 38230 4530
rect 38470 4520 38500 4760
rect 37690 4430 38500 4520
rect 37690 4290 38230 4430
rect 31100 4200 38230 4290
rect 31100 3960 31180 4200
rect 31420 3960 31510 4200
rect 31750 3960 31840 4200
rect 32080 3960 32170 4200
rect 32410 3960 32500 4200
rect 32740 3960 32830 4200
rect 33070 3960 33160 4200
rect 33400 3960 33490 4200
rect 33730 3960 33820 4200
rect 34060 3960 34150 4200
rect 34390 3960 34480 4200
rect 34720 3960 34810 4200
rect 35050 3960 35140 4200
rect 35380 3960 35470 4200
rect 35710 3960 35800 4200
rect 36040 3960 36130 4200
rect 36370 3960 36460 4200
rect 36700 3960 36790 4200
rect 37030 3960 37120 4200
rect 37360 3960 37450 4200
rect 37690 4190 38230 4200
rect 38470 4190 38500 4430
rect 37690 4060 38500 4190
rect 37690 3960 38230 4060
rect 31100 3870 38230 3960
rect 31100 3630 31180 3870
rect 31420 3630 31510 3870
rect 31750 3630 31840 3870
rect 32080 3630 32170 3870
rect 32410 3630 32500 3870
rect 32740 3630 32830 3870
rect 33070 3630 33160 3870
rect 33400 3630 33490 3870
rect 33730 3630 33820 3870
rect 34060 3630 34150 3870
rect 34390 3630 34480 3870
rect 34720 3630 34810 3870
rect 35050 3630 35140 3870
rect 35380 3630 35470 3870
rect 35710 3630 35800 3870
rect 36040 3630 36130 3870
rect 36370 3630 36460 3870
rect 36700 3630 36790 3870
rect 37030 3630 37120 3870
rect 37360 3630 37450 3870
rect 37690 3820 38230 3870
rect 38470 3820 38500 4060
rect 37690 3730 38500 3820
rect 37690 3630 38230 3730
rect 31100 3540 38230 3630
rect 31100 3300 31180 3540
rect 31420 3300 31510 3540
rect 31750 3300 31840 3540
rect 32080 3300 32170 3540
rect 32410 3300 32500 3540
rect 32740 3300 32830 3540
rect 33070 3300 33160 3540
rect 33400 3300 33490 3540
rect 33730 3300 33820 3540
rect 34060 3300 34150 3540
rect 34390 3300 34480 3540
rect 34720 3300 34810 3540
rect 35050 3300 35140 3540
rect 35380 3300 35470 3540
rect 35710 3300 35800 3540
rect 36040 3300 36130 3540
rect 36370 3300 36460 3540
rect 36700 3300 36790 3540
rect 37030 3300 37120 3540
rect 37360 3300 37450 3540
rect 37690 3490 38230 3540
rect 38470 3490 38500 3730
rect 37690 3400 38500 3490
rect 37690 3300 38230 3400
rect 31100 3210 38230 3300
rect 31100 2970 31180 3210
rect 31420 2970 31510 3210
rect 31750 2970 31840 3210
rect 32080 2970 32170 3210
rect 32410 2970 32500 3210
rect 32740 2970 32830 3210
rect 33070 2970 33160 3210
rect 33400 2970 33490 3210
rect 33730 2970 33820 3210
rect 34060 2970 34150 3210
rect 34390 2970 34480 3210
rect 34720 2970 34810 3210
rect 35050 2970 35140 3210
rect 35380 2970 35470 3210
rect 35710 2970 35800 3210
rect 36040 2970 36130 3210
rect 36370 2970 36460 3210
rect 36700 2970 36790 3210
rect 37030 2970 37120 3210
rect 37360 2970 37450 3210
rect 37690 3160 38230 3210
rect 38470 3160 38500 3400
rect 37690 3070 38500 3160
rect 37690 2970 38230 3070
rect 31100 2880 38230 2970
rect 31100 2640 31180 2880
rect 31420 2640 31510 2880
rect 31750 2640 31840 2880
rect 32080 2640 32170 2880
rect 32410 2640 32500 2880
rect 32740 2640 32830 2880
rect 33070 2640 33160 2880
rect 33400 2640 33490 2880
rect 33730 2640 33820 2880
rect 34060 2640 34150 2880
rect 34390 2640 34480 2880
rect 34720 2640 34810 2880
rect 35050 2640 35140 2880
rect 35380 2640 35470 2880
rect 35710 2640 35800 2880
rect 36040 2640 36130 2880
rect 36370 2640 36460 2880
rect 36700 2640 36790 2880
rect 37030 2640 37120 2880
rect 37360 2640 37450 2880
rect 37690 2830 38230 2880
rect 38470 2830 38500 3070
rect 37690 2740 38500 2830
rect 37690 2640 38230 2740
rect 31100 2550 38230 2640
rect 31100 2310 31180 2550
rect 31420 2310 31510 2550
rect 31750 2310 31840 2550
rect 32080 2310 32170 2550
rect 32410 2310 32500 2550
rect 32740 2310 32830 2550
rect 33070 2310 33160 2550
rect 33400 2310 33490 2550
rect 33730 2310 33820 2550
rect 34060 2310 34150 2550
rect 34390 2310 34480 2550
rect 34720 2310 34810 2550
rect 35050 2310 35140 2550
rect 35380 2310 35470 2550
rect 35710 2310 35800 2550
rect 36040 2310 36130 2550
rect 36370 2310 36460 2550
rect 36700 2310 36790 2550
rect 37030 2310 37120 2550
rect 37360 2310 37450 2550
rect 37690 2500 38230 2550
rect 38470 2500 38500 2740
rect 37690 2410 38500 2500
rect 37690 2310 38230 2410
rect 31100 2220 38230 2310
rect 31100 1980 31180 2220
rect 31420 1980 31510 2220
rect 31750 1980 31840 2220
rect 32080 1980 32170 2220
rect 32410 1980 32500 2220
rect 32740 1980 32830 2220
rect 33070 1980 33160 2220
rect 33400 1980 33490 2220
rect 33730 1980 33820 2220
rect 34060 1980 34150 2220
rect 34390 1980 34480 2220
rect 34720 1980 34810 2220
rect 35050 1980 35140 2220
rect 35380 1980 35470 2220
rect 35710 1980 35800 2220
rect 36040 1980 36130 2220
rect 36370 1980 36460 2220
rect 36700 1980 36790 2220
rect 37030 1980 37120 2220
rect 37360 1980 37450 2220
rect 37690 2170 38230 2220
rect 38470 2170 38500 2410
rect 37690 2080 38500 2170
rect 37690 1980 38230 2080
rect 31100 1890 38230 1980
rect 31100 1650 31180 1890
rect 31420 1650 31510 1890
rect 31750 1650 31840 1890
rect 32080 1650 32170 1890
rect 32410 1650 32500 1890
rect 32740 1650 32830 1890
rect 33070 1650 33160 1890
rect 33400 1650 33490 1890
rect 33730 1650 33820 1890
rect 34060 1650 34150 1890
rect 34390 1650 34480 1890
rect 34720 1650 34810 1890
rect 35050 1650 35140 1890
rect 35380 1650 35470 1890
rect 35710 1650 35800 1890
rect 36040 1650 36130 1890
rect 36370 1650 36460 1890
rect 36700 1650 36790 1890
rect 37030 1650 37120 1890
rect 37360 1650 37450 1890
rect 37690 1840 38230 1890
rect 38470 1840 38500 2080
rect 37690 1750 38500 1840
rect 37690 1650 38230 1750
rect 31100 1560 38230 1650
rect 31100 1320 31180 1560
rect 31420 1320 31510 1560
rect 31750 1320 31840 1560
rect 32080 1320 32170 1560
rect 32410 1320 32500 1560
rect 32740 1320 32830 1560
rect 33070 1320 33160 1560
rect 33400 1320 33490 1560
rect 33730 1320 33820 1560
rect 34060 1320 34150 1560
rect 34390 1320 34480 1560
rect 34720 1320 34810 1560
rect 35050 1320 35140 1560
rect 35380 1320 35470 1560
rect 35710 1320 35800 1560
rect 36040 1320 36130 1560
rect 36370 1320 36460 1560
rect 36700 1320 36790 1560
rect 37030 1320 37120 1560
rect 37360 1320 37450 1560
rect 37690 1510 38230 1560
rect 38470 1510 38500 1750
rect 37690 1420 38500 1510
rect 37690 1320 38230 1420
rect 31100 1180 38230 1320
rect 38470 1180 38500 1420
rect 23460 980 23940 1040
rect 23460 740 23510 980
rect 23880 740 23940 980
rect 23460 710 23940 740
rect 25860 980 26340 1040
rect 25860 740 25910 980
rect 26280 740 26340 980
rect 25860 710 26340 740
rect -170 -1840 21610 -1040
rect -6530 -2720 14530 -2160
rect -6530 -2960 1720 -2720
rect 1960 -2960 2050 -2720
rect 2290 -2960 2390 -2720
rect 2630 -2960 2720 -2720
rect 2960 -2960 11940 -2720
rect 12180 -2960 12270 -2720
rect 12510 -2960 12610 -2720
rect 12850 -2960 12940 -2720
rect 13180 -2960 14530 -2720
rect -6530 -11680 -2830 -2960
rect 1540 -2990 3140 -2960
rect 11760 -2990 13360 -2960
rect 17610 -3840 21610 -1840
rect 31100 230 38500 1180
rect 31100 -10 31180 230
rect 31420 -10 31510 230
rect 31750 -10 31840 230
rect 32080 -10 32170 230
rect 32410 -10 32500 230
rect 32740 -10 32830 230
rect 33070 -10 33160 230
rect 33400 -10 33490 230
rect 33730 -10 33820 230
rect 34060 -10 34150 230
rect 34390 -10 34480 230
rect 34720 -10 34810 230
rect 35050 -10 35140 230
rect 35380 -10 35470 230
rect 35710 -10 35800 230
rect 36040 -10 36130 230
rect 36370 -10 36460 230
rect 36700 -10 36790 230
rect 37030 -10 37120 230
rect 37360 -10 37450 230
rect 37690 170 38500 230
rect 37690 -10 38230 170
rect 31100 -70 38230 -10
rect 38470 -70 38500 170
rect 31100 -100 38500 -70
rect 31100 -340 31180 -100
rect 31420 -340 31510 -100
rect 31750 -340 31840 -100
rect 32080 -340 32170 -100
rect 32410 -340 32500 -100
rect 32740 -340 32830 -100
rect 33070 -340 33160 -100
rect 33400 -340 33490 -100
rect 33730 -340 33820 -100
rect 34060 -340 34150 -100
rect 34390 -340 34480 -100
rect 34720 -340 34810 -100
rect 35050 -340 35140 -100
rect 35380 -340 35470 -100
rect 35710 -340 35800 -100
rect 36040 -340 36130 -100
rect 36370 -340 36460 -100
rect 36700 -340 36790 -100
rect 37030 -340 37120 -100
rect 37360 -340 37450 -100
rect 37690 -160 38500 -100
rect 37690 -340 38230 -160
rect 31100 -400 38230 -340
rect 38470 -400 38500 -160
rect 31100 -430 38500 -400
rect 31100 -670 31180 -430
rect 31420 -670 31510 -430
rect 31750 -670 31840 -430
rect 32080 -670 32170 -430
rect 32410 -670 32500 -430
rect 32740 -670 32830 -430
rect 33070 -670 33160 -430
rect 33400 -670 33490 -430
rect 33730 -670 33820 -430
rect 34060 -670 34150 -430
rect 34390 -670 34480 -430
rect 34720 -670 34810 -430
rect 35050 -670 35140 -430
rect 35380 -670 35470 -430
rect 35710 -670 35800 -430
rect 36040 -670 36130 -430
rect 36370 -670 36460 -430
rect 36700 -670 36790 -430
rect 37030 -670 37120 -430
rect 37360 -670 37450 -430
rect 37690 -530 38500 -430
rect 37690 -670 38230 -530
rect 31100 -760 38230 -670
rect 31100 -1000 31180 -760
rect 31420 -1000 31510 -760
rect 31750 -1000 31840 -760
rect 32080 -1000 32170 -760
rect 32410 -1000 32500 -760
rect 32740 -1000 32830 -760
rect 33070 -1000 33160 -760
rect 33400 -1000 33490 -760
rect 33730 -1000 33820 -760
rect 34060 -1000 34150 -760
rect 34390 -1000 34480 -760
rect 34720 -1000 34810 -760
rect 35050 -1000 35140 -760
rect 35380 -1000 35470 -760
rect 35710 -1000 35800 -760
rect 36040 -1000 36130 -760
rect 36370 -1000 36460 -760
rect 36700 -1000 36790 -760
rect 37030 -1000 37120 -760
rect 37360 -1000 37450 -760
rect 37690 -770 38230 -760
rect 38470 -770 38500 -530
rect 37690 -860 38500 -770
rect 37690 -1000 38230 -860
rect 31100 -1090 38230 -1000
rect 31100 -1330 31180 -1090
rect 31420 -1330 31510 -1090
rect 31750 -1330 31840 -1090
rect 32080 -1330 32170 -1090
rect 32410 -1330 32500 -1090
rect 32740 -1330 32830 -1090
rect 33070 -1330 33160 -1090
rect 33400 -1330 33490 -1090
rect 33730 -1330 33820 -1090
rect 34060 -1330 34150 -1090
rect 34390 -1330 34480 -1090
rect 34720 -1330 34810 -1090
rect 35050 -1330 35140 -1090
rect 35380 -1330 35470 -1090
rect 35710 -1330 35800 -1090
rect 36040 -1330 36130 -1090
rect 36370 -1330 36460 -1090
rect 36700 -1330 36790 -1090
rect 37030 -1330 37120 -1090
rect 37360 -1330 37450 -1090
rect 37690 -1100 38230 -1090
rect 38470 -1100 38500 -860
rect 37690 -1190 38500 -1100
rect 37690 -1330 38230 -1190
rect 31100 -1420 38230 -1330
rect 31100 -1660 31180 -1420
rect 31420 -1660 31510 -1420
rect 31750 -1660 31840 -1420
rect 32080 -1660 32170 -1420
rect 32410 -1660 32500 -1420
rect 32740 -1660 32830 -1420
rect 33070 -1660 33160 -1420
rect 33400 -1660 33490 -1420
rect 33730 -1660 33820 -1420
rect 34060 -1660 34150 -1420
rect 34390 -1660 34480 -1420
rect 34720 -1660 34810 -1420
rect 35050 -1660 35140 -1420
rect 35380 -1660 35470 -1420
rect 35710 -1660 35800 -1420
rect 36040 -1660 36130 -1420
rect 36370 -1660 36460 -1420
rect 36700 -1660 36790 -1420
rect 37030 -1660 37120 -1420
rect 37360 -1660 37450 -1420
rect 37690 -1430 38230 -1420
rect 38470 -1430 38500 -1190
rect 37690 -1520 38500 -1430
rect 37690 -1660 38230 -1520
rect 31100 -1750 38230 -1660
rect 31100 -1990 31180 -1750
rect 31420 -1990 31510 -1750
rect 31750 -1990 31840 -1750
rect 32080 -1990 32170 -1750
rect 32410 -1990 32500 -1750
rect 32740 -1990 32830 -1750
rect 33070 -1990 33160 -1750
rect 33400 -1990 33490 -1750
rect 33730 -1990 33820 -1750
rect 34060 -1990 34150 -1750
rect 34390 -1990 34480 -1750
rect 34720 -1990 34810 -1750
rect 35050 -1990 35140 -1750
rect 35380 -1990 35470 -1750
rect 35710 -1990 35800 -1750
rect 36040 -1990 36130 -1750
rect 36370 -1990 36460 -1750
rect 36700 -1990 36790 -1750
rect 37030 -1990 37120 -1750
rect 37360 -1990 37450 -1750
rect 37690 -1760 38230 -1750
rect 38470 -1760 38500 -1520
rect 37690 -1850 38500 -1760
rect 37690 -1990 38230 -1850
rect 31100 -2080 38230 -1990
rect 31100 -2320 31180 -2080
rect 31420 -2320 31510 -2080
rect 31750 -2320 31840 -2080
rect 32080 -2320 32170 -2080
rect 32410 -2320 32500 -2080
rect 32740 -2320 32830 -2080
rect 33070 -2320 33160 -2080
rect 33400 -2320 33490 -2080
rect 33730 -2320 33820 -2080
rect 34060 -2320 34150 -2080
rect 34390 -2320 34480 -2080
rect 34720 -2320 34810 -2080
rect 35050 -2320 35140 -2080
rect 35380 -2320 35470 -2080
rect 35710 -2320 35800 -2080
rect 36040 -2320 36130 -2080
rect 36370 -2320 36460 -2080
rect 36700 -2320 36790 -2080
rect 37030 -2320 37120 -2080
rect 37360 -2320 37450 -2080
rect 37690 -2090 38230 -2080
rect 38470 -2090 38500 -1850
rect 37690 -2180 38500 -2090
rect 37690 -2320 38230 -2180
rect 31100 -2410 38230 -2320
rect 31100 -2650 31180 -2410
rect 31420 -2650 31510 -2410
rect 31750 -2650 31840 -2410
rect 32080 -2650 32170 -2410
rect 32410 -2650 32500 -2410
rect 32740 -2650 32830 -2410
rect 33070 -2650 33160 -2410
rect 33400 -2650 33490 -2410
rect 33730 -2650 33820 -2410
rect 34060 -2650 34150 -2410
rect 34390 -2650 34480 -2410
rect 34720 -2650 34810 -2410
rect 35050 -2650 35140 -2410
rect 35380 -2650 35470 -2410
rect 35710 -2650 35800 -2410
rect 36040 -2650 36130 -2410
rect 36370 -2650 36460 -2410
rect 36700 -2650 36790 -2410
rect 37030 -2650 37120 -2410
rect 37360 -2650 37450 -2410
rect 37690 -2420 38230 -2410
rect 38470 -2420 38500 -2180
rect 37690 -2510 38500 -2420
rect 37690 -2650 38230 -2510
rect 31100 -2740 38230 -2650
rect 31100 -2980 31180 -2740
rect 31420 -2980 31510 -2740
rect 31750 -2980 31840 -2740
rect 32080 -2980 32170 -2740
rect 32410 -2980 32500 -2740
rect 32740 -2980 32830 -2740
rect 33070 -2980 33160 -2740
rect 33400 -2980 33490 -2740
rect 33730 -2980 33820 -2740
rect 34060 -2980 34150 -2740
rect 34390 -2980 34480 -2740
rect 34720 -2980 34810 -2740
rect 35050 -2980 35140 -2740
rect 35380 -2980 35470 -2740
rect 35710 -2980 35800 -2740
rect 36040 -2980 36130 -2740
rect 36370 -2980 36460 -2740
rect 36700 -2980 36790 -2740
rect 37030 -2980 37120 -2740
rect 37360 -2980 37450 -2740
rect 37690 -2750 38230 -2740
rect 38470 -2750 38500 -2510
rect 37690 -2840 38500 -2750
rect 37690 -2980 38230 -2840
rect 31100 -3070 38230 -2980
rect 31100 -3310 31180 -3070
rect 31420 -3310 31510 -3070
rect 31750 -3310 31840 -3070
rect 32080 -3310 32170 -3070
rect 32410 -3310 32500 -3070
rect 32740 -3310 32830 -3070
rect 33070 -3310 33160 -3070
rect 33400 -3310 33490 -3070
rect 33730 -3310 33820 -3070
rect 34060 -3310 34150 -3070
rect 34390 -3310 34480 -3070
rect 34720 -3310 34810 -3070
rect 35050 -3310 35140 -3070
rect 35380 -3310 35470 -3070
rect 35710 -3310 35800 -3070
rect 36040 -3310 36130 -3070
rect 36370 -3310 36460 -3070
rect 36700 -3310 36790 -3070
rect 37030 -3310 37120 -3070
rect 37360 -3310 37450 -3070
rect 37690 -3080 38230 -3070
rect 38470 -3080 38500 -2840
rect 37690 -3170 38500 -3080
rect 37690 -3310 38230 -3170
rect 31100 -3400 38230 -3310
rect 31100 -3640 31180 -3400
rect 31420 -3640 31510 -3400
rect 31750 -3640 31840 -3400
rect 32080 -3640 32170 -3400
rect 32410 -3640 32500 -3400
rect 32740 -3640 32830 -3400
rect 33070 -3640 33160 -3400
rect 33400 -3640 33490 -3400
rect 33730 -3640 33820 -3400
rect 34060 -3640 34150 -3400
rect 34390 -3640 34480 -3400
rect 34720 -3640 34810 -3400
rect 35050 -3640 35140 -3400
rect 35380 -3640 35470 -3400
rect 35710 -3640 35800 -3400
rect 36040 -3640 36130 -3400
rect 36370 -3640 36460 -3400
rect 36700 -3640 36790 -3400
rect 37030 -3640 37120 -3400
rect 37360 -3640 37450 -3400
rect 37690 -3410 38230 -3400
rect 38470 -3410 38500 -3170
rect 37690 -3540 38500 -3410
rect 37690 -3640 38230 -3540
rect 22420 -3690 22900 -3660
rect 22420 -3840 22480 -3690
rect 17610 -3930 22480 -3840
rect 22850 -3840 22900 -3690
rect 26900 -3690 27380 -3660
rect 26900 -3840 26960 -3690
rect 22850 -3930 26960 -3840
rect 27330 -3840 27380 -3690
rect 31100 -3730 38230 -3640
rect 31100 -3840 31180 -3730
rect 27330 -3850 29220 -3840
rect 30380 -3850 31180 -3840
rect 27330 -3930 31180 -3850
rect 17610 -3970 31180 -3930
rect 31420 -3970 31510 -3730
rect 31750 -3970 31840 -3730
rect 32080 -3970 32170 -3730
rect 32410 -3970 32500 -3730
rect 32740 -3970 32830 -3730
rect 33070 -3970 33160 -3730
rect 33400 -3970 33490 -3730
rect 33730 -3970 33820 -3730
rect 34060 -3970 34150 -3730
rect 34390 -3970 34480 -3730
rect 34720 -3970 34810 -3730
rect 35050 -3970 35140 -3730
rect 35380 -3970 35470 -3730
rect 35710 -3970 35800 -3730
rect 36040 -3970 36130 -3730
rect 36370 -3970 36460 -3730
rect 36700 -3970 36790 -3730
rect 37030 -3970 37120 -3730
rect 37360 -3970 37450 -3730
rect 37690 -3780 38230 -3730
rect 38470 -3780 38500 -3540
rect 37690 -3870 38500 -3780
rect 37690 -3970 38230 -3870
rect 17610 -4060 38230 -3970
rect 17610 -4240 31180 -4060
rect -1350 -4840 260 -4630
rect -1350 -5080 -1180 -4840
rect -940 -5080 -850 -4840
rect -610 -5080 -520 -4840
rect -280 -5080 -190 -4840
rect 50 -5080 260 -4840
rect -1350 -5170 260 -5080
rect -1350 -5410 -1180 -5170
rect -940 -5410 -850 -5170
rect -610 -5410 -520 -5170
rect -280 -5410 -190 -5170
rect 50 -5410 260 -5170
rect -1350 -5500 260 -5410
rect -1350 -5740 -1180 -5500
rect -940 -5740 -850 -5500
rect -610 -5740 -520 -5500
rect -280 -5740 -190 -5500
rect 50 -5740 260 -5500
rect -1350 -5830 260 -5740
rect -1350 -6070 -1180 -5830
rect -940 -6070 -850 -5830
rect -610 -6070 -520 -5830
rect -280 -6070 -190 -5830
rect 50 -6070 260 -5830
rect -1350 -6370 260 -6070
rect -1350 -6610 -1170 -6370
rect -930 -6610 -840 -6370
rect -600 -6610 -510 -6370
rect -270 -6610 -180 -6370
rect 60 -6610 260 -6370
rect -1350 -6640 260 -6610
rect 14520 -4840 16130 -4630
rect 14520 -5080 14730 -4840
rect 14970 -5080 15060 -4840
rect 15300 -5080 15390 -4840
rect 15630 -5080 15720 -4840
rect 15960 -5080 16130 -4840
rect 14520 -5170 16130 -5080
rect 14520 -5410 14730 -5170
rect 14970 -5410 15060 -5170
rect 15300 -5410 15390 -5170
rect 15630 -5410 15720 -5170
rect 15960 -5410 16130 -5170
rect 14520 -5500 16130 -5410
rect 14520 -5740 14730 -5500
rect 14970 -5740 15060 -5500
rect 15300 -5740 15390 -5500
rect 15630 -5740 15720 -5500
rect 15960 -5740 16130 -5500
rect 14520 -5830 16130 -5740
rect 14520 -6070 14730 -5830
rect 14970 -6070 15060 -5830
rect 15300 -6070 15390 -5830
rect 15630 -6070 15720 -5830
rect 15960 -6070 16130 -5830
rect 14520 -6370 16130 -6070
rect 14520 -6610 14720 -6370
rect 14960 -6610 15050 -6370
rect 15290 -6610 15380 -6370
rect 15620 -6610 15710 -6370
rect 15950 -6610 16130 -6370
rect 14520 -6640 16130 -6610
rect 17610 -8330 21610 -4240
rect 29220 -4250 30380 -4240
rect 31100 -4300 31180 -4240
rect 31420 -4300 31510 -4060
rect 31750 -4300 31840 -4060
rect 32080 -4300 32170 -4060
rect 32410 -4300 32500 -4060
rect 32740 -4300 32830 -4060
rect 33070 -4300 33160 -4060
rect 33400 -4300 33490 -4060
rect 33730 -4300 33820 -4060
rect 34060 -4300 34150 -4060
rect 34390 -4300 34480 -4060
rect 34720 -4300 34810 -4060
rect 35050 -4300 35140 -4060
rect 35380 -4300 35470 -4060
rect 35710 -4300 35800 -4060
rect 36040 -4300 36130 -4060
rect 36370 -4300 36460 -4060
rect 36700 -4300 36790 -4060
rect 37030 -4300 37120 -4060
rect 37360 -4300 37450 -4060
rect 37690 -4110 38230 -4060
rect 38470 -4110 38500 -3870
rect 37690 -4200 38500 -4110
rect 37690 -4300 38230 -4200
rect 31100 -4390 38230 -4300
rect 31100 -4630 31180 -4390
rect 31420 -4630 31510 -4390
rect 31750 -4630 31840 -4390
rect 32080 -4630 32170 -4390
rect 32410 -4630 32500 -4390
rect 32740 -4630 32830 -4390
rect 33070 -4630 33160 -4390
rect 33400 -4630 33490 -4390
rect 33730 -4630 33820 -4390
rect 34060 -4630 34150 -4390
rect 34390 -4630 34480 -4390
rect 34720 -4630 34810 -4390
rect 35050 -4630 35140 -4390
rect 35380 -4630 35470 -4390
rect 35710 -4630 35800 -4390
rect 36040 -4630 36130 -4390
rect 36370 -4630 36460 -4390
rect 36700 -4630 36790 -4390
rect 37030 -4630 37120 -4390
rect 37360 -4630 37450 -4390
rect 37690 -4440 38230 -4390
rect 38470 -4440 38500 -4200
rect 37690 -4530 38500 -4440
rect 37690 -4630 38230 -4530
rect 31100 -4720 38230 -4630
rect 31100 -4960 31180 -4720
rect 31420 -4960 31510 -4720
rect 31750 -4960 31840 -4720
rect 32080 -4960 32170 -4720
rect 32410 -4960 32500 -4720
rect 32740 -4960 32830 -4720
rect 33070 -4960 33160 -4720
rect 33400 -4960 33490 -4720
rect 33730 -4960 33820 -4720
rect 34060 -4960 34150 -4720
rect 34390 -4960 34480 -4720
rect 34720 -4960 34810 -4720
rect 35050 -4960 35140 -4720
rect 35380 -4960 35470 -4720
rect 35710 -4960 35800 -4720
rect 36040 -4960 36130 -4720
rect 36370 -4960 36460 -4720
rect 36700 -4960 36790 -4720
rect 37030 -4960 37120 -4720
rect 37360 -4960 37450 -4720
rect 37690 -4770 38230 -4720
rect 38470 -4770 38500 -4530
rect 37690 -4860 38500 -4770
rect 37690 -4960 38230 -4860
rect 31100 -5050 38230 -4960
rect 31100 -5290 31180 -5050
rect 31420 -5290 31510 -5050
rect 31750 -5290 31840 -5050
rect 32080 -5290 32170 -5050
rect 32410 -5290 32500 -5050
rect 32740 -5290 32830 -5050
rect 33070 -5290 33160 -5050
rect 33400 -5290 33490 -5050
rect 33730 -5290 33820 -5050
rect 34060 -5290 34150 -5050
rect 34390 -5290 34480 -5050
rect 34720 -5290 34810 -5050
rect 35050 -5290 35140 -5050
rect 35380 -5290 35470 -5050
rect 35710 -5290 35800 -5050
rect 36040 -5290 36130 -5050
rect 36370 -5290 36460 -5050
rect 36700 -5290 36790 -5050
rect 37030 -5290 37120 -5050
rect 37360 -5290 37450 -5050
rect 37690 -5100 38230 -5050
rect 38470 -5100 38500 -4860
rect 37690 -5190 38500 -5100
rect 37690 -5290 38230 -5190
rect 31100 -5380 38230 -5290
rect 31100 -5620 31180 -5380
rect 31420 -5620 31510 -5380
rect 31750 -5620 31840 -5380
rect 32080 -5620 32170 -5380
rect 32410 -5620 32500 -5380
rect 32740 -5620 32830 -5380
rect 33070 -5620 33160 -5380
rect 33400 -5620 33490 -5380
rect 33730 -5620 33820 -5380
rect 34060 -5620 34150 -5380
rect 34390 -5620 34480 -5380
rect 34720 -5620 34810 -5380
rect 35050 -5620 35140 -5380
rect 35380 -5620 35470 -5380
rect 35710 -5620 35800 -5380
rect 36040 -5620 36130 -5380
rect 36370 -5620 36460 -5380
rect 36700 -5620 36790 -5380
rect 37030 -5620 37120 -5380
rect 37360 -5620 37450 -5380
rect 37690 -5430 38230 -5380
rect 38470 -5430 38500 -5190
rect 37690 -5520 38500 -5430
rect 37690 -5620 38230 -5520
rect 31100 -5710 38230 -5620
rect 31100 -5950 31180 -5710
rect 31420 -5950 31510 -5710
rect 31750 -5950 31840 -5710
rect 32080 -5950 32170 -5710
rect 32410 -5950 32500 -5710
rect 32740 -5950 32830 -5710
rect 33070 -5950 33160 -5710
rect 33400 -5950 33490 -5710
rect 33730 -5950 33820 -5710
rect 34060 -5950 34150 -5710
rect 34390 -5950 34480 -5710
rect 34720 -5950 34810 -5710
rect 35050 -5950 35140 -5710
rect 35380 -5950 35470 -5710
rect 35710 -5950 35800 -5710
rect 36040 -5950 36130 -5710
rect 36370 -5950 36460 -5710
rect 36700 -5950 36790 -5710
rect 37030 -5950 37120 -5710
rect 37360 -5950 37450 -5710
rect 37690 -5760 38230 -5710
rect 38470 -5760 38500 -5520
rect 37690 -5850 38500 -5760
rect 37690 -5950 38230 -5850
rect 31100 -6040 38230 -5950
rect 31100 -6280 31180 -6040
rect 31420 -6280 31510 -6040
rect 31750 -6280 31840 -6040
rect 32080 -6280 32170 -6040
rect 32410 -6280 32500 -6040
rect 32740 -6280 32830 -6040
rect 33070 -6280 33160 -6040
rect 33400 -6280 33490 -6040
rect 33730 -6280 33820 -6040
rect 34060 -6280 34150 -6040
rect 34390 -6280 34480 -6040
rect 34720 -6280 34810 -6040
rect 35050 -6280 35140 -6040
rect 35380 -6280 35470 -6040
rect 35710 -6280 35800 -6040
rect 36040 -6280 36130 -6040
rect 36370 -6280 36460 -6040
rect 36700 -6280 36790 -6040
rect 37030 -6280 37120 -6040
rect 37360 -6280 37450 -6040
rect 37690 -6090 38230 -6040
rect 38470 -6090 38500 -5850
rect 37690 -6180 38500 -6090
rect 37690 -6280 38230 -6180
rect 31100 -6420 38230 -6280
rect 38470 -6420 38500 -6180
rect 31100 -6450 38500 -6420
rect 17610 -8370 21930 -8330
rect 17610 -8610 21650 -8370
rect 21890 -8610 21930 -8370
rect 17610 -8650 21930 -8610
rect 17610 -9970 21610 -8650
rect 26880 -9970 30100 -9600
rect 1080 -10340 2680 -10310
rect 1080 -10560 1260 -10340
rect 40 -10580 1260 -10560
rect 1500 -10580 1590 -10340
rect 1830 -10580 1930 -10340
rect 2170 -10580 2260 -10340
rect 2500 -10560 2680 -10340
rect 12220 -10370 13820 -10340
rect 12220 -10560 12400 -10370
rect 2500 -10580 12400 -10560
rect 40 -10610 12400 -10580
rect 12640 -10610 12730 -10370
rect 12970 -10610 13070 -10370
rect 13310 -10610 13400 -10370
rect 13640 -10560 13820 -10370
rect 17610 -10370 30100 -9970
rect 17610 -10560 21610 -10370
rect 13640 -10610 21610 -10560
rect 40 -11360 21610 -10610
rect -6530 -12240 13390 -11680
rect -6530 -12480 1690 -12240
rect 1930 -12480 2020 -12240
rect 2260 -12480 2360 -12240
rect 2600 -12480 2690 -12240
rect 2930 -12480 11970 -12240
rect 12210 -12480 12300 -12240
rect 12540 -12480 12640 -12240
rect 12880 -12480 12970 -12240
rect 13210 -12480 13390 -12240
rect 1510 -12510 3110 -12480
rect 11790 -12510 13390 -12480
rect 17610 -13990 21610 -11360
rect 17610 -14030 21930 -13990
rect 17610 -14270 21650 -14030
rect 21890 -14270 21930 -14030
rect 17610 -14310 21930 -14270
rect 17610 -15860 21610 -14310
rect 27160 -15860 30380 -15460
rect 17610 -16260 30380 -15860
rect 17610 -20070 21610 -16260
rect 17610 -20110 21930 -20070
rect 17610 -20350 21650 -20110
rect 21890 -20350 21930 -20110
rect 17610 -20390 21930 -20350
rect 17610 -21680 21610 -20390
rect 26960 -21680 30180 -21340
rect 17610 -22080 30180 -21680
rect 1550 -22660 3150 -22630
rect 1550 -22670 1730 -22660
rect -6530 -22900 1730 -22670
rect 1970 -22900 2060 -22660
rect 2300 -22900 2400 -22660
rect 2640 -22900 2730 -22660
rect 2970 -22670 3150 -22660
rect 11750 -22660 13350 -22630
rect 11750 -22670 11930 -22660
rect 2970 -22900 11930 -22670
rect 12170 -22900 12260 -22660
rect 12500 -22900 12600 -22660
rect 12840 -22900 12930 -22660
rect 13170 -22670 13350 -22660
rect 17610 -22670 21610 -22080
rect 13170 -22900 21610 -22670
rect -6530 -23700 21610 -22900
use sf  sf_0
timestamp 1640986451
transform 1 0 12590 0 1 -29850
box -11690 7000 1410 17380
use core  core_1
timestamp 1637735227
transform 1 0 7320 0 1 -7060
box -7320 -2490 7580 4060
use core  core_0
timestamp 1637735227
transform 1 0 7320 0 1 2520
box -7320 -2490 7580 4060
use cmfb  cmfb_0
timestamp 1634684585
transform 1 0 25700 0 1 2690
box -3910 -30 2310 4270
use cmfb  cmfb_1
timestamp 1634684585
transform 1 0 25700 0 1 -3610
box -3910 -30 2310 4270
use mirror_1  mirror_1_0
timestamp 1635749472
transform 1 0 20860 0 1 -9070
box 840 -570 9240 3290
use mirror_4  mirror_4_0
timestamp 1635749603
transform 1 0 20940 0 1 -20790
box 760 -570 9240 3290
use mirror_3  mirror_3_0
timestamp 1635750117
transform 1 0 21140 0 1 -14930
box 560 -570 9240 3290
<< labels >>
rlabel metal1 13060 40 13060 40 1 GND
port 7 n
rlabel metal5 -2700 7440 -2700 7440 1 VDD
port 1 n
rlabel metal3 8330 2730 8330 2730 1 Vop
rlabel metal3 6540 2730 6540 2730 1 Von
rlabel metal2 7400 360 7400 360 1 Vcm1
rlabel metal3 8870 -6850 8870 -6850 1 pre_Vout_n
rlabel metal3 6040 -6890 6040 -6890 1 pre_Vout_p
rlabel metal2 7420 -9350 7420 -9350 1 Vcm2
rlabel metal2 7620 -3520 7620 -3520 1 Vcmfb2
rlabel metal2 7470 6130 7470 6130 1 Vcmfb1
rlabel metal5 29100 7420 29100 7420 1 VDD
port 1 n
rlabel metal5 -6360 -23210 -6360 -23210 1 GND
port 7 n
rlabel metal4 39610 8360 39610 8360 1 Vb5
port 20 n
rlabel metal4 30970 -10670 30970 -10670 1 Vb1_
port 21 n
rlabel metal4 30890 -16530 30890 -16530 1 Vb3_
port 22 n
rlabel metal4 30660 -22400 30660 -22400 1 Vb4_
port 23 n
rlabel space 7450 21850 7450 21850 1 MIDDLE_TOP
rlabel metal4 21200 8860 21200 8860 1 Vb2
port 19 n
rlabel metal4 8280 8530 8280 8530 1 Vinn
rlabel metal5 20440 21510 20440 21510 1 Iin_n
port 26 n
rlabel metal4 6600 8530 6600 8530 1 Vinp
rlabel metal5 -5530 21540 -5530 21540 1 Iin_p
port 25 n
rlabel metal3 5090 -23580 5090 -23580 1 Vout_p
port 18 n
rlabel metal3 9790 -23610 9790 -23610 1 Vout_n
port 17 n
<< end >>
