* NGSPICE file created from dnwcell.ext - technology: sky130A

.subckt dnwcell Source Gate Drain
X0 Source Gate Drain Source sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

