* NGSPICE file created from sf_half_test.ext - technology: sky130A

.subckt sf_half_test Vout g_u VDD
X0 Vout g_u VDD Vout sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+07u l=320000u M=26
.ends

