magic
tech sky130A
timestamp 1640251702
<< dnwell >>
rect -105 -105 2815 2390
<< isosubstrate >>
rect -155 2430 2865 2440
rect -155 -145 -145 2430
rect 2855 -145 2865 2430
rect -155 -155 2865 -145
<< nwell >>
rect -145 2285 2855 2430
rect -145 0 0 2285
rect 2710 0 2855 2285
rect -145 -145 2855 0
<< pwell >>
rect 0 0 2710 2285
<< nmos >>
rect 105 -345 2605 -300
rect 105 -440 2605 -395
rect 105 -535 2605 -490
rect 105 -630 2605 -585
rect 105 -725 2605 -680
rect 105 -820 2605 -775
rect 105 -915 2605 -870
rect 105 -1010 2605 -965
rect 105 -1105 2605 -1060
rect 105 -1200 2605 -1155
rect 105 -1295 2605 -1250
rect 105 -1390 2605 -1345
rect 105 -1485 2605 -1440
rect 105 -1580 2605 -1535
rect 105 -1675 2605 -1630
rect 105 -1770 2605 -1725
rect 105 -1865 2605 -1820
rect 105 -1960 2605 -1915
rect 105 -2055 2605 -2010
rect 105 -2150 2605 -2105
rect 105 -2245 2605 -2200
rect 105 -2340 2605 -2295
rect 105 -2435 2605 -2390
rect 105 -2530 2605 -2485
rect 105 -2625 2605 -2580
rect 105 -2720 2605 -2675
<< nmoslvt >>
rect 175 2150 2675 2182
rect 175 2068 2675 2100
rect 175 1986 2675 2018
rect 175 1904 2675 1936
rect 175 1822 2675 1854
rect 175 1740 2675 1772
rect 175 1658 2675 1690
rect 175 1576 2675 1608
rect 175 1494 2675 1526
rect 175 1412 2675 1444
rect 175 1330 2675 1362
rect 175 1248 2675 1280
rect 175 1166 2675 1198
rect 175 1084 2675 1116
rect 175 1002 2675 1034
rect 175 920 2675 952
rect 175 838 2675 870
rect 175 756 2675 788
rect 175 674 2675 706
rect 175 592 2675 624
rect 175 510 2675 542
rect 175 428 2675 460
rect 175 346 2675 378
rect 175 264 2675 296
rect 175 182 2675 214
rect 175 100 2675 132
<< ndiff >>
rect 175 2217 2675 2230
rect 175 2197 200 2217
rect 220 2197 240 2217
rect 260 2197 280 2217
rect 300 2197 320 2217
rect 340 2197 360 2217
rect 380 2197 400 2217
rect 420 2197 440 2217
rect 460 2197 480 2217
rect 500 2197 520 2217
rect 540 2197 560 2217
rect 580 2197 600 2217
rect 620 2197 640 2217
rect 660 2197 680 2217
rect 700 2197 720 2217
rect 740 2197 760 2217
rect 780 2197 800 2217
rect 820 2197 840 2217
rect 860 2197 880 2217
rect 900 2197 920 2217
rect 940 2197 960 2217
rect 980 2197 1000 2217
rect 1020 2197 1040 2217
rect 1060 2197 1080 2217
rect 1100 2197 1120 2217
rect 1140 2197 1160 2217
rect 1180 2197 1200 2217
rect 1220 2197 1240 2217
rect 1260 2197 1280 2217
rect 1300 2197 1320 2217
rect 1340 2197 1360 2217
rect 1380 2197 1400 2217
rect 1420 2197 1440 2217
rect 1460 2197 1480 2217
rect 1500 2197 1520 2217
rect 1540 2197 1560 2217
rect 1580 2197 1600 2217
rect 1620 2197 1640 2217
rect 1660 2197 1680 2217
rect 1700 2197 1720 2217
rect 1740 2197 1760 2217
rect 1780 2197 1800 2217
rect 1820 2197 1840 2217
rect 1860 2197 1880 2217
rect 1900 2197 1920 2217
rect 1940 2197 1960 2217
rect 1980 2197 2000 2217
rect 2020 2197 2040 2217
rect 2060 2197 2080 2217
rect 2100 2197 2120 2217
rect 2140 2197 2160 2217
rect 2180 2197 2200 2217
rect 2220 2197 2240 2217
rect 2260 2197 2280 2217
rect 2300 2197 2320 2217
rect 2340 2197 2360 2217
rect 2380 2197 2400 2217
rect 2420 2197 2440 2217
rect 2460 2197 2480 2217
rect 2500 2197 2520 2217
rect 2540 2197 2560 2217
rect 2580 2197 2600 2217
rect 2620 2197 2640 2217
rect 2660 2197 2675 2217
rect 175 2182 2675 2197
rect 175 2135 2675 2150
rect 175 2115 200 2135
rect 220 2115 240 2135
rect 260 2115 280 2135
rect 300 2115 320 2135
rect 340 2115 360 2135
rect 380 2115 400 2135
rect 420 2115 440 2135
rect 460 2115 480 2135
rect 500 2115 520 2135
rect 540 2115 560 2135
rect 580 2115 600 2135
rect 620 2115 640 2135
rect 660 2115 680 2135
rect 700 2115 720 2135
rect 740 2115 760 2135
rect 780 2115 800 2135
rect 820 2115 840 2135
rect 860 2115 880 2135
rect 900 2115 920 2135
rect 940 2115 960 2135
rect 980 2115 1000 2135
rect 1020 2115 1040 2135
rect 1060 2115 1080 2135
rect 1100 2115 1120 2135
rect 1140 2115 1160 2135
rect 1180 2115 1200 2135
rect 1220 2115 1240 2135
rect 1260 2115 1280 2135
rect 1300 2115 1320 2135
rect 1340 2115 1360 2135
rect 1380 2115 1400 2135
rect 1420 2115 1440 2135
rect 1460 2115 1480 2135
rect 1500 2115 1520 2135
rect 1540 2115 1560 2135
rect 1580 2115 1600 2135
rect 1620 2115 1640 2135
rect 1660 2115 1680 2135
rect 1700 2115 1720 2135
rect 1740 2115 1760 2135
rect 1780 2115 1800 2135
rect 1820 2115 1840 2135
rect 1860 2115 1880 2135
rect 1900 2115 1920 2135
rect 1940 2115 1960 2135
rect 1980 2115 2000 2135
rect 2020 2115 2040 2135
rect 2060 2115 2080 2135
rect 2100 2115 2120 2135
rect 2140 2115 2160 2135
rect 2180 2115 2200 2135
rect 2220 2115 2240 2135
rect 2260 2115 2280 2135
rect 2300 2115 2320 2135
rect 2340 2115 2360 2135
rect 2380 2115 2400 2135
rect 2420 2115 2440 2135
rect 2460 2115 2480 2135
rect 2500 2115 2520 2135
rect 2540 2115 2560 2135
rect 2580 2115 2600 2135
rect 2620 2115 2640 2135
rect 2660 2115 2675 2135
rect 175 2100 2675 2115
rect 175 2053 2675 2068
rect 175 2033 200 2053
rect 220 2033 240 2053
rect 260 2033 280 2053
rect 300 2033 320 2053
rect 340 2033 360 2053
rect 380 2033 400 2053
rect 420 2033 440 2053
rect 460 2033 480 2053
rect 500 2033 520 2053
rect 540 2033 560 2053
rect 580 2033 600 2053
rect 620 2033 640 2053
rect 660 2033 680 2053
rect 700 2033 720 2053
rect 740 2033 760 2053
rect 780 2033 800 2053
rect 820 2033 840 2053
rect 860 2033 880 2053
rect 900 2033 920 2053
rect 940 2033 960 2053
rect 980 2033 1000 2053
rect 1020 2033 1040 2053
rect 1060 2033 1080 2053
rect 1100 2033 1120 2053
rect 1140 2033 1160 2053
rect 1180 2033 1200 2053
rect 1220 2033 1240 2053
rect 1260 2033 1280 2053
rect 1300 2033 1320 2053
rect 1340 2033 1360 2053
rect 1380 2033 1400 2053
rect 1420 2033 1440 2053
rect 1460 2033 1480 2053
rect 1500 2033 1520 2053
rect 1540 2033 1560 2053
rect 1580 2033 1600 2053
rect 1620 2033 1640 2053
rect 1660 2033 1680 2053
rect 1700 2033 1720 2053
rect 1740 2033 1760 2053
rect 1780 2033 1800 2053
rect 1820 2033 1840 2053
rect 1860 2033 1880 2053
rect 1900 2033 1920 2053
rect 1940 2033 1960 2053
rect 1980 2033 2000 2053
rect 2020 2033 2040 2053
rect 2060 2033 2080 2053
rect 2100 2033 2120 2053
rect 2140 2033 2160 2053
rect 2180 2033 2200 2053
rect 2220 2033 2240 2053
rect 2260 2033 2280 2053
rect 2300 2033 2320 2053
rect 2340 2033 2360 2053
rect 2380 2033 2400 2053
rect 2420 2033 2440 2053
rect 2460 2033 2480 2053
rect 2500 2033 2520 2053
rect 2540 2033 2560 2053
rect 2580 2033 2600 2053
rect 2620 2033 2640 2053
rect 2660 2033 2675 2053
rect 175 2018 2675 2033
rect 175 1971 2675 1986
rect 175 1951 200 1971
rect 220 1951 240 1971
rect 260 1951 280 1971
rect 300 1951 320 1971
rect 340 1951 360 1971
rect 380 1951 400 1971
rect 420 1951 440 1971
rect 460 1951 480 1971
rect 500 1951 520 1971
rect 540 1951 560 1971
rect 580 1951 600 1971
rect 620 1951 640 1971
rect 660 1951 680 1971
rect 700 1951 720 1971
rect 740 1951 760 1971
rect 780 1951 800 1971
rect 820 1951 840 1971
rect 860 1951 880 1971
rect 900 1951 920 1971
rect 940 1951 960 1971
rect 980 1951 1000 1971
rect 1020 1951 1040 1971
rect 1060 1951 1080 1971
rect 1100 1951 1120 1971
rect 1140 1951 1160 1971
rect 1180 1951 1200 1971
rect 1220 1951 1240 1971
rect 1260 1951 1280 1971
rect 1300 1951 1320 1971
rect 1340 1951 1360 1971
rect 1380 1951 1400 1971
rect 1420 1951 1440 1971
rect 1460 1951 1480 1971
rect 1500 1951 1520 1971
rect 1540 1951 1560 1971
rect 1580 1951 1600 1971
rect 1620 1951 1640 1971
rect 1660 1951 1680 1971
rect 1700 1951 1720 1971
rect 1740 1951 1760 1971
rect 1780 1951 1800 1971
rect 1820 1951 1840 1971
rect 1860 1951 1880 1971
rect 1900 1951 1920 1971
rect 1940 1951 1960 1971
rect 1980 1951 2000 1971
rect 2020 1951 2040 1971
rect 2060 1951 2080 1971
rect 2100 1951 2120 1971
rect 2140 1951 2160 1971
rect 2180 1951 2200 1971
rect 2220 1951 2240 1971
rect 2260 1951 2280 1971
rect 2300 1951 2320 1971
rect 2340 1951 2360 1971
rect 2380 1951 2400 1971
rect 2420 1951 2440 1971
rect 2460 1951 2480 1971
rect 2500 1951 2520 1971
rect 2540 1951 2560 1971
rect 2580 1951 2600 1971
rect 2620 1951 2640 1971
rect 2660 1951 2675 1971
rect 175 1936 2675 1951
rect 175 1889 2675 1904
rect 175 1869 200 1889
rect 220 1869 240 1889
rect 260 1869 280 1889
rect 300 1869 320 1889
rect 340 1869 360 1889
rect 380 1869 400 1889
rect 420 1869 440 1889
rect 460 1869 480 1889
rect 500 1869 520 1889
rect 540 1869 560 1889
rect 580 1869 600 1889
rect 620 1869 640 1889
rect 660 1869 680 1889
rect 700 1869 720 1889
rect 740 1869 760 1889
rect 780 1869 800 1889
rect 820 1869 840 1889
rect 860 1869 880 1889
rect 900 1869 920 1889
rect 940 1869 960 1889
rect 980 1869 1000 1889
rect 1020 1869 1040 1889
rect 1060 1869 1080 1889
rect 1100 1869 1120 1889
rect 1140 1869 1160 1889
rect 1180 1869 1200 1889
rect 1220 1869 1240 1889
rect 1260 1869 1280 1889
rect 1300 1869 1320 1889
rect 1340 1869 1360 1889
rect 1380 1869 1400 1889
rect 1420 1869 1440 1889
rect 1460 1869 1480 1889
rect 1500 1869 1520 1889
rect 1540 1869 1560 1889
rect 1580 1869 1600 1889
rect 1620 1869 1640 1889
rect 1660 1869 1680 1889
rect 1700 1869 1720 1889
rect 1740 1869 1760 1889
rect 1780 1869 1800 1889
rect 1820 1869 1840 1889
rect 1860 1869 1880 1889
rect 1900 1869 1920 1889
rect 1940 1869 1960 1889
rect 1980 1869 2000 1889
rect 2020 1869 2040 1889
rect 2060 1869 2080 1889
rect 2100 1869 2120 1889
rect 2140 1869 2160 1889
rect 2180 1869 2200 1889
rect 2220 1869 2240 1889
rect 2260 1869 2280 1889
rect 2300 1869 2320 1889
rect 2340 1869 2360 1889
rect 2380 1869 2400 1889
rect 2420 1869 2440 1889
rect 2460 1869 2480 1889
rect 2500 1869 2520 1889
rect 2540 1869 2560 1889
rect 2580 1869 2600 1889
rect 2620 1869 2640 1889
rect 2660 1869 2675 1889
rect 175 1854 2675 1869
rect 175 1807 2675 1822
rect 175 1787 200 1807
rect 220 1787 240 1807
rect 260 1787 280 1807
rect 300 1787 320 1807
rect 340 1787 360 1807
rect 380 1787 400 1807
rect 420 1787 440 1807
rect 460 1787 480 1807
rect 500 1787 520 1807
rect 540 1787 560 1807
rect 580 1787 600 1807
rect 620 1787 640 1807
rect 660 1787 680 1807
rect 700 1787 720 1807
rect 740 1787 760 1807
rect 780 1787 800 1807
rect 820 1787 840 1807
rect 860 1787 880 1807
rect 900 1787 920 1807
rect 940 1787 960 1807
rect 980 1787 1000 1807
rect 1020 1787 1040 1807
rect 1060 1787 1080 1807
rect 1100 1787 1120 1807
rect 1140 1787 1160 1807
rect 1180 1787 1200 1807
rect 1220 1787 1240 1807
rect 1260 1787 1280 1807
rect 1300 1787 1320 1807
rect 1340 1787 1360 1807
rect 1380 1787 1400 1807
rect 1420 1787 1440 1807
rect 1460 1787 1480 1807
rect 1500 1787 1520 1807
rect 1540 1787 1560 1807
rect 1580 1787 1600 1807
rect 1620 1787 1640 1807
rect 1660 1787 1680 1807
rect 1700 1787 1720 1807
rect 1740 1787 1760 1807
rect 1780 1787 1800 1807
rect 1820 1787 1840 1807
rect 1860 1787 1880 1807
rect 1900 1787 1920 1807
rect 1940 1787 1960 1807
rect 1980 1787 2000 1807
rect 2020 1787 2040 1807
rect 2060 1787 2080 1807
rect 2100 1787 2120 1807
rect 2140 1787 2160 1807
rect 2180 1787 2200 1807
rect 2220 1787 2240 1807
rect 2260 1787 2280 1807
rect 2300 1787 2320 1807
rect 2340 1787 2360 1807
rect 2380 1787 2400 1807
rect 2420 1787 2440 1807
rect 2460 1787 2480 1807
rect 2500 1787 2520 1807
rect 2540 1787 2560 1807
rect 2580 1787 2600 1807
rect 2620 1787 2640 1807
rect 2660 1787 2675 1807
rect 175 1772 2675 1787
rect 175 1725 2675 1740
rect 175 1705 200 1725
rect 220 1705 240 1725
rect 260 1705 280 1725
rect 300 1705 320 1725
rect 340 1705 360 1725
rect 380 1705 400 1725
rect 420 1705 440 1725
rect 460 1705 480 1725
rect 500 1705 520 1725
rect 540 1705 560 1725
rect 580 1705 600 1725
rect 620 1705 640 1725
rect 660 1705 680 1725
rect 700 1705 720 1725
rect 740 1705 760 1725
rect 780 1705 800 1725
rect 820 1705 840 1725
rect 860 1705 880 1725
rect 900 1705 920 1725
rect 940 1705 960 1725
rect 980 1705 1000 1725
rect 1020 1705 1040 1725
rect 1060 1705 1080 1725
rect 1100 1705 1120 1725
rect 1140 1705 1160 1725
rect 1180 1705 1200 1725
rect 1220 1705 1240 1725
rect 1260 1705 1280 1725
rect 1300 1705 1320 1725
rect 1340 1705 1360 1725
rect 1380 1705 1400 1725
rect 1420 1705 1440 1725
rect 1460 1705 1480 1725
rect 1500 1705 1520 1725
rect 1540 1705 1560 1725
rect 1580 1705 1600 1725
rect 1620 1705 1640 1725
rect 1660 1705 1680 1725
rect 1700 1705 1720 1725
rect 1740 1705 1760 1725
rect 1780 1705 1800 1725
rect 1820 1705 1840 1725
rect 1860 1705 1880 1725
rect 1900 1705 1920 1725
rect 1940 1705 1960 1725
rect 1980 1705 2000 1725
rect 2020 1705 2040 1725
rect 2060 1705 2080 1725
rect 2100 1705 2120 1725
rect 2140 1705 2160 1725
rect 2180 1705 2200 1725
rect 2220 1705 2240 1725
rect 2260 1705 2280 1725
rect 2300 1705 2320 1725
rect 2340 1705 2360 1725
rect 2380 1705 2400 1725
rect 2420 1705 2440 1725
rect 2460 1705 2480 1725
rect 2500 1705 2520 1725
rect 2540 1705 2560 1725
rect 2580 1705 2600 1725
rect 2620 1705 2640 1725
rect 2660 1705 2675 1725
rect 175 1690 2675 1705
rect 175 1643 2675 1658
rect 175 1623 200 1643
rect 220 1623 240 1643
rect 260 1623 280 1643
rect 300 1623 320 1643
rect 340 1623 360 1643
rect 380 1623 400 1643
rect 420 1623 440 1643
rect 460 1623 480 1643
rect 500 1623 520 1643
rect 540 1623 560 1643
rect 580 1623 600 1643
rect 620 1623 640 1643
rect 660 1623 680 1643
rect 700 1623 720 1643
rect 740 1623 760 1643
rect 780 1623 800 1643
rect 820 1623 840 1643
rect 860 1623 880 1643
rect 900 1623 920 1643
rect 940 1623 960 1643
rect 980 1623 1000 1643
rect 1020 1623 1040 1643
rect 1060 1623 1080 1643
rect 1100 1623 1120 1643
rect 1140 1623 1160 1643
rect 1180 1623 1200 1643
rect 1220 1623 1240 1643
rect 1260 1623 1280 1643
rect 1300 1623 1320 1643
rect 1340 1623 1360 1643
rect 1380 1623 1400 1643
rect 1420 1623 1440 1643
rect 1460 1623 1480 1643
rect 1500 1623 1520 1643
rect 1540 1623 1560 1643
rect 1580 1623 1600 1643
rect 1620 1623 1640 1643
rect 1660 1623 1680 1643
rect 1700 1623 1720 1643
rect 1740 1623 1760 1643
rect 1780 1623 1800 1643
rect 1820 1623 1840 1643
rect 1860 1623 1880 1643
rect 1900 1623 1920 1643
rect 1940 1623 1960 1643
rect 1980 1623 2000 1643
rect 2020 1623 2040 1643
rect 2060 1623 2080 1643
rect 2100 1623 2120 1643
rect 2140 1623 2160 1643
rect 2180 1623 2200 1643
rect 2220 1623 2240 1643
rect 2260 1623 2280 1643
rect 2300 1623 2320 1643
rect 2340 1623 2360 1643
rect 2380 1623 2400 1643
rect 2420 1623 2440 1643
rect 2460 1623 2480 1643
rect 2500 1623 2520 1643
rect 2540 1623 2560 1643
rect 2580 1623 2600 1643
rect 2620 1623 2640 1643
rect 2660 1623 2675 1643
rect 175 1608 2675 1623
rect 175 1561 2675 1576
rect 175 1541 200 1561
rect 220 1541 240 1561
rect 260 1541 280 1561
rect 300 1541 320 1561
rect 340 1541 360 1561
rect 380 1541 400 1561
rect 420 1541 440 1561
rect 460 1541 480 1561
rect 500 1541 520 1561
rect 540 1541 560 1561
rect 580 1541 600 1561
rect 620 1541 640 1561
rect 660 1541 680 1561
rect 700 1541 720 1561
rect 740 1541 760 1561
rect 780 1541 800 1561
rect 820 1541 840 1561
rect 860 1541 880 1561
rect 900 1541 920 1561
rect 940 1541 960 1561
rect 980 1541 1000 1561
rect 1020 1541 1040 1561
rect 1060 1541 1080 1561
rect 1100 1541 1120 1561
rect 1140 1541 1160 1561
rect 1180 1541 1200 1561
rect 1220 1541 1240 1561
rect 1260 1541 1280 1561
rect 1300 1541 1320 1561
rect 1340 1541 1360 1561
rect 1380 1541 1400 1561
rect 1420 1541 1440 1561
rect 1460 1541 1480 1561
rect 1500 1541 1520 1561
rect 1540 1541 1560 1561
rect 1580 1541 1600 1561
rect 1620 1541 1640 1561
rect 1660 1541 1680 1561
rect 1700 1541 1720 1561
rect 1740 1541 1760 1561
rect 1780 1541 1800 1561
rect 1820 1541 1840 1561
rect 1860 1541 1880 1561
rect 1900 1541 1920 1561
rect 1940 1541 1960 1561
rect 1980 1541 2000 1561
rect 2020 1541 2040 1561
rect 2060 1541 2080 1561
rect 2100 1541 2120 1561
rect 2140 1541 2160 1561
rect 2180 1541 2200 1561
rect 2220 1541 2240 1561
rect 2260 1541 2280 1561
rect 2300 1541 2320 1561
rect 2340 1541 2360 1561
rect 2380 1541 2400 1561
rect 2420 1541 2440 1561
rect 2460 1541 2480 1561
rect 2500 1541 2520 1561
rect 2540 1541 2560 1561
rect 2580 1541 2600 1561
rect 2620 1541 2640 1561
rect 2660 1541 2675 1561
rect 175 1526 2675 1541
rect 175 1479 2675 1494
rect 175 1459 200 1479
rect 220 1459 240 1479
rect 260 1459 280 1479
rect 300 1459 320 1479
rect 340 1459 360 1479
rect 380 1459 400 1479
rect 420 1459 440 1479
rect 460 1459 480 1479
rect 500 1459 520 1479
rect 540 1459 560 1479
rect 580 1459 600 1479
rect 620 1459 640 1479
rect 660 1459 680 1479
rect 700 1459 720 1479
rect 740 1459 760 1479
rect 780 1459 800 1479
rect 820 1459 840 1479
rect 860 1459 880 1479
rect 900 1459 920 1479
rect 940 1459 960 1479
rect 980 1459 1000 1479
rect 1020 1459 1040 1479
rect 1060 1459 1080 1479
rect 1100 1459 1120 1479
rect 1140 1459 1160 1479
rect 1180 1459 1200 1479
rect 1220 1459 1240 1479
rect 1260 1459 1280 1479
rect 1300 1459 1320 1479
rect 1340 1459 1360 1479
rect 1380 1459 1400 1479
rect 1420 1459 1440 1479
rect 1460 1459 1480 1479
rect 1500 1459 1520 1479
rect 1540 1459 1560 1479
rect 1580 1459 1600 1479
rect 1620 1459 1640 1479
rect 1660 1459 1680 1479
rect 1700 1459 1720 1479
rect 1740 1459 1760 1479
rect 1780 1459 1800 1479
rect 1820 1459 1840 1479
rect 1860 1459 1880 1479
rect 1900 1459 1920 1479
rect 1940 1459 1960 1479
rect 1980 1459 2000 1479
rect 2020 1459 2040 1479
rect 2060 1459 2080 1479
rect 2100 1459 2120 1479
rect 2140 1459 2160 1479
rect 2180 1459 2200 1479
rect 2220 1459 2240 1479
rect 2260 1459 2280 1479
rect 2300 1459 2320 1479
rect 2340 1459 2360 1479
rect 2380 1459 2400 1479
rect 2420 1459 2440 1479
rect 2460 1459 2480 1479
rect 2500 1459 2520 1479
rect 2540 1459 2560 1479
rect 2580 1459 2600 1479
rect 2620 1459 2640 1479
rect 2660 1459 2675 1479
rect 175 1444 2675 1459
rect 175 1397 2675 1412
rect 175 1377 200 1397
rect 220 1377 240 1397
rect 260 1377 280 1397
rect 300 1377 320 1397
rect 340 1377 360 1397
rect 380 1377 400 1397
rect 420 1377 440 1397
rect 460 1377 480 1397
rect 500 1377 520 1397
rect 540 1377 560 1397
rect 580 1377 600 1397
rect 620 1377 640 1397
rect 660 1377 680 1397
rect 700 1377 720 1397
rect 740 1377 760 1397
rect 780 1377 800 1397
rect 820 1377 840 1397
rect 860 1377 880 1397
rect 900 1377 920 1397
rect 940 1377 960 1397
rect 980 1377 1000 1397
rect 1020 1377 1040 1397
rect 1060 1377 1080 1397
rect 1100 1377 1120 1397
rect 1140 1377 1160 1397
rect 1180 1377 1200 1397
rect 1220 1377 1240 1397
rect 1260 1377 1280 1397
rect 1300 1377 1320 1397
rect 1340 1377 1360 1397
rect 1380 1377 1400 1397
rect 1420 1377 1440 1397
rect 1460 1377 1480 1397
rect 1500 1377 1520 1397
rect 1540 1377 1560 1397
rect 1580 1377 1600 1397
rect 1620 1377 1640 1397
rect 1660 1377 1680 1397
rect 1700 1377 1720 1397
rect 1740 1377 1760 1397
rect 1780 1377 1800 1397
rect 1820 1377 1840 1397
rect 1860 1377 1880 1397
rect 1900 1377 1920 1397
rect 1940 1377 1960 1397
rect 1980 1377 2000 1397
rect 2020 1377 2040 1397
rect 2060 1377 2080 1397
rect 2100 1377 2120 1397
rect 2140 1377 2160 1397
rect 2180 1377 2200 1397
rect 2220 1377 2240 1397
rect 2260 1377 2280 1397
rect 2300 1377 2320 1397
rect 2340 1377 2360 1397
rect 2380 1377 2400 1397
rect 2420 1377 2440 1397
rect 2460 1377 2480 1397
rect 2500 1377 2520 1397
rect 2540 1377 2560 1397
rect 2580 1377 2600 1397
rect 2620 1377 2640 1397
rect 2660 1377 2675 1397
rect 175 1362 2675 1377
rect 175 1315 2675 1330
rect 175 1295 200 1315
rect 220 1295 240 1315
rect 260 1295 280 1315
rect 300 1295 320 1315
rect 340 1295 360 1315
rect 380 1295 400 1315
rect 420 1295 440 1315
rect 460 1295 480 1315
rect 500 1295 520 1315
rect 540 1295 560 1315
rect 580 1295 600 1315
rect 620 1295 640 1315
rect 660 1295 680 1315
rect 700 1295 720 1315
rect 740 1295 760 1315
rect 780 1295 800 1315
rect 820 1295 840 1315
rect 860 1295 880 1315
rect 900 1295 920 1315
rect 940 1295 960 1315
rect 980 1295 1000 1315
rect 1020 1295 1040 1315
rect 1060 1295 1080 1315
rect 1100 1295 1120 1315
rect 1140 1295 1160 1315
rect 1180 1295 1200 1315
rect 1220 1295 1240 1315
rect 1260 1295 1280 1315
rect 1300 1295 1320 1315
rect 1340 1295 1360 1315
rect 1380 1295 1400 1315
rect 1420 1295 1440 1315
rect 1460 1295 1480 1315
rect 1500 1295 1520 1315
rect 1540 1295 1560 1315
rect 1580 1295 1600 1315
rect 1620 1295 1640 1315
rect 1660 1295 1680 1315
rect 1700 1295 1720 1315
rect 1740 1295 1760 1315
rect 1780 1295 1800 1315
rect 1820 1295 1840 1315
rect 1860 1295 1880 1315
rect 1900 1295 1920 1315
rect 1940 1295 1960 1315
rect 1980 1295 2000 1315
rect 2020 1295 2040 1315
rect 2060 1295 2080 1315
rect 2100 1295 2120 1315
rect 2140 1295 2160 1315
rect 2180 1295 2200 1315
rect 2220 1295 2240 1315
rect 2260 1295 2280 1315
rect 2300 1295 2320 1315
rect 2340 1295 2360 1315
rect 2380 1295 2400 1315
rect 2420 1295 2440 1315
rect 2460 1295 2480 1315
rect 2500 1295 2520 1315
rect 2540 1295 2560 1315
rect 2580 1295 2600 1315
rect 2620 1295 2640 1315
rect 2660 1295 2675 1315
rect 175 1280 2675 1295
rect 175 1233 2675 1248
rect 175 1213 200 1233
rect 220 1213 240 1233
rect 260 1213 280 1233
rect 300 1213 320 1233
rect 340 1213 360 1233
rect 380 1213 400 1233
rect 420 1213 440 1233
rect 460 1213 480 1233
rect 500 1213 520 1233
rect 540 1213 560 1233
rect 580 1213 600 1233
rect 620 1213 640 1233
rect 660 1213 680 1233
rect 700 1213 720 1233
rect 740 1213 760 1233
rect 780 1213 800 1233
rect 820 1213 840 1233
rect 860 1213 880 1233
rect 900 1213 920 1233
rect 940 1213 960 1233
rect 980 1213 1000 1233
rect 1020 1213 1040 1233
rect 1060 1213 1080 1233
rect 1100 1213 1120 1233
rect 1140 1213 1160 1233
rect 1180 1213 1200 1233
rect 1220 1213 1240 1233
rect 1260 1213 1280 1233
rect 1300 1213 1320 1233
rect 1340 1213 1360 1233
rect 1380 1213 1400 1233
rect 1420 1213 1440 1233
rect 1460 1213 1480 1233
rect 1500 1213 1520 1233
rect 1540 1213 1560 1233
rect 1580 1213 1600 1233
rect 1620 1213 1640 1233
rect 1660 1213 1680 1233
rect 1700 1213 1720 1233
rect 1740 1213 1760 1233
rect 1780 1213 1800 1233
rect 1820 1213 1840 1233
rect 1860 1213 1880 1233
rect 1900 1213 1920 1233
rect 1940 1213 1960 1233
rect 1980 1213 2000 1233
rect 2020 1213 2040 1233
rect 2060 1213 2080 1233
rect 2100 1213 2120 1233
rect 2140 1213 2160 1233
rect 2180 1213 2200 1233
rect 2220 1213 2240 1233
rect 2260 1213 2280 1233
rect 2300 1213 2320 1233
rect 2340 1213 2360 1233
rect 2380 1213 2400 1233
rect 2420 1213 2440 1233
rect 2460 1213 2480 1233
rect 2500 1213 2520 1233
rect 2540 1213 2560 1233
rect 2580 1213 2600 1233
rect 2620 1213 2640 1233
rect 2660 1213 2675 1233
rect 175 1198 2675 1213
rect 175 1151 2675 1166
rect 175 1131 200 1151
rect 220 1131 240 1151
rect 260 1131 280 1151
rect 300 1131 320 1151
rect 340 1131 360 1151
rect 380 1131 400 1151
rect 420 1131 440 1151
rect 460 1131 480 1151
rect 500 1131 520 1151
rect 540 1131 560 1151
rect 580 1131 600 1151
rect 620 1131 640 1151
rect 660 1131 680 1151
rect 700 1131 720 1151
rect 740 1131 760 1151
rect 780 1131 800 1151
rect 820 1131 840 1151
rect 860 1131 880 1151
rect 900 1131 920 1151
rect 940 1131 960 1151
rect 980 1131 1000 1151
rect 1020 1131 1040 1151
rect 1060 1131 1080 1151
rect 1100 1131 1120 1151
rect 1140 1131 1160 1151
rect 1180 1131 1200 1151
rect 1220 1131 1240 1151
rect 1260 1131 1280 1151
rect 1300 1131 1320 1151
rect 1340 1131 1360 1151
rect 1380 1131 1400 1151
rect 1420 1131 1440 1151
rect 1460 1131 1480 1151
rect 1500 1131 1520 1151
rect 1540 1131 1560 1151
rect 1580 1131 1600 1151
rect 1620 1131 1640 1151
rect 1660 1131 1680 1151
rect 1700 1131 1720 1151
rect 1740 1131 1760 1151
rect 1780 1131 1800 1151
rect 1820 1131 1840 1151
rect 1860 1131 1880 1151
rect 1900 1131 1920 1151
rect 1940 1131 1960 1151
rect 1980 1131 2000 1151
rect 2020 1131 2040 1151
rect 2060 1131 2080 1151
rect 2100 1131 2120 1151
rect 2140 1131 2160 1151
rect 2180 1131 2200 1151
rect 2220 1131 2240 1151
rect 2260 1131 2280 1151
rect 2300 1131 2320 1151
rect 2340 1131 2360 1151
rect 2380 1131 2400 1151
rect 2420 1131 2440 1151
rect 2460 1131 2480 1151
rect 2500 1131 2520 1151
rect 2540 1131 2560 1151
rect 2580 1131 2600 1151
rect 2620 1131 2640 1151
rect 2660 1131 2675 1151
rect 175 1116 2675 1131
rect 175 1069 2675 1084
rect 175 1049 200 1069
rect 220 1049 240 1069
rect 260 1049 280 1069
rect 300 1049 320 1069
rect 340 1049 360 1069
rect 380 1049 400 1069
rect 420 1049 440 1069
rect 460 1049 480 1069
rect 500 1049 520 1069
rect 540 1049 560 1069
rect 580 1049 600 1069
rect 620 1049 640 1069
rect 660 1049 680 1069
rect 700 1049 720 1069
rect 740 1049 760 1069
rect 780 1049 800 1069
rect 820 1049 840 1069
rect 860 1049 880 1069
rect 900 1049 920 1069
rect 940 1049 960 1069
rect 980 1049 1000 1069
rect 1020 1049 1040 1069
rect 1060 1049 1080 1069
rect 1100 1049 1120 1069
rect 1140 1049 1160 1069
rect 1180 1049 1200 1069
rect 1220 1049 1240 1069
rect 1260 1049 1280 1069
rect 1300 1049 1320 1069
rect 1340 1049 1360 1069
rect 1380 1049 1400 1069
rect 1420 1049 1440 1069
rect 1460 1049 1480 1069
rect 1500 1049 1520 1069
rect 1540 1049 1560 1069
rect 1580 1049 1600 1069
rect 1620 1049 1640 1069
rect 1660 1049 1680 1069
rect 1700 1049 1720 1069
rect 1740 1049 1760 1069
rect 1780 1049 1800 1069
rect 1820 1049 1840 1069
rect 1860 1049 1880 1069
rect 1900 1049 1920 1069
rect 1940 1049 1960 1069
rect 1980 1049 2000 1069
rect 2020 1049 2040 1069
rect 2060 1049 2080 1069
rect 2100 1049 2120 1069
rect 2140 1049 2160 1069
rect 2180 1049 2200 1069
rect 2220 1049 2240 1069
rect 2260 1049 2280 1069
rect 2300 1049 2320 1069
rect 2340 1049 2360 1069
rect 2380 1049 2400 1069
rect 2420 1049 2440 1069
rect 2460 1049 2480 1069
rect 2500 1049 2520 1069
rect 2540 1049 2560 1069
rect 2580 1049 2600 1069
rect 2620 1049 2640 1069
rect 2660 1049 2675 1069
rect 175 1034 2675 1049
rect 175 987 2675 1002
rect 175 967 200 987
rect 220 967 240 987
rect 260 967 280 987
rect 300 967 320 987
rect 340 967 360 987
rect 380 967 400 987
rect 420 967 440 987
rect 460 967 480 987
rect 500 967 520 987
rect 540 967 560 987
rect 580 967 600 987
rect 620 967 640 987
rect 660 967 680 987
rect 700 967 720 987
rect 740 967 760 987
rect 780 967 800 987
rect 820 967 840 987
rect 860 967 880 987
rect 900 967 920 987
rect 940 967 960 987
rect 980 967 1000 987
rect 1020 967 1040 987
rect 1060 967 1080 987
rect 1100 967 1120 987
rect 1140 967 1160 987
rect 1180 967 1200 987
rect 1220 967 1240 987
rect 1260 967 1280 987
rect 1300 967 1320 987
rect 1340 967 1360 987
rect 1380 967 1400 987
rect 1420 967 1440 987
rect 1460 967 1480 987
rect 1500 967 1520 987
rect 1540 967 1560 987
rect 1580 967 1600 987
rect 1620 967 1640 987
rect 1660 967 1680 987
rect 1700 967 1720 987
rect 1740 967 1760 987
rect 1780 967 1800 987
rect 1820 967 1840 987
rect 1860 967 1880 987
rect 1900 967 1920 987
rect 1940 967 1960 987
rect 1980 967 2000 987
rect 2020 967 2040 987
rect 2060 967 2080 987
rect 2100 967 2120 987
rect 2140 967 2160 987
rect 2180 967 2200 987
rect 2220 967 2240 987
rect 2260 967 2280 987
rect 2300 967 2320 987
rect 2340 967 2360 987
rect 2380 967 2400 987
rect 2420 967 2440 987
rect 2460 967 2480 987
rect 2500 967 2520 987
rect 2540 967 2560 987
rect 2580 967 2600 987
rect 2620 967 2640 987
rect 2660 967 2675 987
rect 175 952 2675 967
rect 175 905 2675 920
rect 175 885 200 905
rect 220 885 240 905
rect 260 885 280 905
rect 300 885 320 905
rect 340 885 360 905
rect 380 885 400 905
rect 420 885 440 905
rect 460 885 480 905
rect 500 885 520 905
rect 540 885 560 905
rect 580 885 600 905
rect 620 885 640 905
rect 660 885 680 905
rect 700 885 720 905
rect 740 885 760 905
rect 780 885 800 905
rect 820 885 840 905
rect 860 885 880 905
rect 900 885 920 905
rect 940 885 960 905
rect 980 885 1000 905
rect 1020 885 1040 905
rect 1060 885 1080 905
rect 1100 885 1120 905
rect 1140 885 1160 905
rect 1180 885 1200 905
rect 1220 885 1240 905
rect 1260 885 1280 905
rect 1300 885 1320 905
rect 1340 885 1360 905
rect 1380 885 1400 905
rect 1420 885 1440 905
rect 1460 885 1480 905
rect 1500 885 1520 905
rect 1540 885 1560 905
rect 1580 885 1600 905
rect 1620 885 1640 905
rect 1660 885 1680 905
rect 1700 885 1720 905
rect 1740 885 1760 905
rect 1780 885 1800 905
rect 1820 885 1840 905
rect 1860 885 1880 905
rect 1900 885 1920 905
rect 1940 885 1960 905
rect 1980 885 2000 905
rect 2020 885 2040 905
rect 2060 885 2080 905
rect 2100 885 2120 905
rect 2140 885 2160 905
rect 2180 885 2200 905
rect 2220 885 2240 905
rect 2260 885 2280 905
rect 2300 885 2320 905
rect 2340 885 2360 905
rect 2380 885 2400 905
rect 2420 885 2440 905
rect 2460 885 2480 905
rect 2500 885 2520 905
rect 2540 885 2560 905
rect 2580 885 2600 905
rect 2620 885 2640 905
rect 2660 885 2675 905
rect 175 870 2675 885
rect 175 823 2675 838
rect 175 803 200 823
rect 220 803 240 823
rect 260 803 280 823
rect 300 803 320 823
rect 340 803 360 823
rect 380 803 400 823
rect 420 803 440 823
rect 460 803 480 823
rect 500 803 520 823
rect 540 803 560 823
rect 580 803 600 823
rect 620 803 640 823
rect 660 803 680 823
rect 700 803 720 823
rect 740 803 760 823
rect 780 803 800 823
rect 820 803 840 823
rect 860 803 880 823
rect 900 803 920 823
rect 940 803 960 823
rect 980 803 1000 823
rect 1020 803 1040 823
rect 1060 803 1080 823
rect 1100 803 1120 823
rect 1140 803 1160 823
rect 1180 803 1200 823
rect 1220 803 1240 823
rect 1260 803 1280 823
rect 1300 803 1320 823
rect 1340 803 1360 823
rect 1380 803 1400 823
rect 1420 803 1440 823
rect 1460 803 1480 823
rect 1500 803 1520 823
rect 1540 803 1560 823
rect 1580 803 1600 823
rect 1620 803 1640 823
rect 1660 803 1680 823
rect 1700 803 1720 823
rect 1740 803 1760 823
rect 1780 803 1800 823
rect 1820 803 1840 823
rect 1860 803 1880 823
rect 1900 803 1920 823
rect 1940 803 1960 823
rect 1980 803 2000 823
rect 2020 803 2040 823
rect 2060 803 2080 823
rect 2100 803 2120 823
rect 2140 803 2160 823
rect 2180 803 2200 823
rect 2220 803 2240 823
rect 2260 803 2280 823
rect 2300 803 2320 823
rect 2340 803 2360 823
rect 2380 803 2400 823
rect 2420 803 2440 823
rect 2460 803 2480 823
rect 2500 803 2520 823
rect 2540 803 2560 823
rect 2580 803 2600 823
rect 2620 803 2640 823
rect 2660 803 2675 823
rect 175 788 2675 803
rect 175 741 2675 756
rect 175 721 200 741
rect 220 721 240 741
rect 260 721 280 741
rect 300 721 320 741
rect 340 721 360 741
rect 380 721 400 741
rect 420 721 440 741
rect 460 721 480 741
rect 500 721 520 741
rect 540 721 560 741
rect 580 721 600 741
rect 620 721 640 741
rect 660 721 680 741
rect 700 721 720 741
rect 740 721 760 741
rect 780 721 800 741
rect 820 721 840 741
rect 860 721 880 741
rect 900 721 920 741
rect 940 721 960 741
rect 980 721 1000 741
rect 1020 721 1040 741
rect 1060 721 1080 741
rect 1100 721 1120 741
rect 1140 721 1160 741
rect 1180 721 1200 741
rect 1220 721 1240 741
rect 1260 721 1280 741
rect 1300 721 1320 741
rect 1340 721 1360 741
rect 1380 721 1400 741
rect 1420 721 1440 741
rect 1460 721 1480 741
rect 1500 721 1520 741
rect 1540 721 1560 741
rect 1580 721 1600 741
rect 1620 721 1640 741
rect 1660 721 1680 741
rect 1700 721 1720 741
rect 1740 721 1760 741
rect 1780 721 1800 741
rect 1820 721 1840 741
rect 1860 721 1880 741
rect 1900 721 1920 741
rect 1940 721 1960 741
rect 1980 721 2000 741
rect 2020 721 2040 741
rect 2060 721 2080 741
rect 2100 721 2120 741
rect 2140 721 2160 741
rect 2180 721 2200 741
rect 2220 721 2240 741
rect 2260 721 2280 741
rect 2300 721 2320 741
rect 2340 721 2360 741
rect 2380 721 2400 741
rect 2420 721 2440 741
rect 2460 721 2480 741
rect 2500 721 2520 741
rect 2540 721 2560 741
rect 2580 721 2600 741
rect 2620 721 2640 741
rect 2660 721 2675 741
rect 175 706 2675 721
rect 175 659 2675 674
rect 175 639 200 659
rect 220 639 240 659
rect 260 639 280 659
rect 300 639 320 659
rect 340 639 360 659
rect 380 639 400 659
rect 420 639 440 659
rect 460 639 480 659
rect 500 639 520 659
rect 540 639 560 659
rect 580 639 600 659
rect 620 639 640 659
rect 660 639 680 659
rect 700 639 720 659
rect 740 639 760 659
rect 780 639 800 659
rect 820 639 840 659
rect 860 639 880 659
rect 900 639 920 659
rect 940 639 960 659
rect 980 639 1000 659
rect 1020 639 1040 659
rect 1060 639 1080 659
rect 1100 639 1120 659
rect 1140 639 1160 659
rect 1180 639 1200 659
rect 1220 639 1240 659
rect 1260 639 1280 659
rect 1300 639 1320 659
rect 1340 639 1360 659
rect 1380 639 1400 659
rect 1420 639 1440 659
rect 1460 639 1480 659
rect 1500 639 1520 659
rect 1540 639 1560 659
rect 1580 639 1600 659
rect 1620 639 1640 659
rect 1660 639 1680 659
rect 1700 639 1720 659
rect 1740 639 1760 659
rect 1780 639 1800 659
rect 1820 639 1840 659
rect 1860 639 1880 659
rect 1900 639 1920 659
rect 1940 639 1960 659
rect 1980 639 2000 659
rect 2020 639 2040 659
rect 2060 639 2080 659
rect 2100 639 2120 659
rect 2140 639 2160 659
rect 2180 639 2200 659
rect 2220 639 2240 659
rect 2260 639 2280 659
rect 2300 639 2320 659
rect 2340 639 2360 659
rect 2380 639 2400 659
rect 2420 639 2440 659
rect 2460 639 2480 659
rect 2500 639 2520 659
rect 2540 639 2560 659
rect 2580 639 2600 659
rect 2620 639 2640 659
rect 2660 639 2675 659
rect 175 624 2675 639
rect 175 577 2675 592
rect 175 557 200 577
rect 220 557 240 577
rect 260 557 280 577
rect 300 557 320 577
rect 340 557 360 577
rect 380 557 400 577
rect 420 557 440 577
rect 460 557 480 577
rect 500 557 520 577
rect 540 557 560 577
rect 580 557 600 577
rect 620 557 640 577
rect 660 557 680 577
rect 700 557 720 577
rect 740 557 760 577
rect 780 557 800 577
rect 820 557 840 577
rect 860 557 880 577
rect 900 557 920 577
rect 940 557 960 577
rect 980 557 1000 577
rect 1020 557 1040 577
rect 1060 557 1080 577
rect 1100 557 1120 577
rect 1140 557 1160 577
rect 1180 557 1200 577
rect 1220 557 1240 577
rect 1260 557 1280 577
rect 1300 557 1320 577
rect 1340 557 1360 577
rect 1380 557 1400 577
rect 1420 557 1440 577
rect 1460 557 1480 577
rect 1500 557 1520 577
rect 1540 557 1560 577
rect 1580 557 1600 577
rect 1620 557 1640 577
rect 1660 557 1680 577
rect 1700 557 1720 577
rect 1740 557 1760 577
rect 1780 557 1800 577
rect 1820 557 1840 577
rect 1860 557 1880 577
rect 1900 557 1920 577
rect 1940 557 1960 577
rect 1980 557 2000 577
rect 2020 557 2040 577
rect 2060 557 2080 577
rect 2100 557 2120 577
rect 2140 557 2160 577
rect 2180 557 2200 577
rect 2220 557 2240 577
rect 2260 557 2280 577
rect 2300 557 2320 577
rect 2340 557 2360 577
rect 2380 557 2400 577
rect 2420 557 2440 577
rect 2460 557 2480 577
rect 2500 557 2520 577
rect 2540 557 2560 577
rect 2580 557 2600 577
rect 2620 557 2640 577
rect 2660 557 2675 577
rect 175 542 2675 557
rect 175 495 2675 510
rect 175 475 200 495
rect 220 475 240 495
rect 260 475 280 495
rect 300 475 320 495
rect 340 475 360 495
rect 380 475 400 495
rect 420 475 440 495
rect 460 475 480 495
rect 500 475 520 495
rect 540 475 560 495
rect 580 475 600 495
rect 620 475 640 495
rect 660 475 680 495
rect 700 475 720 495
rect 740 475 760 495
rect 780 475 800 495
rect 820 475 840 495
rect 860 475 880 495
rect 900 475 920 495
rect 940 475 960 495
rect 980 475 1000 495
rect 1020 475 1040 495
rect 1060 475 1080 495
rect 1100 475 1120 495
rect 1140 475 1160 495
rect 1180 475 1200 495
rect 1220 475 1240 495
rect 1260 475 1280 495
rect 1300 475 1320 495
rect 1340 475 1360 495
rect 1380 475 1400 495
rect 1420 475 1440 495
rect 1460 475 1480 495
rect 1500 475 1520 495
rect 1540 475 1560 495
rect 1580 475 1600 495
rect 1620 475 1640 495
rect 1660 475 1680 495
rect 1700 475 1720 495
rect 1740 475 1760 495
rect 1780 475 1800 495
rect 1820 475 1840 495
rect 1860 475 1880 495
rect 1900 475 1920 495
rect 1940 475 1960 495
rect 1980 475 2000 495
rect 2020 475 2040 495
rect 2060 475 2080 495
rect 2100 475 2120 495
rect 2140 475 2160 495
rect 2180 475 2200 495
rect 2220 475 2240 495
rect 2260 475 2280 495
rect 2300 475 2320 495
rect 2340 475 2360 495
rect 2380 475 2400 495
rect 2420 475 2440 495
rect 2460 475 2480 495
rect 2500 475 2520 495
rect 2540 475 2560 495
rect 2580 475 2600 495
rect 2620 475 2640 495
rect 2660 475 2675 495
rect 175 460 2675 475
rect 175 413 2675 428
rect 175 393 200 413
rect 220 393 240 413
rect 260 393 280 413
rect 300 393 320 413
rect 340 393 360 413
rect 380 393 400 413
rect 420 393 440 413
rect 460 393 480 413
rect 500 393 520 413
rect 540 393 560 413
rect 580 393 600 413
rect 620 393 640 413
rect 660 393 680 413
rect 700 393 720 413
rect 740 393 760 413
rect 780 393 800 413
rect 820 393 840 413
rect 860 393 880 413
rect 900 393 920 413
rect 940 393 960 413
rect 980 393 1000 413
rect 1020 393 1040 413
rect 1060 393 1080 413
rect 1100 393 1120 413
rect 1140 393 1160 413
rect 1180 393 1200 413
rect 1220 393 1240 413
rect 1260 393 1280 413
rect 1300 393 1320 413
rect 1340 393 1360 413
rect 1380 393 1400 413
rect 1420 393 1440 413
rect 1460 393 1480 413
rect 1500 393 1520 413
rect 1540 393 1560 413
rect 1580 393 1600 413
rect 1620 393 1640 413
rect 1660 393 1680 413
rect 1700 393 1720 413
rect 1740 393 1760 413
rect 1780 393 1800 413
rect 1820 393 1840 413
rect 1860 393 1880 413
rect 1900 393 1920 413
rect 1940 393 1960 413
rect 1980 393 2000 413
rect 2020 393 2040 413
rect 2060 393 2080 413
rect 2100 393 2120 413
rect 2140 393 2160 413
rect 2180 393 2200 413
rect 2220 393 2240 413
rect 2260 393 2280 413
rect 2300 393 2320 413
rect 2340 393 2360 413
rect 2380 393 2400 413
rect 2420 393 2440 413
rect 2460 393 2480 413
rect 2500 393 2520 413
rect 2540 393 2560 413
rect 2580 393 2600 413
rect 2620 393 2640 413
rect 2660 393 2675 413
rect 175 378 2675 393
rect 175 331 2675 346
rect 175 311 200 331
rect 220 311 240 331
rect 260 311 280 331
rect 300 311 320 331
rect 340 311 360 331
rect 380 311 400 331
rect 420 311 440 331
rect 460 311 480 331
rect 500 311 520 331
rect 540 311 560 331
rect 580 311 600 331
rect 620 311 640 331
rect 660 311 680 331
rect 700 311 720 331
rect 740 311 760 331
rect 780 311 800 331
rect 820 311 840 331
rect 860 311 880 331
rect 900 311 920 331
rect 940 311 960 331
rect 980 311 1000 331
rect 1020 311 1040 331
rect 1060 311 1080 331
rect 1100 311 1120 331
rect 1140 311 1160 331
rect 1180 311 1200 331
rect 1220 311 1240 331
rect 1260 311 1280 331
rect 1300 311 1320 331
rect 1340 311 1360 331
rect 1380 311 1400 331
rect 1420 311 1440 331
rect 1460 311 1480 331
rect 1500 311 1520 331
rect 1540 311 1560 331
rect 1580 311 1600 331
rect 1620 311 1640 331
rect 1660 311 1680 331
rect 1700 311 1720 331
rect 1740 311 1760 331
rect 1780 311 1800 331
rect 1820 311 1840 331
rect 1860 311 1880 331
rect 1900 311 1920 331
rect 1940 311 1960 331
rect 1980 311 2000 331
rect 2020 311 2040 331
rect 2060 311 2080 331
rect 2100 311 2120 331
rect 2140 311 2160 331
rect 2180 311 2200 331
rect 2220 311 2240 331
rect 2260 311 2280 331
rect 2300 311 2320 331
rect 2340 311 2360 331
rect 2380 311 2400 331
rect 2420 311 2440 331
rect 2460 311 2480 331
rect 2500 311 2520 331
rect 2540 311 2560 331
rect 2580 311 2600 331
rect 2620 311 2640 331
rect 2660 311 2675 331
rect 175 296 2675 311
rect 175 249 2675 264
rect 175 229 200 249
rect 220 229 240 249
rect 260 229 280 249
rect 300 229 320 249
rect 340 229 360 249
rect 380 229 400 249
rect 420 229 440 249
rect 460 229 480 249
rect 500 229 520 249
rect 540 229 560 249
rect 580 229 600 249
rect 620 229 640 249
rect 660 229 680 249
rect 700 229 720 249
rect 740 229 760 249
rect 780 229 800 249
rect 820 229 840 249
rect 860 229 880 249
rect 900 229 920 249
rect 940 229 960 249
rect 980 229 1000 249
rect 1020 229 1040 249
rect 1060 229 1080 249
rect 1100 229 1120 249
rect 1140 229 1160 249
rect 1180 229 1200 249
rect 1220 229 1240 249
rect 1260 229 1280 249
rect 1300 229 1320 249
rect 1340 229 1360 249
rect 1380 229 1400 249
rect 1420 229 1440 249
rect 1460 229 1480 249
rect 1500 229 1520 249
rect 1540 229 1560 249
rect 1580 229 1600 249
rect 1620 229 1640 249
rect 1660 229 1680 249
rect 1700 229 1720 249
rect 1740 229 1760 249
rect 1780 229 1800 249
rect 1820 229 1840 249
rect 1860 229 1880 249
rect 1900 229 1920 249
rect 1940 229 1960 249
rect 1980 229 2000 249
rect 2020 229 2040 249
rect 2060 229 2080 249
rect 2100 229 2120 249
rect 2140 229 2160 249
rect 2180 229 2200 249
rect 2220 229 2240 249
rect 2260 229 2280 249
rect 2300 229 2320 249
rect 2340 229 2360 249
rect 2380 229 2400 249
rect 2420 229 2440 249
rect 2460 229 2480 249
rect 2500 229 2520 249
rect 2540 229 2560 249
rect 2580 229 2600 249
rect 2620 229 2640 249
rect 2660 229 2675 249
rect 175 214 2675 229
rect 175 167 2675 182
rect 175 147 200 167
rect 220 147 240 167
rect 260 147 280 167
rect 300 147 320 167
rect 340 147 360 167
rect 380 147 400 167
rect 420 147 440 167
rect 460 147 480 167
rect 500 147 520 167
rect 540 147 560 167
rect 580 147 600 167
rect 620 147 640 167
rect 660 147 680 167
rect 700 147 720 167
rect 740 147 760 167
rect 780 147 800 167
rect 820 147 840 167
rect 860 147 880 167
rect 900 147 920 167
rect 940 147 960 167
rect 980 147 1000 167
rect 1020 147 1040 167
rect 1060 147 1080 167
rect 1100 147 1120 167
rect 1140 147 1160 167
rect 1180 147 1200 167
rect 1220 147 1240 167
rect 1260 147 1280 167
rect 1300 147 1320 167
rect 1340 147 1360 167
rect 1380 147 1400 167
rect 1420 147 1440 167
rect 1460 147 1480 167
rect 1500 147 1520 167
rect 1540 147 1560 167
rect 1580 147 1600 167
rect 1620 147 1640 167
rect 1660 147 1680 167
rect 1700 147 1720 167
rect 1740 147 1760 167
rect 1780 147 1800 167
rect 1820 147 1840 167
rect 1860 147 1880 167
rect 1900 147 1920 167
rect 1940 147 1960 167
rect 1980 147 2000 167
rect 2020 147 2040 167
rect 2060 147 2080 167
rect 2100 147 2120 167
rect 2140 147 2160 167
rect 2180 147 2200 167
rect 2220 147 2240 167
rect 2260 147 2280 167
rect 2300 147 2320 167
rect 2340 147 2360 167
rect 2380 147 2400 167
rect 2420 147 2440 167
rect 2460 147 2480 167
rect 2500 147 2520 167
rect 2540 147 2560 167
rect 2580 147 2600 167
rect 2620 147 2640 167
rect 2660 147 2675 167
rect 175 132 2675 147
rect 175 85 2675 100
rect 175 65 200 85
rect 220 65 240 85
rect 260 65 280 85
rect 300 65 320 85
rect 340 65 360 85
rect 380 65 400 85
rect 420 65 440 85
rect 460 65 480 85
rect 500 65 520 85
rect 540 65 560 85
rect 580 65 600 85
rect 620 65 640 85
rect 660 65 680 85
rect 700 65 720 85
rect 740 65 760 85
rect 780 65 800 85
rect 820 65 840 85
rect 860 65 880 85
rect 900 65 920 85
rect 940 65 960 85
rect 980 65 1000 85
rect 1020 65 1040 85
rect 1060 65 1080 85
rect 1100 65 1120 85
rect 1140 65 1160 85
rect 1180 65 1200 85
rect 1220 65 1240 85
rect 1260 65 1280 85
rect 1300 65 1320 85
rect 1340 65 1360 85
rect 1380 65 1400 85
rect 1420 65 1440 85
rect 1460 65 1480 85
rect 1500 65 1520 85
rect 1540 65 1560 85
rect 1580 65 1600 85
rect 1620 65 1640 85
rect 1660 65 1680 85
rect 1700 65 1720 85
rect 1740 65 1760 85
rect 1780 65 1800 85
rect 1820 65 1840 85
rect 1860 65 1880 85
rect 1900 65 1920 85
rect 1940 65 1960 85
rect 1980 65 2000 85
rect 2020 65 2040 85
rect 2060 65 2080 85
rect 2100 65 2120 85
rect 2140 65 2160 85
rect 2180 65 2200 85
rect 2220 65 2240 85
rect 2260 65 2280 85
rect 2300 65 2320 85
rect 2340 65 2360 85
rect 2380 65 2400 85
rect 2420 65 2440 85
rect 2460 65 2480 85
rect 2500 65 2520 85
rect 2540 65 2560 85
rect 2580 65 2600 85
rect 2620 65 2640 85
rect 2660 65 2675 85
rect 175 55 2675 65
rect 105 -265 2605 -255
rect 105 -285 120 -265
rect 140 -285 160 -265
rect 180 -285 200 -265
rect 220 -285 240 -265
rect 260 -285 280 -265
rect 300 -285 320 -265
rect 340 -285 360 -265
rect 380 -285 400 -265
rect 420 -285 440 -265
rect 460 -285 480 -265
rect 500 -285 520 -265
rect 540 -285 560 -265
rect 580 -285 600 -265
rect 620 -285 640 -265
rect 660 -285 680 -265
rect 700 -285 720 -265
rect 740 -285 760 -265
rect 780 -285 800 -265
rect 820 -285 840 -265
rect 860 -285 880 -265
rect 900 -285 920 -265
rect 940 -285 960 -265
rect 980 -285 1000 -265
rect 1020 -285 1040 -265
rect 1060 -285 1080 -265
rect 1100 -285 1120 -265
rect 1140 -285 1160 -265
rect 1180 -285 1200 -265
rect 1220 -285 1240 -265
rect 1260 -285 1280 -265
rect 1300 -285 1320 -265
rect 1340 -285 1360 -265
rect 1380 -285 1400 -265
rect 1420 -285 1440 -265
rect 1460 -285 1480 -265
rect 1500 -285 1520 -265
rect 1540 -285 1560 -265
rect 1580 -285 1600 -265
rect 1620 -285 1640 -265
rect 1660 -285 1680 -265
rect 1700 -285 1720 -265
rect 1740 -285 1760 -265
rect 1780 -285 1800 -265
rect 1820 -285 1840 -265
rect 1860 -285 1880 -265
rect 1900 -285 1920 -265
rect 1940 -285 1960 -265
rect 1980 -285 2000 -265
rect 2020 -285 2040 -265
rect 2060 -285 2080 -265
rect 2100 -285 2120 -265
rect 2140 -285 2160 -265
rect 2180 -285 2200 -265
rect 2220 -285 2240 -265
rect 2260 -285 2280 -265
rect 2300 -285 2320 -265
rect 2340 -285 2360 -265
rect 2380 -285 2400 -265
rect 2420 -285 2440 -265
rect 2460 -285 2480 -265
rect 2500 -285 2520 -265
rect 2540 -285 2560 -265
rect 2590 -285 2605 -265
rect 105 -300 2605 -285
rect 105 -360 2605 -345
rect 105 -380 120 -360
rect 140 -380 160 -360
rect 180 -380 200 -360
rect 220 -380 240 -360
rect 260 -380 280 -360
rect 300 -380 320 -360
rect 340 -380 360 -360
rect 380 -380 400 -360
rect 420 -380 440 -360
rect 460 -380 480 -360
rect 500 -380 520 -360
rect 540 -380 560 -360
rect 580 -380 600 -360
rect 620 -380 640 -360
rect 660 -380 680 -360
rect 700 -380 720 -360
rect 740 -380 760 -360
rect 780 -380 800 -360
rect 820 -380 840 -360
rect 860 -380 880 -360
rect 900 -380 920 -360
rect 940 -380 960 -360
rect 980 -380 1000 -360
rect 1020 -380 1040 -360
rect 1060 -380 1080 -360
rect 1100 -380 1120 -360
rect 1140 -380 1160 -360
rect 1180 -380 1200 -360
rect 1220 -380 1240 -360
rect 1260 -380 1280 -360
rect 1300 -380 1320 -360
rect 1340 -380 1360 -360
rect 1380 -380 1400 -360
rect 1420 -380 1440 -360
rect 1460 -380 1480 -360
rect 1500 -380 1520 -360
rect 1540 -380 1560 -360
rect 1580 -380 1600 -360
rect 1620 -380 1640 -360
rect 1660 -380 1680 -360
rect 1700 -380 1720 -360
rect 1740 -380 1760 -360
rect 1780 -380 1800 -360
rect 1820 -380 1840 -360
rect 1860 -380 1880 -360
rect 1900 -380 1920 -360
rect 1940 -380 1960 -360
rect 1980 -380 2000 -360
rect 2020 -380 2040 -360
rect 2060 -380 2080 -360
rect 2100 -380 2120 -360
rect 2140 -380 2160 -360
rect 2180 -380 2200 -360
rect 2220 -380 2240 -360
rect 2260 -380 2280 -360
rect 2300 -380 2320 -360
rect 2340 -380 2360 -360
rect 2380 -380 2400 -360
rect 2420 -380 2440 -360
rect 2460 -380 2480 -360
rect 2500 -380 2520 -360
rect 2540 -380 2560 -360
rect 2590 -380 2605 -360
rect 105 -395 2605 -380
rect 105 -455 2605 -440
rect 105 -475 120 -455
rect 140 -475 160 -455
rect 180 -475 200 -455
rect 220 -475 240 -455
rect 260 -475 280 -455
rect 300 -475 320 -455
rect 340 -475 360 -455
rect 380 -475 400 -455
rect 420 -475 440 -455
rect 460 -475 480 -455
rect 500 -475 520 -455
rect 540 -475 560 -455
rect 580 -475 600 -455
rect 620 -475 640 -455
rect 660 -475 680 -455
rect 700 -475 720 -455
rect 740 -475 760 -455
rect 780 -475 800 -455
rect 820 -475 840 -455
rect 860 -475 880 -455
rect 900 -475 920 -455
rect 940 -475 960 -455
rect 980 -475 1000 -455
rect 1020 -475 1040 -455
rect 1060 -475 1080 -455
rect 1100 -475 1120 -455
rect 1140 -475 1160 -455
rect 1180 -475 1200 -455
rect 1220 -475 1240 -455
rect 1260 -475 1280 -455
rect 1300 -475 1320 -455
rect 1340 -475 1360 -455
rect 1380 -475 1400 -455
rect 1420 -475 1440 -455
rect 1460 -475 1480 -455
rect 1500 -475 1520 -455
rect 1540 -475 1560 -455
rect 1580 -475 1600 -455
rect 1620 -475 1640 -455
rect 1660 -475 1680 -455
rect 1700 -475 1720 -455
rect 1740 -475 1760 -455
rect 1780 -475 1800 -455
rect 1820 -475 1840 -455
rect 1860 -475 1880 -455
rect 1900 -475 1920 -455
rect 1940 -475 1960 -455
rect 1980 -475 2000 -455
rect 2020 -475 2040 -455
rect 2060 -475 2080 -455
rect 2100 -475 2120 -455
rect 2140 -475 2160 -455
rect 2180 -475 2200 -455
rect 2220 -475 2240 -455
rect 2260 -475 2280 -455
rect 2300 -475 2320 -455
rect 2340 -475 2360 -455
rect 2380 -475 2400 -455
rect 2420 -475 2440 -455
rect 2460 -475 2480 -455
rect 2500 -475 2520 -455
rect 2540 -475 2560 -455
rect 2590 -475 2605 -455
rect 105 -490 2605 -475
rect 105 -550 2605 -535
rect 105 -570 120 -550
rect 140 -570 160 -550
rect 180 -570 200 -550
rect 220 -570 240 -550
rect 260 -570 280 -550
rect 300 -570 320 -550
rect 340 -570 360 -550
rect 380 -570 400 -550
rect 420 -570 440 -550
rect 460 -570 480 -550
rect 500 -570 520 -550
rect 540 -570 560 -550
rect 580 -570 600 -550
rect 620 -570 640 -550
rect 660 -570 680 -550
rect 700 -570 720 -550
rect 740 -570 760 -550
rect 780 -570 800 -550
rect 820 -570 840 -550
rect 860 -570 880 -550
rect 900 -570 920 -550
rect 940 -570 960 -550
rect 980 -570 1000 -550
rect 1020 -570 1040 -550
rect 1060 -570 1080 -550
rect 1100 -570 1120 -550
rect 1140 -570 1160 -550
rect 1180 -570 1200 -550
rect 1220 -570 1240 -550
rect 1260 -570 1280 -550
rect 1300 -570 1320 -550
rect 1340 -570 1360 -550
rect 1380 -570 1400 -550
rect 1420 -570 1440 -550
rect 1460 -570 1480 -550
rect 1500 -570 1520 -550
rect 1540 -570 1560 -550
rect 1580 -570 1600 -550
rect 1620 -570 1640 -550
rect 1660 -570 1680 -550
rect 1700 -570 1720 -550
rect 1740 -570 1760 -550
rect 1780 -570 1800 -550
rect 1820 -570 1840 -550
rect 1860 -570 1880 -550
rect 1900 -570 1920 -550
rect 1940 -570 1960 -550
rect 1980 -570 2000 -550
rect 2020 -570 2040 -550
rect 2060 -570 2080 -550
rect 2100 -570 2120 -550
rect 2140 -570 2160 -550
rect 2180 -570 2200 -550
rect 2220 -570 2240 -550
rect 2260 -570 2280 -550
rect 2300 -570 2320 -550
rect 2340 -570 2360 -550
rect 2380 -570 2400 -550
rect 2420 -570 2440 -550
rect 2460 -570 2480 -550
rect 2500 -570 2520 -550
rect 2540 -570 2560 -550
rect 2590 -570 2605 -550
rect 105 -585 2605 -570
rect 105 -645 2605 -630
rect 105 -665 120 -645
rect 140 -665 160 -645
rect 180 -665 200 -645
rect 220 -665 240 -645
rect 260 -665 280 -645
rect 300 -665 320 -645
rect 340 -665 360 -645
rect 380 -665 400 -645
rect 420 -665 440 -645
rect 460 -665 480 -645
rect 500 -665 520 -645
rect 540 -665 560 -645
rect 580 -665 600 -645
rect 620 -665 640 -645
rect 660 -665 680 -645
rect 700 -665 720 -645
rect 740 -665 760 -645
rect 780 -665 800 -645
rect 820 -665 840 -645
rect 860 -665 880 -645
rect 900 -665 920 -645
rect 940 -665 960 -645
rect 980 -665 1000 -645
rect 1020 -665 1040 -645
rect 1060 -665 1080 -645
rect 1100 -665 1120 -645
rect 1140 -665 1160 -645
rect 1180 -665 1200 -645
rect 1220 -665 1240 -645
rect 1260 -665 1280 -645
rect 1300 -665 1320 -645
rect 1340 -665 1360 -645
rect 1380 -665 1400 -645
rect 1420 -665 1440 -645
rect 1460 -665 1480 -645
rect 1500 -665 1520 -645
rect 1540 -665 1560 -645
rect 1580 -665 1600 -645
rect 1620 -665 1640 -645
rect 1660 -665 1680 -645
rect 1700 -665 1720 -645
rect 1740 -665 1760 -645
rect 1780 -665 1800 -645
rect 1820 -665 1840 -645
rect 1860 -665 1880 -645
rect 1900 -665 1920 -645
rect 1940 -665 1960 -645
rect 1980 -665 2000 -645
rect 2020 -665 2040 -645
rect 2060 -665 2080 -645
rect 2100 -665 2120 -645
rect 2140 -665 2160 -645
rect 2180 -665 2200 -645
rect 2220 -665 2240 -645
rect 2260 -665 2280 -645
rect 2300 -665 2320 -645
rect 2340 -665 2360 -645
rect 2380 -665 2400 -645
rect 2420 -665 2440 -645
rect 2460 -665 2480 -645
rect 2500 -665 2520 -645
rect 2540 -665 2560 -645
rect 2590 -665 2605 -645
rect 105 -680 2605 -665
rect 105 -740 2605 -725
rect 105 -760 120 -740
rect 140 -760 160 -740
rect 180 -760 200 -740
rect 220 -760 240 -740
rect 260 -760 280 -740
rect 300 -760 320 -740
rect 340 -760 360 -740
rect 380 -760 400 -740
rect 420 -760 440 -740
rect 460 -760 480 -740
rect 500 -760 520 -740
rect 540 -760 560 -740
rect 580 -760 600 -740
rect 620 -760 640 -740
rect 660 -760 680 -740
rect 700 -760 720 -740
rect 740 -760 760 -740
rect 780 -760 800 -740
rect 820 -760 840 -740
rect 860 -760 880 -740
rect 900 -760 920 -740
rect 940 -760 960 -740
rect 980 -760 1000 -740
rect 1020 -760 1040 -740
rect 1060 -760 1080 -740
rect 1100 -760 1120 -740
rect 1140 -760 1160 -740
rect 1180 -760 1200 -740
rect 1220 -760 1240 -740
rect 1260 -760 1280 -740
rect 1300 -760 1320 -740
rect 1340 -760 1360 -740
rect 1380 -760 1400 -740
rect 1420 -760 1440 -740
rect 1460 -760 1480 -740
rect 1500 -760 1520 -740
rect 1540 -760 1560 -740
rect 1580 -760 1600 -740
rect 1620 -760 1640 -740
rect 1660 -760 1680 -740
rect 1700 -760 1720 -740
rect 1740 -760 1760 -740
rect 1780 -760 1800 -740
rect 1820 -760 1840 -740
rect 1860 -760 1880 -740
rect 1900 -760 1920 -740
rect 1940 -760 1960 -740
rect 1980 -760 2000 -740
rect 2020 -760 2040 -740
rect 2060 -760 2080 -740
rect 2100 -760 2120 -740
rect 2140 -760 2160 -740
rect 2180 -760 2200 -740
rect 2220 -760 2240 -740
rect 2260 -760 2280 -740
rect 2300 -760 2320 -740
rect 2340 -760 2360 -740
rect 2380 -760 2400 -740
rect 2420 -760 2440 -740
rect 2460 -760 2480 -740
rect 2500 -760 2520 -740
rect 2540 -760 2560 -740
rect 2590 -760 2605 -740
rect 105 -775 2605 -760
rect 105 -835 2605 -820
rect 105 -855 120 -835
rect 140 -855 160 -835
rect 180 -855 200 -835
rect 220 -855 240 -835
rect 260 -855 280 -835
rect 300 -855 320 -835
rect 340 -855 360 -835
rect 380 -855 400 -835
rect 420 -855 440 -835
rect 460 -855 480 -835
rect 500 -855 520 -835
rect 540 -855 560 -835
rect 580 -855 600 -835
rect 620 -855 640 -835
rect 660 -855 680 -835
rect 700 -855 720 -835
rect 740 -855 760 -835
rect 780 -855 800 -835
rect 820 -855 840 -835
rect 860 -855 880 -835
rect 900 -855 920 -835
rect 940 -855 960 -835
rect 980 -855 1000 -835
rect 1020 -855 1040 -835
rect 1060 -855 1080 -835
rect 1100 -855 1120 -835
rect 1140 -855 1160 -835
rect 1180 -855 1200 -835
rect 1220 -855 1240 -835
rect 1260 -855 1280 -835
rect 1300 -855 1320 -835
rect 1340 -855 1360 -835
rect 1380 -855 1400 -835
rect 1420 -855 1440 -835
rect 1460 -855 1480 -835
rect 1500 -855 1520 -835
rect 1540 -855 1560 -835
rect 1580 -855 1600 -835
rect 1620 -855 1640 -835
rect 1660 -855 1680 -835
rect 1700 -855 1720 -835
rect 1740 -855 1760 -835
rect 1780 -855 1800 -835
rect 1820 -855 1840 -835
rect 1860 -855 1880 -835
rect 1900 -855 1920 -835
rect 1940 -855 1960 -835
rect 1980 -855 2000 -835
rect 2020 -855 2040 -835
rect 2060 -855 2080 -835
rect 2100 -855 2120 -835
rect 2140 -855 2160 -835
rect 2180 -855 2200 -835
rect 2220 -855 2240 -835
rect 2260 -855 2280 -835
rect 2300 -855 2320 -835
rect 2340 -855 2360 -835
rect 2380 -855 2400 -835
rect 2420 -855 2440 -835
rect 2460 -855 2480 -835
rect 2500 -855 2520 -835
rect 2540 -855 2560 -835
rect 2590 -855 2605 -835
rect 105 -870 2605 -855
rect 105 -930 2605 -915
rect 105 -950 120 -930
rect 140 -950 160 -930
rect 180 -950 200 -930
rect 220 -950 240 -930
rect 260 -950 280 -930
rect 300 -950 320 -930
rect 340 -950 360 -930
rect 380 -950 400 -930
rect 420 -950 440 -930
rect 460 -950 480 -930
rect 500 -950 520 -930
rect 540 -950 560 -930
rect 580 -950 600 -930
rect 620 -950 640 -930
rect 660 -950 680 -930
rect 700 -950 720 -930
rect 740 -950 760 -930
rect 780 -950 800 -930
rect 820 -950 840 -930
rect 860 -950 880 -930
rect 900 -950 920 -930
rect 940 -950 960 -930
rect 980 -950 1000 -930
rect 1020 -950 1040 -930
rect 1060 -950 1080 -930
rect 1100 -950 1120 -930
rect 1140 -950 1160 -930
rect 1180 -950 1200 -930
rect 1220 -950 1240 -930
rect 1260 -950 1280 -930
rect 1300 -950 1320 -930
rect 1340 -950 1360 -930
rect 1380 -950 1400 -930
rect 1420 -950 1440 -930
rect 1460 -950 1480 -930
rect 1500 -950 1520 -930
rect 1540 -950 1560 -930
rect 1580 -950 1600 -930
rect 1620 -950 1640 -930
rect 1660 -950 1680 -930
rect 1700 -950 1720 -930
rect 1740 -950 1760 -930
rect 1780 -950 1800 -930
rect 1820 -950 1840 -930
rect 1860 -950 1880 -930
rect 1900 -950 1920 -930
rect 1940 -950 1960 -930
rect 1980 -950 2000 -930
rect 2020 -950 2040 -930
rect 2060 -950 2080 -930
rect 2100 -950 2120 -930
rect 2140 -950 2160 -930
rect 2180 -950 2200 -930
rect 2220 -950 2240 -930
rect 2260 -950 2280 -930
rect 2300 -950 2320 -930
rect 2340 -950 2360 -930
rect 2380 -950 2400 -930
rect 2420 -950 2440 -930
rect 2460 -950 2480 -930
rect 2500 -950 2520 -930
rect 2540 -950 2560 -930
rect 2590 -950 2605 -930
rect 105 -965 2605 -950
rect 105 -1025 2605 -1010
rect 105 -1045 120 -1025
rect 140 -1045 160 -1025
rect 180 -1045 200 -1025
rect 220 -1045 240 -1025
rect 260 -1045 280 -1025
rect 300 -1045 320 -1025
rect 340 -1045 360 -1025
rect 380 -1045 400 -1025
rect 420 -1045 440 -1025
rect 460 -1045 480 -1025
rect 500 -1045 520 -1025
rect 540 -1045 560 -1025
rect 580 -1045 600 -1025
rect 620 -1045 640 -1025
rect 660 -1045 680 -1025
rect 700 -1045 720 -1025
rect 740 -1045 760 -1025
rect 780 -1045 800 -1025
rect 820 -1045 840 -1025
rect 860 -1045 880 -1025
rect 900 -1045 920 -1025
rect 940 -1045 960 -1025
rect 980 -1045 1000 -1025
rect 1020 -1045 1040 -1025
rect 1060 -1045 1080 -1025
rect 1100 -1045 1120 -1025
rect 1140 -1045 1160 -1025
rect 1180 -1045 1200 -1025
rect 1220 -1045 1240 -1025
rect 1260 -1045 1280 -1025
rect 1300 -1045 1320 -1025
rect 1340 -1045 1360 -1025
rect 1380 -1045 1400 -1025
rect 1420 -1045 1440 -1025
rect 1460 -1045 1480 -1025
rect 1500 -1045 1520 -1025
rect 1540 -1045 1560 -1025
rect 1580 -1045 1600 -1025
rect 1620 -1045 1640 -1025
rect 1660 -1045 1680 -1025
rect 1700 -1045 1720 -1025
rect 1740 -1045 1760 -1025
rect 1780 -1045 1800 -1025
rect 1820 -1045 1840 -1025
rect 1860 -1045 1880 -1025
rect 1900 -1045 1920 -1025
rect 1940 -1045 1960 -1025
rect 1980 -1045 2000 -1025
rect 2020 -1045 2040 -1025
rect 2060 -1045 2080 -1025
rect 2100 -1045 2120 -1025
rect 2140 -1045 2160 -1025
rect 2180 -1045 2200 -1025
rect 2220 -1045 2240 -1025
rect 2260 -1045 2280 -1025
rect 2300 -1045 2320 -1025
rect 2340 -1045 2360 -1025
rect 2380 -1045 2400 -1025
rect 2420 -1045 2440 -1025
rect 2460 -1045 2480 -1025
rect 2500 -1045 2520 -1025
rect 2540 -1045 2560 -1025
rect 2590 -1045 2605 -1025
rect 105 -1060 2605 -1045
rect 105 -1120 2605 -1105
rect 105 -1140 120 -1120
rect 140 -1140 160 -1120
rect 180 -1140 200 -1120
rect 220 -1140 240 -1120
rect 260 -1140 280 -1120
rect 300 -1140 320 -1120
rect 340 -1140 360 -1120
rect 380 -1140 400 -1120
rect 420 -1140 440 -1120
rect 460 -1140 480 -1120
rect 500 -1140 520 -1120
rect 540 -1140 560 -1120
rect 580 -1140 600 -1120
rect 620 -1140 640 -1120
rect 660 -1140 680 -1120
rect 700 -1140 720 -1120
rect 740 -1140 760 -1120
rect 780 -1140 800 -1120
rect 820 -1140 840 -1120
rect 860 -1140 880 -1120
rect 900 -1140 920 -1120
rect 940 -1140 960 -1120
rect 980 -1140 1000 -1120
rect 1020 -1140 1040 -1120
rect 1060 -1140 1080 -1120
rect 1100 -1140 1120 -1120
rect 1140 -1140 1160 -1120
rect 1180 -1140 1200 -1120
rect 1220 -1140 1240 -1120
rect 1260 -1140 1280 -1120
rect 1300 -1140 1320 -1120
rect 1340 -1140 1360 -1120
rect 1380 -1140 1400 -1120
rect 1420 -1140 1440 -1120
rect 1460 -1140 1480 -1120
rect 1500 -1140 1520 -1120
rect 1540 -1140 1560 -1120
rect 1580 -1140 1600 -1120
rect 1620 -1140 1640 -1120
rect 1660 -1140 1680 -1120
rect 1700 -1140 1720 -1120
rect 1740 -1140 1760 -1120
rect 1780 -1140 1800 -1120
rect 1820 -1140 1840 -1120
rect 1860 -1140 1880 -1120
rect 1900 -1140 1920 -1120
rect 1940 -1140 1960 -1120
rect 1980 -1140 2000 -1120
rect 2020 -1140 2040 -1120
rect 2060 -1140 2080 -1120
rect 2100 -1140 2120 -1120
rect 2140 -1140 2160 -1120
rect 2180 -1140 2200 -1120
rect 2220 -1140 2240 -1120
rect 2260 -1140 2280 -1120
rect 2300 -1140 2320 -1120
rect 2340 -1140 2360 -1120
rect 2380 -1140 2400 -1120
rect 2420 -1140 2440 -1120
rect 2460 -1140 2480 -1120
rect 2500 -1140 2520 -1120
rect 2540 -1140 2560 -1120
rect 2590 -1140 2605 -1120
rect 105 -1155 2605 -1140
rect 105 -1215 2605 -1200
rect 105 -1235 120 -1215
rect 140 -1235 160 -1215
rect 180 -1235 200 -1215
rect 220 -1235 240 -1215
rect 260 -1235 280 -1215
rect 300 -1235 320 -1215
rect 340 -1235 360 -1215
rect 380 -1235 400 -1215
rect 420 -1235 440 -1215
rect 460 -1235 480 -1215
rect 500 -1235 520 -1215
rect 540 -1235 560 -1215
rect 580 -1235 600 -1215
rect 620 -1235 640 -1215
rect 660 -1235 680 -1215
rect 700 -1235 720 -1215
rect 740 -1235 760 -1215
rect 780 -1235 800 -1215
rect 820 -1235 840 -1215
rect 860 -1235 880 -1215
rect 900 -1235 920 -1215
rect 940 -1235 960 -1215
rect 980 -1235 1000 -1215
rect 1020 -1235 1040 -1215
rect 1060 -1235 1080 -1215
rect 1100 -1235 1120 -1215
rect 1140 -1235 1160 -1215
rect 1180 -1235 1200 -1215
rect 1220 -1235 1240 -1215
rect 1260 -1235 1280 -1215
rect 1300 -1235 1320 -1215
rect 1340 -1235 1360 -1215
rect 1380 -1235 1400 -1215
rect 1420 -1235 1440 -1215
rect 1460 -1235 1480 -1215
rect 1500 -1235 1520 -1215
rect 1540 -1235 1560 -1215
rect 1580 -1235 1600 -1215
rect 1620 -1235 1640 -1215
rect 1660 -1235 1680 -1215
rect 1700 -1235 1720 -1215
rect 1740 -1235 1760 -1215
rect 1780 -1235 1800 -1215
rect 1820 -1235 1840 -1215
rect 1860 -1235 1880 -1215
rect 1900 -1235 1920 -1215
rect 1940 -1235 1960 -1215
rect 1980 -1235 2000 -1215
rect 2020 -1235 2040 -1215
rect 2060 -1235 2080 -1215
rect 2100 -1235 2120 -1215
rect 2140 -1235 2160 -1215
rect 2180 -1235 2200 -1215
rect 2220 -1235 2240 -1215
rect 2260 -1235 2280 -1215
rect 2300 -1235 2320 -1215
rect 2340 -1235 2360 -1215
rect 2380 -1235 2400 -1215
rect 2420 -1235 2440 -1215
rect 2460 -1235 2480 -1215
rect 2500 -1235 2520 -1215
rect 2540 -1235 2560 -1215
rect 2590 -1235 2605 -1215
rect 105 -1250 2605 -1235
rect 105 -1310 2605 -1295
rect 105 -1330 120 -1310
rect 140 -1330 160 -1310
rect 180 -1330 200 -1310
rect 220 -1330 240 -1310
rect 260 -1330 280 -1310
rect 300 -1330 320 -1310
rect 340 -1330 360 -1310
rect 380 -1330 400 -1310
rect 420 -1330 440 -1310
rect 460 -1330 480 -1310
rect 500 -1330 520 -1310
rect 540 -1330 560 -1310
rect 580 -1330 600 -1310
rect 620 -1330 640 -1310
rect 660 -1330 680 -1310
rect 700 -1330 720 -1310
rect 740 -1330 760 -1310
rect 780 -1330 800 -1310
rect 820 -1330 840 -1310
rect 860 -1330 880 -1310
rect 900 -1330 920 -1310
rect 940 -1330 960 -1310
rect 980 -1330 1000 -1310
rect 1020 -1330 1040 -1310
rect 1060 -1330 1080 -1310
rect 1100 -1330 1120 -1310
rect 1140 -1330 1160 -1310
rect 1180 -1330 1200 -1310
rect 1220 -1330 1240 -1310
rect 1260 -1330 1280 -1310
rect 1300 -1330 1320 -1310
rect 1340 -1330 1360 -1310
rect 1380 -1330 1400 -1310
rect 1420 -1330 1440 -1310
rect 1460 -1330 1480 -1310
rect 1500 -1330 1520 -1310
rect 1540 -1330 1560 -1310
rect 1580 -1330 1600 -1310
rect 1620 -1330 1640 -1310
rect 1660 -1330 1680 -1310
rect 1700 -1330 1720 -1310
rect 1740 -1330 1760 -1310
rect 1780 -1330 1800 -1310
rect 1820 -1330 1840 -1310
rect 1860 -1330 1880 -1310
rect 1900 -1330 1920 -1310
rect 1940 -1330 1960 -1310
rect 1980 -1330 2000 -1310
rect 2020 -1330 2040 -1310
rect 2060 -1330 2080 -1310
rect 2100 -1330 2120 -1310
rect 2140 -1330 2160 -1310
rect 2180 -1330 2200 -1310
rect 2220 -1330 2240 -1310
rect 2260 -1330 2280 -1310
rect 2300 -1330 2320 -1310
rect 2340 -1330 2360 -1310
rect 2380 -1330 2400 -1310
rect 2420 -1330 2440 -1310
rect 2460 -1330 2480 -1310
rect 2500 -1330 2520 -1310
rect 2540 -1330 2560 -1310
rect 2590 -1330 2605 -1310
rect 105 -1345 2605 -1330
rect 105 -1405 2605 -1390
rect 105 -1425 120 -1405
rect 140 -1425 160 -1405
rect 180 -1425 200 -1405
rect 220 -1425 240 -1405
rect 260 -1425 280 -1405
rect 300 -1425 320 -1405
rect 340 -1425 360 -1405
rect 380 -1425 400 -1405
rect 420 -1425 440 -1405
rect 460 -1425 480 -1405
rect 500 -1425 520 -1405
rect 540 -1425 560 -1405
rect 580 -1425 600 -1405
rect 620 -1425 640 -1405
rect 660 -1425 680 -1405
rect 700 -1425 720 -1405
rect 740 -1425 760 -1405
rect 780 -1425 800 -1405
rect 820 -1425 840 -1405
rect 860 -1425 880 -1405
rect 900 -1425 920 -1405
rect 940 -1425 960 -1405
rect 980 -1425 1000 -1405
rect 1020 -1425 1040 -1405
rect 1060 -1425 1080 -1405
rect 1100 -1425 1120 -1405
rect 1140 -1425 1160 -1405
rect 1180 -1425 1200 -1405
rect 1220 -1425 1240 -1405
rect 1260 -1425 1280 -1405
rect 1300 -1425 1320 -1405
rect 1340 -1425 1360 -1405
rect 1380 -1425 1400 -1405
rect 1420 -1425 1440 -1405
rect 1460 -1425 1480 -1405
rect 1500 -1425 1520 -1405
rect 1540 -1425 1560 -1405
rect 1580 -1425 1600 -1405
rect 1620 -1425 1640 -1405
rect 1660 -1425 1680 -1405
rect 1700 -1425 1720 -1405
rect 1740 -1425 1760 -1405
rect 1780 -1425 1800 -1405
rect 1820 -1425 1840 -1405
rect 1860 -1425 1880 -1405
rect 1900 -1425 1920 -1405
rect 1940 -1425 1960 -1405
rect 1980 -1425 2000 -1405
rect 2020 -1425 2040 -1405
rect 2060 -1425 2080 -1405
rect 2100 -1425 2120 -1405
rect 2140 -1425 2160 -1405
rect 2180 -1425 2200 -1405
rect 2220 -1425 2240 -1405
rect 2260 -1425 2280 -1405
rect 2300 -1425 2320 -1405
rect 2340 -1425 2360 -1405
rect 2380 -1425 2400 -1405
rect 2420 -1425 2440 -1405
rect 2460 -1425 2480 -1405
rect 2500 -1425 2520 -1405
rect 2540 -1425 2560 -1405
rect 2590 -1425 2605 -1405
rect 105 -1440 2605 -1425
rect 105 -1500 2605 -1485
rect 105 -1520 120 -1500
rect 140 -1520 160 -1500
rect 180 -1520 200 -1500
rect 220 -1520 240 -1500
rect 260 -1520 280 -1500
rect 300 -1520 320 -1500
rect 340 -1520 360 -1500
rect 380 -1520 400 -1500
rect 420 -1520 440 -1500
rect 460 -1520 480 -1500
rect 500 -1520 520 -1500
rect 540 -1520 560 -1500
rect 580 -1520 600 -1500
rect 620 -1520 640 -1500
rect 660 -1520 680 -1500
rect 700 -1520 720 -1500
rect 740 -1520 760 -1500
rect 780 -1520 800 -1500
rect 820 -1520 840 -1500
rect 860 -1520 880 -1500
rect 900 -1520 920 -1500
rect 940 -1520 960 -1500
rect 980 -1520 1000 -1500
rect 1020 -1520 1040 -1500
rect 1060 -1520 1080 -1500
rect 1100 -1520 1120 -1500
rect 1140 -1520 1160 -1500
rect 1180 -1520 1200 -1500
rect 1220 -1520 1240 -1500
rect 1260 -1520 1280 -1500
rect 1300 -1520 1320 -1500
rect 1340 -1520 1360 -1500
rect 1380 -1520 1400 -1500
rect 1420 -1520 1440 -1500
rect 1460 -1520 1480 -1500
rect 1500 -1520 1520 -1500
rect 1540 -1520 1560 -1500
rect 1580 -1520 1600 -1500
rect 1620 -1520 1640 -1500
rect 1660 -1520 1680 -1500
rect 1700 -1520 1720 -1500
rect 1740 -1520 1760 -1500
rect 1780 -1520 1800 -1500
rect 1820 -1520 1840 -1500
rect 1860 -1520 1880 -1500
rect 1900 -1520 1920 -1500
rect 1940 -1520 1960 -1500
rect 1980 -1520 2000 -1500
rect 2020 -1520 2040 -1500
rect 2060 -1520 2080 -1500
rect 2100 -1520 2120 -1500
rect 2140 -1520 2160 -1500
rect 2180 -1520 2200 -1500
rect 2220 -1520 2240 -1500
rect 2260 -1520 2280 -1500
rect 2300 -1520 2320 -1500
rect 2340 -1520 2360 -1500
rect 2380 -1520 2400 -1500
rect 2420 -1520 2440 -1500
rect 2460 -1520 2480 -1500
rect 2500 -1520 2520 -1500
rect 2540 -1520 2560 -1500
rect 2590 -1520 2605 -1500
rect 105 -1535 2605 -1520
rect 105 -1595 2605 -1580
rect 105 -1615 120 -1595
rect 140 -1615 160 -1595
rect 180 -1615 200 -1595
rect 220 -1615 240 -1595
rect 260 -1615 280 -1595
rect 300 -1615 320 -1595
rect 340 -1615 360 -1595
rect 380 -1615 400 -1595
rect 420 -1615 440 -1595
rect 460 -1615 480 -1595
rect 500 -1615 520 -1595
rect 540 -1615 560 -1595
rect 580 -1615 600 -1595
rect 620 -1615 640 -1595
rect 660 -1615 680 -1595
rect 700 -1615 720 -1595
rect 740 -1615 760 -1595
rect 780 -1615 800 -1595
rect 820 -1615 840 -1595
rect 860 -1615 880 -1595
rect 900 -1615 920 -1595
rect 940 -1615 960 -1595
rect 980 -1615 1000 -1595
rect 1020 -1615 1040 -1595
rect 1060 -1615 1080 -1595
rect 1100 -1615 1120 -1595
rect 1140 -1615 1160 -1595
rect 1180 -1615 1200 -1595
rect 1220 -1615 1240 -1595
rect 1260 -1615 1280 -1595
rect 1300 -1615 1320 -1595
rect 1340 -1615 1360 -1595
rect 1380 -1615 1400 -1595
rect 1420 -1615 1440 -1595
rect 1460 -1615 1480 -1595
rect 1500 -1615 1520 -1595
rect 1540 -1615 1560 -1595
rect 1580 -1615 1600 -1595
rect 1620 -1615 1640 -1595
rect 1660 -1615 1680 -1595
rect 1700 -1615 1720 -1595
rect 1740 -1615 1760 -1595
rect 1780 -1615 1800 -1595
rect 1820 -1615 1840 -1595
rect 1860 -1615 1880 -1595
rect 1900 -1615 1920 -1595
rect 1940 -1615 1960 -1595
rect 1980 -1615 2000 -1595
rect 2020 -1615 2040 -1595
rect 2060 -1615 2080 -1595
rect 2100 -1615 2120 -1595
rect 2140 -1615 2160 -1595
rect 2180 -1615 2200 -1595
rect 2220 -1615 2240 -1595
rect 2260 -1615 2280 -1595
rect 2300 -1615 2320 -1595
rect 2340 -1615 2360 -1595
rect 2380 -1615 2400 -1595
rect 2420 -1615 2440 -1595
rect 2460 -1615 2480 -1595
rect 2500 -1615 2520 -1595
rect 2540 -1615 2560 -1595
rect 2590 -1615 2605 -1595
rect 105 -1630 2605 -1615
rect 105 -1690 2605 -1675
rect 105 -1710 120 -1690
rect 140 -1710 160 -1690
rect 180 -1710 200 -1690
rect 220 -1710 240 -1690
rect 260 -1710 280 -1690
rect 300 -1710 320 -1690
rect 340 -1710 360 -1690
rect 380 -1710 400 -1690
rect 420 -1710 440 -1690
rect 460 -1710 480 -1690
rect 500 -1710 520 -1690
rect 540 -1710 560 -1690
rect 580 -1710 600 -1690
rect 620 -1710 640 -1690
rect 660 -1710 680 -1690
rect 700 -1710 720 -1690
rect 740 -1710 760 -1690
rect 780 -1710 800 -1690
rect 820 -1710 840 -1690
rect 860 -1710 880 -1690
rect 900 -1710 920 -1690
rect 940 -1710 960 -1690
rect 980 -1710 1000 -1690
rect 1020 -1710 1040 -1690
rect 1060 -1710 1080 -1690
rect 1100 -1710 1120 -1690
rect 1140 -1710 1160 -1690
rect 1180 -1710 1200 -1690
rect 1220 -1710 1240 -1690
rect 1260 -1710 1280 -1690
rect 1300 -1710 1320 -1690
rect 1340 -1710 1360 -1690
rect 1380 -1710 1400 -1690
rect 1420 -1710 1440 -1690
rect 1460 -1710 1480 -1690
rect 1500 -1710 1520 -1690
rect 1540 -1710 1560 -1690
rect 1580 -1710 1600 -1690
rect 1620 -1710 1640 -1690
rect 1660 -1710 1680 -1690
rect 1700 -1710 1720 -1690
rect 1740 -1710 1760 -1690
rect 1780 -1710 1800 -1690
rect 1820 -1710 1840 -1690
rect 1860 -1710 1880 -1690
rect 1900 -1710 1920 -1690
rect 1940 -1710 1960 -1690
rect 1980 -1710 2000 -1690
rect 2020 -1710 2040 -1690
rect 2060 -1710 2080 -1690
rect 2100 -1710 2120 -1690
rect 2140 -1710 2160 -1690
rect 2180 -1710 2200 -1690
rect 2220 -1710 2240 -1690
rect 2260 -1710 2280 -1690
rect 2300 -1710 2320 -1690
rect 2340 -1710 2360 -1690
rect 2380 -1710 2400 -1690
rect 2420 -1710 2440 -1690
rect 2460 -1710 2480 -1690
rect 2500 -1710 2520 -1690
rect 2540 -1710 2560 -1690
rect 2590 -1710 2605 -1690
rect 105 -1725 2605 -1710
rect 105 -1785 2605 -1770
rect 105 -1805 120 -1785
rect 140 -1805 160 -1785
rect 180 -1805 200 -1785
rect 220 -1805 240 -1785
rect 260 -1805 280 -1785
rect 300 -1805 320 -1785
rect 340 -1805 360 -1785
rect 380 -1805 400 -1785
rect 420 -1805 440 -1785
rect 460 -1805 480 -1785
rect 500 -1805 520 -1785
rect 540 -1805 560 -1785
rect 580 -1805 600 -1785
rect 620 -1805 640 -1785
rect 660 -1805 680 -1785
rect 700 -1805 720 -1785
rect 740 -1805 760 -1785
rect 780 -1805 800 -1785
rect 820 -1805 840 -1785
rect 860 -1805 880 -1785
rect 900 -1805 920 -1785
rect 940 -1805 960 -1785
rect 980 -1805 1000 -1785
rect 1020 -1805 1040 -1785
rect 1060 -1805 1080 -1785
rect 1100 -1805 1120 -1785
rect 1140 -1805 1160 -1785
rect 1180 -1805 1200 -1785
rect 1220 -1805 1240 -1785
rect 1260 -1805 1280 -1785
rect 1300 -1805 1320 -1785
rect 1340 -1805 1360 -1785
rect 1380 -1805 1400 -1785
rect 1420 -1805 1440 -1785
rect 1460 -1805 1480 -1785
rect 1500 -1805 1520 -1785
rect 1540 -1805 1560 -1785
rect 1580 -1805 1600 -1785
rect 1620 -1805 1640 -1785
rect 1660 -1805 1680 -1785
rect 1700 -1805 1720 -1785
rect 1740 -1805 1760 -1785
rect 1780 -1805 1800 -1785
rect 1820 -1805 1840 -1785
rect 1860 -1805 1880 -1785
rect 1900 -1805 1920 -1785
rect 1940 -1805 1960 -1785
rect 1980 -1805 2000 -1785
rect 2020 -1805 2040 -1785
rect 2060 -1805 2080 -1785
rect 2100 -1805 2120 -1785
rect 2140 -1805 2160 -1785
rect 2180 -1805 2200 -1785
rect 2220 -1805 2240 -1785
rect 2260 -1805 2280 -1785
rect 2300 -1805 2320 -1785
rect 2340 -1805 2360 -1785
rect 2380 -1805 2400 -1785
rect 2420 -1805 2440 -1785
rect 2460 -1805 2480 -1785
rect 2500 -1805 2520 -1785
rect 2540 -1805 2560 -1785
rect 2590 -1805 2605 -1785
rect 105 -1820 2605 -1805
rect 105 -1880 2605 -1865
rect 105 -1900 120 -1880
rect 140 -1900 160 -1880
rect 180 -1900 200 -1880
rect 220 -1900 240 -1880
rect 260 -1900 280 -1880
rect 300 -1900 320 -1880
rect 340 -1900 360 -1880
rect 380 -1900 400 -1880
rect 420 -1900 440 -1880
rect 460 -1900 480 -1880
rect 500 -1900 520 -1880
rect 540 -1900 560 -1880
rect 580 -1900 600 -1880
rect 620 -1900 640 -1880
rect 660 -1900 680 -1880
rect 700 -1900 720 -1880
rect 740 -1900 760 -1880
rect 780 -1900 800 -1880
rect 820 -1900 840 -1880
rect 860 -1900 880 -1880
rect 900 -1900 920 -1880
rect 940 -1900 960 -1880
rect 980 -1900 1000 -1880
rect 1020 -1900 1040 -1880
rect 1060 -1900 1080 -1880
rect 1100 -1900 1120 -1880
rect 1140 -1900 1160 -1880
rect 1180 -1900 1200 -1880
rect 1220 -1900 1240 -1880
rect 1260 -1900 1280 -1880
rect 1300 -1900 1320 -1880
rect 1340 -1900 1360 -1880
rect 1380 -1900 1400 -1880
rect 1420 -1900 1440 -1880
rect 1460 -1900 1480 -1880
rect 1500 -1900 1520 -1880
rect 1540 -1900 1560 -1880
rect 1580 -1900 1600 -1880
rect 1620 -1900 1640 -1880
rect 1660 -1900 1680 -1880
rect 1700 -1900 1720 -1880
rect 1740 -1900 1760 -1880
rect 1780 -1900 1800 -1880
rect 1820 -1900 1840 -1880
rect 1860 -1900 1880 -1880
rect 1900 -1900 1920 -1880
rect 1940 -1900 1960 -1880
rect 1980 -1900 2000 -1880
rect 2020 -1900 2040 -1880
rect 2060 -1900 2080 -1880
rect 2100 -1900 2120 -1880
rect 2140 -1900 2160 -1880
rect 2180 -1900 2200 -1880
rect 2220 -1900 2240 -1880
rect 2260 -1900 2280 -1880
rect 2300 -1900 2320 -1880
rect 2340 -1900 2360 -1880
rect 2380 -1900 2400 -1880
rect 2420 -1900 2440 -1880
rect 2460 -1900 2480 -1880
rect 2500 -1900 2520 -1880
rect 2540 -1900 2560 -1880
rect 2590 -1900 2605 -1880
rect 105 -1915 2605 -1900
rect 105 -1975 2605 -1960
rect 105 -1995 120 -1975
rect 140 -1995 160 -1975
rect 180 -1995 200 -1975
rect 220 -1995 240 -1975
rect 260 -1995 280 -1975
rect 300 -1995 320 -1975
rect 340 -1995 360 -1975
rect 380 -1995 400 -1975
rect 420 -1995 440 -1975
rect 460 -1995 480 -1975
rect 500 -1995 520 -1975
rect 540 -1995 560 -1975
rect 580 -1995 600 -1975
rect 620 -1995 640 -1975
rect 660 -1995 680 -1975
rect 700 -1995 720 -1975
rect 740 -1995 760 -1975
rect 780 -1995 800 -1975
rect 820 -1995 840 -1975
rect 860 -1995 880 -1975
rect 900 -1995 920 -1975
rect 940 -1995 960 -1975
rect 980 -1995 1000 -1975
rect 1020 -1995 1040 -1975
rect 1060 -1995 1080 -1975
rect 1100 -1995 1120 -1975
rect 1140 -1995 1160 -1975
rect 1180 -1995 1200 -1975
rect 1220 -1995 1240 -1975
rect 1260 -1995 1280 -1975
rect 1300 -1995 1320 -1975
rect 1340 -1995 1360 -1975
rect 1380 -1995 1400 -1975
rect 1420 -1995 1440 -1975
rect 1460 -1995 1480 -1975
rect 1500 -1995 1520 -1975
rect 1540 -1995 1560 -1975
rect 1580 -1995 1600 -1975
rect 1620 -1995 1640 -1975
rect 1660 -1995 1680 -1975
rect 1700 -1995 1720 -1975
rect 1740 -1995 1760 -1975
rect 1780 -1995 1800 -1975
rect 1820 -1995 1840 -1975
rect 1860 -1995 1880 -1975
rect 1900 -1995 1920 -1975
rect 1940 -1995 1960 -1975
rect 1980 -1995 2000 -1975
rect 2020 -1995 2040 -1975
rect 2060 -1995 2080 -1975
rect 2100 -1995 2120 -1975
rect 2140 -1995 2160 -1975
rect 2180 -1995 2200 -1975
rect 2220 -1995 2240 -1975
rect 2260 -1995 2280 -1975
rect 2300 -1995 2320 -1975
rect 2340 -1995 2360 -1975
rect 2380 -1995 2400 -1975
rect 2420 -1995 2440 -1975
rect 2460 -1995 2480 -1975
rect 2500 -1995 2520 -1975
rect 2540 -1995 2560 -1975
rect 2590 -1995 2605 -1975
rect 105 -2010 2605 -1995
rect 105 -2070 2605 -2055
rect 105 -2090 120 -2070
rect 140 -2090 160 -2070
rect 180 -2090 200 -2070
rect 220 -2090 240 -2070
rect 260 -2090 280 -2070
rect 300 -2090 320 -2070
rect 340 -2090 360 -2070
rect 380 -2090 400 -2070
rect 420 -2090 440 -2070
rect 460 -2090 480 -2070
rect 500 -2090 520 -2070
rect 540 -2090 560 -2070
rect 580 -2090 600 -2070
rect 620 -2090 640 -2070
rect 660 -2090 680 -2070
rect 700 -2090 720 -2070
rect 740 -2090 760 -2070
rect 780 -2090 800 -2070
rect 820 -2090 840 -2070
rect 860 -2090 880 -2070
rect 900 -2090 920 -2070
rect 940 -2090 960 -2070
rect 980 -2090 1000 -2070
rect 1020 -2090 1040 -2070
rect 1060 -2090 1080 -2070
rect 1100 -2090 1120 -2070
rect 1140 -2090 1160 -2070
rect 1180 -2090 1200 -2070
rect 1220 -2090 1240 -2070
rect 1260 -2090 1280 -2070
rect 1300 -2090 1320 -2070
rect 1340 -2090 1360 -2070
rect 1380 -2090 1400 -2070
rect 1420 -2090 1440 -2070
rect 1460 -2090 1480 -2070
rect 1500 -2090 1520 -2070
rect 1540 -2090 1560 -2070
rect 1580 -2090 1600 -2070
rect 1620 -2090 1640 -2070
rect 1660 -2090 1680 -2070
rect 1700 -2090 1720 -2070
rect 1740 -2090 1760 -2070
rect 1780 -2090 1800 -2070
rect 1820 -2090 1840 -2070
rect 1860 -2090 1880 -2070
rect 1900 -2090 1920 -2070
rect 1940 -2090 1960 -2070
rect 1980 -2090 2000 -2070
rect 2020 -2090 2040 -2070
rect 2060 -2090 2080 -2070
rect 2100 -2090 2120 -2070
rect 2140 -2090 2160 -2070
rect 2180 -2090 2200 -2070
rect 2220 -2090 2240 -2070
rect 2260 -2090 2280 -2070
rect 2300 -2090 2320 -2070
rect 2340 -2090 2360 -2070
rect 2380 -2090 2400 -2070
rect 2420 -2090 2440 -2070
rect 2460 -2090 2480 -2070
rect 2500 -2090 2520 -2070
rect 2540 -2090 2560 -2070
rect 2590 -2090 2605 -2070
rect 105 -2105 2605 -2090
rect 105 -2165 2605 -2150
rect 105 -2185 120 -2165
rect 140 -2185 160 -2165
rect 180 -2185 200 -2165
rect 220 -2185 240 -2165
rect 260 -2185 280 -2165
rect 300 -2185 320 -2165
rect 340 -2185 360 -2165
rect 380 -2185 400 -2165
rect 420 -2185 440 -2165
rect 460 -2185 480 -2165
rect 500 -2185 520 -2165
rect 540 -2185 560 -2165
rect 580 -2185 600 -2165
rect 620 -2185 640 -2165
rect 660 -2185 680 -2165
rect 700 -2185 720 -2165
rect 740 -2185 760 -2165
rect 780 -2185 800 -2165
rect 820 -2185 840 -2165
rect 860 -2185 880 -2165
rect 900 -2185 920 -2165
rect 940 -2185 960 -2165
rect 980 -2185 1000 -2165
rect 1020 -2185 1040 -2165
rect 1060 -2185 1080 -2165
rect 1100 -2185 1120 -2165
rect 1140 -2185 1160 -2165
rect 1180 -2185 1200 -2165
rect 1220 -2185 1240 -2165
rect 1260 -2185 1280 -2165
rect 1300 -2185 1320 -2165
rect 1340 -2185 1360 -2165
rect 1380 -2185 1400 -2165
rect 1420 -2185 1440 -2165
rect 1460 -2185 1480 -2165
rect 1500 -2185 1520 -2165
rect 1540 -2185 1560 -2165
rect 1580 -2185 1600 -2165
rect 1620 -2185 1640 -2165
rect 1660 -2185 1680 -2165
rect 1700 -2185 1720 -2165
rect 1740 -2185 1760 -2165
rect 1780 -2185 1800 -2165
rect 1820 -2185 1840 -2165
rect 1860 -2185 1880 -2165
rect 1900 -2185 1920 -2165
rect 1940 -2185 1960 -2165
rect 1980 -2185 2000 -2165
rect 2020 -2185 2040 -2165
rect 2060 -2185 2080 -2165
rect 2100 -2185 2120 -2165
rect 2140 -2185 2160 -2165
rect 2180 -2185 2200 -2165
rect 2220 -2185 2240 -2165
rect 2260 -2185 2280 -2165
rect 2300 -2185 2320 -2165
rect 2340 -2185 2360 -2165
rect 2380 -2185 2400 -2165
rect 2420 -2185 2440 -2165
rect 2460 -2185 2480 -2165
rect 2500 -2185 2520 -2165
rect 2540 -2185 2560 -2165
rect 2590 -2185 2605 -2165
rect 105 -2200 2605 -2185
rect 105 -2260 2605 -2245
rect 105 -2280 120 -2260
rect 140 -2280 160 -2260
rect 180 -2280 200 -2260
rect 220 -2280 240 -2260
rect 260 -2280 280 -2260
rect 300 -2280 320 -2260
rect 340 -2280 360 -2260
rect 380 -2280 400 -2260
rect 420 -2280 440 -2260
rect 460 -2280 480 -2260
rect 500 -2280 520 -2260
rect 540 -2280 560 -2260
rect 580 -2280 600 -2260
rect 620 -2280 640 -2260
rect 660 -2280 680 -2260
rect 700 -2280 720 -2260
rect 740 -2280 760 -2260
rect 780 -2280 800 -2260
rect 820 -2280 840 -2260
rect 860 -2280 880 -2260
rect 900 -2280 920 -2260
rect 940 -2280 960 -2260
rect 980 -2280 1000 -2260
rect 1020 -2280 1040 -2260
rect 1060 -2280 1080 -2260
rect 1100 -2280 1120 -2260
rect 1140 -2280 1160 -2260
rect 1180 -2280 1200 -2260
rect 1220 -2280 1240 -2260
rect 1260 -2280 1280 -2260
rect 1300 -2280 1320 -2260
rect 1340 -2280 1360 -2260
rect 1380 -2280 1400 -2260
rect 1420 -2280 1440 -2260
rect 1460 -2280 1480 -2260
rect 1500 -2280 1520 -2260
rect 1540 -2280 1560 -2260
rect 1580 -2280 1600 -2260
rect 1620 -2280 1640 -2260
rect 1660 -2280 1680 -2260
rect 1700 -2280 1720 -2260
rect 1740 -2280 1760 -2260
rect 1780 -2280 1800 -2260
rect 1820 -2280 1840 -2260
rect 1860 -2280 1880 -2260
rect 1900 -2280 1920 -2260
rect 1940 -2280 1960 -2260
rect 1980 -2280 2000 -2260
rect 2020 -2280 2040 -2260
rect 2060 -2280 2080 -2260
rect 2100 -2280 2120 -2260
rect 2140 -2280 2160 -2260
rect 2180 -2280 2200 -2260
rect 2220 -2280 2240 -2260
rect 2260 -2280 2280 -2260
rect 2300 -2280 2320 -2260
rect 2340 -2280 2360 -2260
rect 2380 -2280 2400 -2260
rect 2420 -2280 2440 -2260
rect 2460 -2280 2480 -2260
rect 2500 -2280 2520 -2260
rect 2540 -2280 2560 -2260
rect 2590 -2280 2605 -2260
rect 105 -2295 2605 -2280
rect 105 -2355 2605 -2340
rect 105 -2375 120 -2355
rect 140 -2375 160 -2355
rect 180 -2375 200 -2355
rect 220 -2375 240 -2355
rect 260 -2375 280 -2355
rect 300 -2375 320 -2355
rect 340 -2375 360 -2355
rect 380 -2375 400 -2355
rect 420 -2375 440 -2355
rect 460 -2375 480 -2355
rect 500 -2375 520 -2355
rect 540 -2375 560 -2355
rect 580 -2375 600 -2355
rect 620 -2375 640 -2355
rect 660 -2375 680 -2355
rect 700 -2375 720 -2355
rect 740 -2375 760 -2355
rect 780 -2375 800 -2355
rect 820 -2375 840 -2355
rect 860 -2375 880 -2355
rect 900 -2375 920 -2355
rect 940 -2375 960 -2355
rect 980 -2375 1000 -2355
rect 1020 -2375 1040 -2355
rect 1060 -2375 1080 -2355
rect 1100 -2375 1120 -2355
rect 1140 -2375 1160 -2355
rect 1180 -2375 1200 -2355
rect 1220 -2375 1240 -2355
rect 1260 -2375 1280 -2355
rect 1300 -2375 1320 -2355
rect 1340 -2375 1360 -2355
rect 1380 -2375 1400 -2355
rect 1420 -2375 1440 -2355
rect 1460 -2375 1480 -2355
rect 1500 -2375 1520 -2355
rect 1540 -2375 1560 -2355
rect 1580 -2375 1600 -2355
rect 1620 -2375 1640 -2355
rect 1660 -2375 1680 -2355
rect 1700 -2375 1720 -2355
rect 1740 -2375 1760 -2355
rect 1780 -2375 1800 -2355
rect 1820 -2375 1840 -2355
rect 1860 -2375 1880 -2355
rect 1900 -2375 1920 -2355
rect 1940 -2375 1960 -2355
rect 1980 -2375 2000 -2355
rect 2020 -2375 2040 -2355
rect 2060 -2375 2080 -2355
rect 2100 -2375 2120 -2355
rect 2140 -2375 2160 -2355
rect 2180 -2375 2200 -2355
rect 2220 -2375 2240 -2355
rect 2260 -2375 2280 -2355
rect 2300 -2375 2320 -2355
rect 2340 -2375 2360 -2355
rect 2380 -2375 2400 -2355
rect 2420 -2375 2440 -2355
rect 2460 -2375 2480 -2355
rect 2500 -2375 2520 -2355
rect 2540 -2375 2560 -2355
rect 2590 -2375 2605 -2355
rect 105 -2390 2605 -2375
rect 105 -2450 2605 -2435
rect 105 -2470 120 -2450
rect 140 -2470 160 -2450
rect 180 -2470 200 -2450
rect 220 -2470 240 -2450
rect 260 -2470 280 -2450
rect 300 -2470 320 -2450
rect 340 -2470 360 -2450
rect 380 -2470 400 -2450
rect 420 -2470 440 -2450
rect 460 -2470 480 -2450
rect 500 -2470 520 -2450
rect 540 -2470 560 -2450
rect 580 -2470 600 -2450
rect 620 -2470 640 -2450
rect 660 -2470 680 -2450
rect 700 -2470 720 -2450
rect 740 -2470 760 -2450
rect 780 -2470 800 -2450
rect 820 -2470 840 -2450
rect 860 -2470 880 -2450
rect 900 -2470 920 -2450
rect 940 -2470 960 -2450
rect 980 -2470 1000 -2450
rect 1020 -2470 1040 -2450
rect 1060 -2470 1080 -2450
rect 1100 -2470 1120 -2450
rect 1140 -2470 1160 -2450
rect 1180 -2470 1200 -2450
rect 1220 -2470 1240 -2450
rect 1260 -2470 1280 -2450
rect 1300 -2470 1320 -2450
rect 1340 -2470 1360 -2450
rect 1380 -2470 1400 -2450
rect 1420 -2470 1440 -2450
rect 1460 -2470 1480 -2450
rect 1500 -2470 1520 -2450
rect 1540 -2470 1560 -2450
rect 1580 -2470 1600 -2450
rect 1620 -2470 1640 -2450
rect 1660 -2470 1680 -2450
rect 1700 -2470 1720 -2450
rect 1740 -2470 1760 -2450
rect 1780 -2470 1800 -2450
rect 1820 -2470 1840 -2450
rect 1860 -2470 1880 -2450
rect 1900 -2470 1920 -2450
rect 1940 -2470 1960 -2450
rect 1980 -2470 2000 -2450
rect 2020 -2470 2040 -2450
rect 2060 -2470 2080 -2450
rect 2100 -2470 2120 -2450
rect 2140 -2470 2160 -2450
rect 2180 -2470 2200 -2450
rect 2220 -2470 2240 -2450
rect 2260 -2470 2280 -2450
rect 2300 -2470 2320 -2450
rect 2340 -2470 2360 -2450
rect 2380 -2470 2400 -2450
rect 2420 -2470 2440 -2450
rect 2460 -2470 2480 -2450
rect 2500 -2470 2520 -2450
rect 2540 -2470 2560 -2450
rect 2590 -2470 2605 -2450
rect 105 -2485 2605 -2470
rect 105 -2545 2605 -2530
rect 105 -2565 120 -2545
rect 140 -2565 160 -2545
rect 180 -2565 200 -2545
rect 220 -2565 240 -2545
rect 260 -2565 280 -2545
rect 300 -2565 320 -2545
rect 340 -2565 360 -2545
rect 380 -2565 400 -2545
rect 420 -2565 440 -2545
rect 460 -2565 480 -2545
rect 500 -2565 520 -2545
rect 540 -2565 560 -2545
rect 580 -2565 600 -2545
rect 620 -2565 640 -2545
rect 660 -2565 680 -2545
rect 700 -2565 720 -2545
rect 740 -2565 760 -2545
rect 780 -2565 800 -2545
rect 820 -2565 840 -2545
rect 860 -2565 880 -2545
rect 900 -2565 920 -2545
rect 940 -2565 960 -2545
rect 980 -2565 1000 -2545
rect 1020 -2565 1040 -2545
rect 1060 -2565 1080 -2545
rect 1100 -2565 1120 -2545
rect 1140 -2565 1160 -2545
rect 1180 -2565 1200 -2545
rect 1220 -2565 1240 -2545
rect 1260 -2565 1280 -2545
rect 1300 -2565 1320 -2545
rect 1340 -2565 1360 -2545
rect 1380 -2565 1400 -2545
rect 1420 -2565 1440 -2545
rect 1460 -2565 1480 -2545
rect 1500 -2565 1520 -2545
rect 1540 -2565 1560 -2545
rect 1580 -2565 1600 -2545
rect 1620 -2565 1640 -2545
rect 1660 -2565 1680 -2545
rect 1700 -2565 1720 -2545
rect 1740 -2565 1760 -2545
rect 1780 -2565 1800 -2545
rect 1820 -2565 1840 -2545
rect 1860 -2565 1880 -2545
rect 1900 -2565 1920 -2545
rect 1940 -2565 1960 -2545
rect 1980 -2565 2000 -2545
rect 2020 -2565 2040 -2545
rect 2060 -2565 2080 -2545
rect 2100 -2565 2120 -2545
rect 2140 -2565 2160 -2545
rect 2180 -2565 2200 -2545
rect 2220 -2565 2240 -2545
rect 2260 -2565 2280 -2545
rect 2300 -2565 2320 -2545
rect 2340 -2565 2360 -2545
rect 2380 -2565 2400 -2545
rect 2420 -2565 2440 -2545
rect 2460 -2565 2480 -2545
rect 2500 -2565 2520 -2545
rect 2540 -2565 2560 -2545
rect 2590 -2565 2605 -2545
rect 105 -2580 2605 -2565
rect 105 -2640 2605 -2625
rect 105 -2660 120 -2640
rect 140 -2660 160 -2640
rect 180 -2660 200 -2640
rect 220 -2660 240 -2640
rect 260 -2660 280 -2640
rect 300 -2660 320 -2640
rect 340 -2660 360 -2640
rect 380 -2660 400 -2640
rect 420 -2660 440 -2640
rect 460 -2660 480 -2640
rect 500 -2660 520 -2640
rect 540 -2660 560 -2640
rect 580 -2660 600 -2640
rect 620 -2660 640 -2640
rect 660 -2660 680 -2640
rect 700 -2660 720 -2640
rect 740 -2660 760 -2640
rect 780 -2660 800 -2640
rect 820 -2660 840 -2640
rect 860 -2660 880 -2640
rect 900 -2660 920 -2640
rect 940 -2660 960 -2640
rect 980 -2660 1000 -2640
rect 1020 -2660 1040 -2640
rect 1060 -2660 1080 -2640
rect 1100 -2660 1120 -2640
rect 1140 -2660 1160 -2640
rect 1180 -2660 1200 -2640
rect 1220 -2660 1240 -2640
rect 1260 -2660 1280 -2640
rect 1300 -2660 1320 -2640
rect 1340 -2660 1360 -2640
rect 1380 -2660 1400 -2640
rect 1420 -2660 1440 -2640
rect 1460 -2660 1480 -2640
rect 1500 -2660 1520 -2640
rect 1540 -2660 1560 -2640
rect 1580 -2660 1600 -2640
rect 1620 -2660 1640 -2640
rect 1660 -2660 1680 -2640
rect 1700 -2660 1720 -2640
rect 1740 -2660 1760 -2640
rect 1780 -2660 1800 -2640
rect 1820 -2660 1840 -2640
rect 1860 -2660 1880 -2640
rect 1900 -2660 1920 -2640
rect 1940 -2660 1960 -2640
rect 1980 -2660 2000 -2640
rect 2020 -2660 2040 -2640
rect 2060 -2660 2080 -2640
rect 2100 -2660 2120 -2640
rect 2140 -2660 2160 -2640
rect 2180 -2660 2200 -2640
rect 2220 -2660 2240 -2640
rect 2260 -2660 2280 -2640
rect 2300 -2660 2320 -2640
rect 2340 -2660 2360 -2640
rect 2380 -2660 2400 -2640
rect 2420 -2660 2440 -2640
rect 2460 -2660 2480 -2640
rect 2500 -2660 2520 -2640
rect 2540 -2660 2560 -2640
rect 2590 -2660 2605 -2640
rect 105 -2675 2605 -2660
rect 105 -2735 2605 -2720
rect 105 -2755 120 -2735
rect 140 -2755 160 -2735
rect 180 -2755 200 -2735
rect 220 -2755 240 -2735
rect 260 -2755 280 -2735
rect 300 -2755 320 -2735
rect 340 -2755 360 -2735
rect 380 -2755 400 -2735
rect 420 -2755 440 -2735
rect 460 -2755 480 -2735
rect 500 -2755 520 -2735
rect 540 -2755 560 -2735
rect 580 -2755 600 -2735
rect 620 -2755 640 -2735
rect 660 -2755 680 -2735
rect 700 -2755 720 -2735
rect 740 -2755 760 -2735
rect 780 -2755 800 -2735
rect 820 -2755 840 -2735
rect 860 -2755 880 -2735
rect 900 -2755 920 -2735
rect 940 -2755 960 -2735
rect 980 -2755 1000 -2735
rect 1020 -2755 1040 -2735
rect 1060 -2755 1080 -2735
rect 1100 -2755 1120 -2735
rect 1140 -2755 1160 -2735
rect 1180 -2755 1200 -2735
rect 1220 -2755 1240 -2735
rect 1260 -2755 1280 -2735
rect 1300 -2755 1320 -2735
rect 1340 -2755 1360 -2735
rect 1380 -2755 1400 -2735
rect 1420 -2755 1440 -2735
rect 1460 -2755 1480 -2735
rect 1500 -2755 1520 -2735
rect 1540 -2755 1560 -2735
rect 1580 -2755 1600 -2735
rect 1620 -2755 1640 -2735
rect 1660 -2755 1680 -2735
rect 1700 -2755 1720 -2735
rect 1740 -2755 1760 -2735
rect 1780 -2755 1800 -2735
rect 1820 -2755 1840 -2735
rect 1860 -2755 1880 -2735
rect 1900 -2755 1920 -2735
rect 1940 -2755 1960 -2735
rect 1980 -2755 2000 -2735
rect 2020 -2755 2040 -2735
rect 2060 -2755 2080 -2735
rect 2100 -2755 2120 -2735
rect 2140 -2755 2160 -2735
rect 2180 -2755 2200 -2735
rect 2220 -2755 2240 -2735
rect 2260 -2755 2280 -2735
rect 2300 -2755 2320 -2735
rect 2340 -2755 2360 -2735
rect 2380 -2755 2400 -2735
rect 2420 -2755 2440 -2735
rect 2460 -2755 2480 -2735
rect 2500 -2755 2520 -2735
rect 2540 -2755 2560 -2735
rect 2590 -2755 2605 -2735
rect 105 -2765 2605 -2755
<< ndiffc >>
rect 200 2197 220 2217
rect 240 2197 260 2217
rect 280 2197 300 2217
rect 320 2197 340 2217
rect 360 2197 380 2217
rect 400 2197 420 2217
rect 440 2197 460 2217
rect 480 2197 500 2217
rect 520 2197 540 2217
rect 560 2197 580 2217
rect 600 2197 620 2217
rect 640 2197 660 2217
rect 680 2197 700 2217
rect 720 2197 740 2217
rect 760 2197 780 2217
rect 800 2197 820 2217
rect 840 2197 860 2217
rect 880 2197 900 2217
rect 920 2197 940 2217
rect 960 2197 980 2217
rect 1000 2197 1020 2217
rect 1040 2197 1060 2217
rect 1080 2197 1100 2217
rect 1120 2197 1140 2217
rect 1160 2197 1180 2217
rect 1200 2197 1220 2217
rect 1240 2197 1260 2217
rect 1280 2197 1300 2217
rect 1320 2197 1340 2217
rect 1360 2197 1380 2217
rect 1400 2197 1420 2217
rect 1440 2197 1460 2217
rect 1480 2197 1500 2217
rect 1520 2197 1540 2217
rect 1560 2197 1580 2217
rect 1600 2197 1620 2217
rect 1640 2197 1660 2217
rect 1680 2197 1700 2217
rect 1720 2197 1740 2217
rect 1760 2197 1780 2217
rect 1800 2197 1820 2217
rect 1840 2197 1860 2217
rect 1880 2197 1900 2217
rect 1920 2197 1940 2217
rect 1960 2197 1980 2217
rect 2000 2197 2020 2217
rect 2040 2197 2060 2217
rect 2080 2197 2100 2217
rect 2120 2197 2140 2217
rect 2160 2197 2180 2217
rect 2200 2197 2220 2217
rect 2240 2197 2260 2217
rect 2280 2197 2300 2217
rect 2320 2197 2340 2217
rect 2360 2197 2380 2217
rect 2400 2197 2420 2217
rect 2440 2197 2460 2217
rect 2480 2197 2500 2217
rect 2520 2197 2540 2217
rect 2560 2197 2580 2217
rect 2600 2197 2620 2217
rect 2640 2197 2660 2217
rect 200 2115 220 2135
rect 240 2115 260 2135
rect 280 2115 300 2135
rect 320 2115 340 2135
rect 360 2115 380 2135
rect 400 2115 420 2135
rect 440 2115 460 2135
rect 480 2115 500 2135
rect 520 2115 540 2135
rect 560 2115 580 2135
rect 600 2115 620 2135
rect 640 2115 660 2135
rect 680 2115 700 2135
rect 720 2115 740 2135
rect 760 2115 780 2135
rect 800 2115 820 2135
rect 840 2115 860 2135
rect 880 2115 900 2135
rect 920 2115 940 2135
rect 960 2115 980 2135
rect 1000 2115 1020 2135
rect 1040 2115 1060 2135
rect 1080 2115 1100 2135
rect 1120 2115 1140 2135
rect 1160 2115 1180 2135
rect 1200 2115 1220 2135
rect 1240 2115 1260 2135
rect 1280 2115 1300 2135
rect 1320 2115 1340 2135
rect 1360 2115 1380 2135
rect 1400 2115 1420 2135
rect 1440 2115 1460 2135
rect 1480 2115 1500 2135
rect 1520 2115 1540 2135
rect 1560 2115 1580 2135
rect 1600 2115 1620 2135
rect 1640 2115 1660 2135
rect 1680 2115 1700 2135
rect 1720 2115 1740 2135
rect 1760 2115 1780 2135
rect 1800 2115 1820 2135
rect 1840 2115 1860 2135
rect 1880 2115 1900 2135
rect 1920 2115 1940 2135
rect 1960 2115 1980 2135
rect 2000 2115 2020 2135
rect 2040 2115 2060 2135
rect 2080 2115 2100 2135
rect 2120 2115 2140 2135
rect 2160 2115 2180 2135
rect 2200 2115 2220 2135
rect 2240 2115 2260 2135
rect 2280 2115 2300 2135
rect 2320 2115 2340 2135
rect 2360 2115 2380 2135
rect 2400 2115 2420 2135
rect 2440 2115 2460 2135
rect 2480 2115 2500 2135
rect 2520 2115 2540 2135
rect 2560 2115 2580 2135
rect 2600 2115 2620 2135
rect 2640 2115 2660 2135
rect 200 2033 220 2053
rect 240 2033 260 2053
rect 280 2033 300 2053
rect 320 2033 340 2053
rect 360 2033 380 2053
rect 400 2033 420 2053
rect 440 2033 460 2053
rect 480 2033 500 2053
rect 520 2033 540 2053
rect 560 2033 580 2053
rect 600 2033 620 2053
rect 640 2033 660 2053
rect 680 2033 700 2053
rect 720 2033 740 2053
rect 760 2033 780 2053
rect 800 2033 820 2053
rect 840 2033 860 2053
rect 880 2033 900 2053
rect 920 2033 940 2053
rect 960 2033 980 2053
rect 1000 2033 1020 2053
rect 1040 2033 1060 2053
rect 1080 2033 1100 2053
rect 1120 2033 1140 2053
rect 1160 2033 1180 2053
rect 1200 2033 1220 2053
rect 1240 2033 1260 2053
rect 1280 2033 1300 2053
rect 1320 2033 1340 2053
rect 1360 2033 1380 2053
rect 1400 2033 1420 2053
rect 1440 2033 1460 2053
rect 1480 2033 1500 2053
rect 1520 2033 1540 2053
rect 1560 2033 1580 2053
rect 1600 2033 1620 2053
rect 1640 2033 1660 2053
rect 1680 2033 1700 2053
rect 1720 2033 1740 2053
rect 1760 2033 1780 2053
rect 1800 2033 1820 2053
rect 1840 2033 1860 2053
rect 1880 2033 1900 2053
rect 1920 2033 1940 2053
rect 1960 2033 1980 2053
rect 2000 2033 2020 2053
rect 2040 2033 2060 2053
rect 2080 2033 2100 2053
rect 2120 2033 2140 2053
rect 2160 2033 2180 2053
rect 2200 2033 2220 2053
rect 2240 2033 2260 2053
rect 2280 2033 2300 2053
rect 2320 2033 2340 2053
rect 2360 2033 2380 2053
rect 2400 2033 2420 2053
rect 2440 2033 2460 2053
rect 2480 2033 2500 2053
rect 2520 2033 2540 2053
rect 2560 2033 2580 2053
rect 2600 2033 2620 2053
rect 2640 2033 2660 2053
rect 200 1951 220 1971
rect 240 1951 260 1971
rect 280 1951 300 1971
rect 320 1951 340 1971
rect 360 1951 380 1971
rect 400 1951 420 1971
rect 440 1951 460 1971
rect 480 1951 500 1971
rect 520 1951 540 1971
rect 560 1951 580 1971
rect 600 1951 620 1971
rect 640 1951 660 1971
rect 680 1951 700 1971
rect 720 1951 740 1971
rect 760 1951 780 1971
rect 800 1951 820 1971
rect 840 1951 860 1971
rect 880 1951 900 1971
rect 920 1951 940 1971
rect 960 1951 980 1971
rect 1000 1951 1020 1971
rect 1040 1951 1060 1971
rect 1080 1951 1100 1971
rect 1120 1951 1140 1971
rect 1160 1951 1180 1971
rect 1200 1951 1220 1971
rect 1240 1951 1260 1971
rect 1280 1951 1300 1971
rect 1320 1951 1340 1971
rect 1360 1951 1380 1971
rect 1400 1951 1420 1971
rect 1440 1951 1460 1971
rect 1480 1951 1500 1971
rect 1520 1951 1540 1971
rect 1560 1951 1580 1971
rect 1600 1951 1620 1971
rect 1640 1951 1660 1971
rect 1680 1951 1700 1971
rect 1720 1951 1740 1971
rect 1760 1951 1780 1971
rect 1800 1951 1820 1971
rect 1840 1951 1860 1971
rect 1880 1951 1900 1971
rect 1920 1951 1940 1971
rect 1960 1951 1980 1971
rect 2000 1951 2020 1971
rect 2040 1951 2060 1971
rect 2080 1951 2100 1971
rect 2120 1951 2140 1971
rect 2160 1951 2180 1971
rect 2200 1951 2220 1971
rect 2240 1951 2260 1971
rect 2280 1951 2300 1971
rect 2320 1951 2340 1971
rect 2360 1951 2380 1971
rect 2400 1951 2420 1971
rect 2440 1951 2460 1971
rect 2480 1951 2500 1971
rect 2520 1951 2540 1971
rect 2560 1951 2580 1971
rect 2600 1951 2620 1971
rect 2640 1951 2660 1971
rect 200 1869 220 1889
rect 240 1869 260 1889
rect 280 1869 300 1889
rect 320 1869 340 1889
rect 360 1869 380 1889
rect 400 1869 420 1889
rect 440 1869 460 1889
rect 480 1869 500 1889
rect 520 1869 540 1889
rect 560 1869 580 1889
rect 600 1869 620 1889
rect 640 1869 660 1889
rect 680 1869 700 1889
rect 720 1869 740 1889
rect 760 1869 780 1889
rect 800 1869 820 1889
rect 840 1869 860 1889
rect 880 1869 900 1889
rect 920 1869 940 1889
rect 960 1869 980 1889
rect 1000 1869 1020 1889
rect 1040 1869 1060 1889
rect 1080 1869 1100 1889
rect 1120 1869 1140 1889
rect 1160 1869 1180 1889
rect 1200 1869 1220 1889
rect 1240 1869 1260 1889
rect 1280 1869 1300 1889
rect 1320 1869 1340 1889
rect 1360 1869 1380 1889
rect 1400 1869 1420 1889
rect 1440 1869 1460 1889
rect 1480 1869 1500 1889
rect 1520 1869 1540 1889
rect 1560 1869 1580 1889
rect 1600 1869 1620 1889
rect 1640 1869 1660 1889
rect 1680 1869 1700 1889
rect 1720 1869 1740 1889
rect 1760 1869 1780 1889
rect 1800 1869 1820 1889
rect 1840 1869 1860 1889
rect 1880 1869 1900 1889
rect 1920 1869 1940 1889
rect 1960 1869 1980 1889
rect 2000 1869 2020 1889
rect 2040 1869 2060 1889
rect 2080 1869 2100 1889
rect 2120 1869 2140 1889
rect 2160 1869 2180 1889
rect 2200 1869 2220 1889
rect 2240 1869 2260 1889
rect 2280 1869 2300 1889
rect 2320 1869 2340 1889
rect 2360 1869 2380 1889
rect 2400 1869 2420 1889
rect 2440 1869 2460 1889
rect 2480 1869 2500 1889
rect 2520 1869 2540 1889
rect 2560 1869 2580 1889
rect 2600 1869 2620 1889
rect 2640 1869 2660 1889
rect 200 1787 220 1807
rect 240 1787 260 1807
rect 280 1787 300 1807
rect 320 1787 340 1807
rect 360 1787 380 1807
rect 400 1787 420 1807
rect 440 1787 460 1807
rect 480 1787 500 1807
rect 520 1787 540 1807
rect 560 1787 580 1807
rect 600 1787 620 1807
rect 640 1787 660 1807
rect 680 1787 700 1807
rect 720 1787 740 1807
rect 760 1787 780 1807
rect 800 1787 820 1807
rect 840 1787 860 1807
rect 880 1787 900 1807
rect 920 1787 940 1807
rect 960 1787 980 1807
rect 1000 1787 1020 1807
rect 1040 1787 1060 1807
rect 1080 1787 1100 1807
rect 1120 1787 1140 1807
rect 1160 1787 1180 1807
rect 1200 1787 1220 1807
rect 1240 1787 1260 1807
rect 1280 1787 1300 1807
rect 1320 1787 1340 1807
rect 1360 1787 1380 1807
rect 1400 1787 1420 1807
rect 1440 1787 1460 1807
rect 1480 1787 1500 1807
rect 1520 1787 1540 1807
rect 1560 1787 1580 1807
rect 1600 1787 1620 1807
rect 1640 1787 1660 1807
rect 1680 1787 1700 1807
rect 1720 1787 1740 1807
rect 1760 1787 1780 1807
rect 1800 1787 1820 1807
rect 1840 1787 1860 1807
rect 1880 1787 1900 1807
rect 1920 1787 1940 1807
rect 1960 1787 1980 1807
rect 2000 1787 2020 1807
rect 2040 1787 2060 1807
rect 2080 1787 2100 1807
rect 2120 1787 2140 1807
rect 2160 1787 2180 1807
rect 2200 1787 2220 1807
rect 2240 1787 2260 1807
rect 2280 1787 2300 1807
rect 2320 1787 2340 1807
rect 2360 1787 2380 1807
rect 2400 1787 2420 1807
rect 2440 1787 2460 1807
rect 2480 1787 2500 1807
rect 2520 1787 2540 1807
rect 2560 1787 2580 1807
rect 2600 1787 2620 1807
rect 2640 1787 2660 1807
rect 200 1705 220 1725
rect 240 1705 260 1725
rect 280 1705 300 1725
rect 320 1705 340 1725
rect 360 1705 380 1725
rect 400 1705 420 1725
rect 440 1705 460 1725
rect 480 1705 500 1725
rect 520 1705 540 1725
rect 560 1705 580 1725
rect 600 1705 620 1725
rect 640 1705 660 1725
rect 680 1705 700 1725
rect 720 1705 740 1725
rect 760 1705 780 1725
rect 800 1705 820 1725
rect 840 1705 860 1725
rect 880 1705 900 1725
rect 920 1705 940 1725
rect 960 1705 980 1725
rect 1000 1705 1020 1725
rect 1040 1705 1060 1725
rect 1080 1705 1100 1725
rect 1120 1705 1140 1725
rect 1160 1705 1180 1725
rect 1200 1705 1220 1725
rect 1240 1705 1260 1725
rect 1280 1705 1300 1725
rect 1320 1705 1340 1725
rect 1360 1705 1380 1725
rect 1400 1705 1420 1725
rect 1440 1705 1460 1725
rect 1480 1705 1500 1725
rect 1520 1705 1540 1725
rect 1560 1705 1580 1725
rect 1600 1705 1620 1725
rect 1640 1705 1660 1725
rect 1680 1705 1700 1725
rect 1720 1705 1740 1725
rect 1760 1705 1780 1725
rect 1800 1705 1820 1725
rect 1840 1705 1860 1725
rect 1880 1705 1900 1725
rect 1920 1705 1940 1725
rect 1960 1705 1980 1725
rect 2000 1705 2020 1725
rect 2040 1705 2060 1725
rect 2080 1705 2100 1725
rect 2120 1705 2140 1725
rect 2160 1705 2180 1725
rect 2200 1705 2220 1725
rect 2240 1705 2260 1725
rect 2280 1705 2300 1725
rect 2320 1705 2340 1725
rect 2360 1705 2380 1725
rect 2400 1705 2420 1725
rect 2440 1705 2460 1725
rect 2480 1705 2500 1725
rect 2520 1705 2540 1725
rect 2560 1705 2580 1725
rect 2600 1705 2620 1725
rect 2640 1705 2660 1725
rect 200 1623 220 1643
rect 240 1623 260 1643
rect 280 1623 300 1643
rect 320 1623 340 1643
rect 360 1623 380 1643
rect 400 1623 420 1643
rect 440 1623 460 1643
rect 480 1623 500 1643
rect 520 1623 540 1643
rect 560 1623 580 1643
rect 600 1623 620 1643
rect 640 1623 660 1643
rect 680 1623 700 1643
rect 720 1623 740 1643
rect 760 1623 780 1643
rect 800 1623 820 1643
rect 840 1623 860 1643
rect 880 1623 900 1643
rect 920 1623 940 1643
rect 960 1623 980 1643
rect 1000 1623 1020 1643
rect 1040 1623 1060 1643
rect 1080 1623 1100 1643
rect 1120 1623 1140 1643
rect 1160 1623 1180 1643
rect 1200 1623 1220 1643
rect 1240 1623 1260 1643
rect 1280 1623 1300 1643
rect 1320 1623 1340 1643
rect 1360 1623 1380 1643
rect 1400 1623 1420 1643
rect 1440 1623 1460 1643
rect 1480 1623 1500 1643
rect 1520 1623 1540 1643
rect 1560 1623 1580 1643
rect 1600 1623 1620 1643
rect 1640 1623 1660 1643
rect 1680 1623 1700 1643
rect 1720 1623 1740 1643
rect 1760 1623 1780 1643
rect 1800 1623 1820 1643
rect 1840 1623 1860 1643
rect 1880 1623 1900 1643
rect 1920 1623 1940 1643
rect 1960 1623 1980 1643
rect 2000 1623 2020 1643
rect 2040 1623 2060 1643
rect 2080 1623 2100 1643
rect 2120 1623 2140 1643
rect 2160 1623 2180 1643
rect 2200 1623 2220 1643
rect 2240 1623 2260 1643
rect 2280 1623 2300 1643
rect 2320 1623 2340 1643
rect 2360 1623 2380 1643
rect 2400 1623 2420 1643
rect 2440 1623 2460 1643
rect 2480 1623 2500 1643
rect 2520 1623 2540 1643
rect 2560 1623 2580 1643
rect 2600 1623 2620 1643
rect 2640 1623 2660 1643
rect 200 1541 220 1561
rect 240 1541 260 1561
rect 280 1541 300 1561
rect 320 1541 340 1561
rect 360 1541 380 1561
rect 400 1541 420 1561
rect 440 1541 460 1561
rect 480 1541 500 1561
rect 520 1541 540 1561
rect 560 1541 580 1561
rect 600 1541 620 1561
rect 640 1541 660 1561
rect 680 1541 700 1561
rect 720 1541 740 1561
rect 760 1541 780 1561
rect 800 1541 820 1561
rect 840 1541 860 1561
rect 880 1541 900 1561
rect 920 1541 940 1561
rect 960 1541 980 1561
rect 1000 1541 1020 1561
rect 1040 1541 1060 1561
rect 1080 1541 1100 1561
rect 1120 1541 1140 1561
rect 1160 1541 1180 1561
rect 1200 1541 1220 1561
rect 1240 1541 1260 1561
rect 1280 1541 1300 1561
rect 1320 1541 1340 1561
rect 1360 1541 1380 1561
rect 1400 1541 1420 1561
rect 1440 1541 1460 1561
rect 1480 1541 1500 1561
rect 1520 1541 1540 1561
rect 1560 1541 1580 1561
rect 1600 1541 1620 1561
rect 1640 1541 1660 1561
rect 1680 1541 1700 1561
rect 1720 1541 1740 1561
rect 1760 1541 1780 1561
rect 1800 1541 1820 1561
rect 1840 1541 1860 1561
rect 1880 1541 1900 1561
rect 1920 1541 1940 1561
rect 1960 1541 1980 1561
rect 2000 1541 2020 1561
rect 2040 1541 2060 1561
rect 2080 1541 2100 1561
rect 2120 1541 2140 1561
rect 2160 1541 2180 1561
rect 2200 1541 2220 1561
rect 2240 1541 2260 1561
rect 2280 1541 2300 1561
rect 2320 1541 2340 1561
rect 2360 1541 2380 1561
rect 2400 1541 2420 1561
rect 2440 1541 2460 1561
rect 2480 1541 2500 1561
rect 2520 1541 2540 1561
rect 2560 1541 2580 1561
rect 2600 1541 2620 1561
rect 2640 1541 2660 1561
rect 200 1459 220 1479
rect 240 1459 260 1479
rect 280 1459 300 1479
rect 320 1459 340 1479
rect 360 1459 380 1479
rect 400 1459 420 1479
rect 440 1459 460 1479
rect 480 1459 500 1479
rect 520 1459 540 1479
rect 560 1459 580 1479
rect 600 1459 620 1479
rect 640 1459 660 1479
rect 680 1459 700 1479
rect 720 1459 740 1479
rect 760 1459 780 1479
rect 800 1459 820 1479
rect 840 1459 860 1479
rect 880 1459 900 1479
rect 920 1459 940 1479
rect 960 1459 980 1479
rect 1000 1459 1020 1479
rect 1040 1459 1060 1479
rect 1080 1459 1100 1479
rect 1120 1459 1140 1479
rect 1160 1459 1180 1479
rect 1200 1459 1220 1479
rect 1240 1459 1260 1479
rect 1280 1459 1300 1479
rect 1320 1459 1340 1479
rect 1360 1459 1380 1479
rect 1400 1459 1420 1479
rect 1440 1459 1460 1479
rect 1480 1459 1500 1479
rect 1520 1459 1540 1479
rect 1560 1459 1580 1479
rect 1600 1459 1620 1479
rect 1640 1459 1660 1479
rect 1680 1459 1700 1479
rect 1720 1459 1740 1479
rect 1760 1459 1780 1479
rect 1800 1459 1820 1479
rect 1840 1459 1860 1479
rect 1880 1459 1900 1479
rect 1920 1459 1940 1479
rect 1960 1459 1980 1479
rect 2000 1459 2020 1479
rect 2040 1459 2060 1479
rect 2080 1459 2100 1479
rect 2120 1459 2140 1479
rect 2160 1459 2180 1479
rect 2200 1459 2220 1479
rect 2240 1459 2260 1479
rect 2280 1459 2300 1479
rect 2320 1459 2340 1479
rect 2360 1459 2380 1479
rect 2400 1459 2420 1479
rect 2440 1459 2460 1479
rect 2480 1459 2500 1479
rect 2520 1459 2540 1479
rect 2560 1459 2580 1479
rect 2600 1459 2620 1479
rect 2640 1459 2660 1479
rect 200 1377 220 1397
rect 240 1377 260 1397
rect 280 1377 300 1397
rect 320 1377 340 1397
rect 360 1377 380 1397
rect 400 1377 420 1397
rect 440 1377 460 1397
rect 480 1377 500 1397
rect 520 1377 540 1397
rect 560 1377 580 1397
rect 600 1377 620 1397
rect 640 1377 660 1397
rect 680 1377 700 1397
rect 720 1377 740 1397
rect 760 1377 780 1397
rect 800 1377 820 1397
rect 840 1377 860 1397
rect 880 1377 900 1397
rect 920 1377 940 1397
rect 960 1377 980 1397
rect 1000 1377 1020 1397
rect 1040 1377 1060 1397
rect 1080 1377 1100 1397
rect 1120 1377 1140 1397
rect 1160 1377 1180 1397
rect 1200 1377 1220 1397
rect 1240 1377 1260 1397
rect 1280 1377 1300 1397
rect 1320 1377 1340 1397
rect 1360 1377 1380 1397
rect 1400 1377 1420 1397
rect 1440 1377 1460 1397
rect 1480 1377 1500 1397
rect 1520 1377 1540 1397
rect 1560 1377 1580 1397
rect 1600 1377 1620 1397
rect 1640 1377 1660 1397
rect 1680 1377 1700 1397
rect 1720 1377 1740 1397
rect 1760 1377 1780 1397
rect 1800 1377 1820 1397
rect 1840 1377 1860 1397
rect 1880 1377 1900 1397
rect 1920 1377 1940 1397
rect 1960 1377 1980 1397
rect 2000 1377 2020 1397
rect 2040 1377 2060 1397
rect 2080 1377 2100 1397
rect 2120 1377 2140 1397
rect 2160 1377 2180 1397
rect 2200 1377 2220 1397
rect 2240 1377 2260 1397
rect 2280 1377 2300 1397
rect 2320 1377 2340 1397
rect 2360 1377 2380 1397
rect 2400 1377 2420 1397
rect 2440 1377 2460 1397
rect 2480 1377 2500 1397
rect 2520 1377 2540 1397
rect 2560 1377 2580 1397
rect 2600 1377 2620 1397
rect 2640 1377 2660 1397
rect 200 1295 220 1315
rect 240 1295 260 1315
rect 280 1295 300 1315
rect 320 1295 340 1315
rect 360 1295 380 1315
rect 400 1295 420 1315
rect 440 1295 460 1315
rect 480 1295 500 1315
rect 520 1295 540 1315
rect 560 1295 580 1315
rect 600 1295 620 1315
rect 640 1295 660 1315
rect 680 1295 700 1315
rect 720 1295 740 1315
rect 760 1295 780 1315
rect 800 1295 820 1315
rect 840 1295 860 1315
rect 880 1295 900 1315
rect 920 1295 940 1315
rect 960 1295 980 1315
rect 1000 1295 1020 1315
rect 1040 1295 1060 1315
rect 1080 1295 1100 1315
rect 1120 1295 1140 1315
rect 1160 1295 1180 1315
rect 1200 1295 1220 1315
rect 1240 1295 1260 1315
rect 1280 1295 1300 1315
rect 1320 1295 1340 1315
rect 1360 1295 1380 1315
rect 1400 1295 1420 1315
rect 1440 1295 1460 1315
rect 1480 1295 1500 1315
rect 1520 1295 1540 1315
rect 1560 1295 1580 1315
rect 1600 1295 1620 1315
rect 1640 1295 1660 1315
rect 1680 1295 1700 1315
rect 1720 1295 1740 1315
rect 1760 1295 1780 1315
rect 1800 1295 1820 1315
rect 1840 1295 1860 1315
rect 1880 1295 1900 1315
rect 1920 1295 1940 1315
rect 1960 1295 1980 1315
rect 2000 1295 2020 1315
rect 2040 1295 2060 1315
rect 2080 1295 2100 1315
rect 2120 1295 2140 1315
rect 2160 1295 2180 1315
rect 2200 1295 2220 1315
rect 2240 1295 2260 1315
rect 2280 1295 2300 1315
rect 2320 1295 2340 1315
rect 2360 1295 2380 1315
rect 2400 1295 2420 1315
rect 2440 1295 2460 1315
rect 2480 1295 2500 1315
rect 2520 1295 2540 1315
rect 2560 1295 2580 1315
rect 2600 1295 2620 1315
rect 2640 1295 2660 1315
rect 200 1213 220 1233
rect 240 1213 260 1233
rect 280 1213 300 1233
rect 320 1213 340 1233
rect 360 1213 380 1233
rect 400 1213 420 1233
rect 440 1213 460 1233
rect 480 1213 500 1233
rect 520 1213 540 1233
rect 560 1213 580 1233
rect 600 1213 620 1233
rect 640 1213 660 1233
rect 680 1213 700 1233
rect 720 1213 740 1233
rect 760 1213 780 1233
rect 800 1213 820 1233
rect 840 1213 860 1233
rect 880 1213 900 1233
rect 920 1213 940 1233
rect 960 1213 980 1233
rect 1000 1213 1020 1233
rect 1040 1213 1060 1233
rect 1080 1213 1100 1233
rect 1120 1213 1140 1233
rect 1160 1213 1180 1233
rect 1200 1213 1220 1233
rect 1240 1213 1260 1233
rect 1280 1213 1300 1233
rect 1320 1213 1340 1233
rect 1360 1213 1380 1233
rect 1400 1213 1420 1233
rect 1440 1213 1460 1233
rect 1480 1213 1500 1233
rect 1520 1213 1540 1233
rect 1560 1213 1580 1233
rect 1600 1213 1620 1233
rect 1640 1213 1660 1233
rect 1680 1213 1700 1233
rect 1720 1213 1740 1233
rect 1760 1213 1780 1233
rect 1800 1213 1820 1233
rect 1840 1213 1860 1233
rect 1880 1213 1900 1233
rect 1920 1213 1940 1233
rect 1960 1213 1980 1233
rect 2000 1213 2020 1233
rect 2040 1213 2060 1233
rect 2080 1213 2100 1233
rect 2120 1213 2140 1233
rect 2160 1213 2180 1233
rect 2200 1213 2220 1233
rect 2240 1213 2260 1233
rect 2280 1213 2300 1233
rect 2320 1213 2340 1233
rect 2360 1213 2380 1233
rect 2400 1213 2420 1233
rect 2440 1213 2460 1233
rect 2480 1213 2500 1233
rect 2520 1213 2540 1233
rect 2560 1213 2580 1233
rect 2600 1213 2620 1233
rect 2640 1213 2660 1233
rect 200 1131 220 1151
rect 240 1131 260 1151
rect 280 1131 300 1151
rect 320 1131 340 1151
rect 360 1131 380 1151
rect 400 1131 420 1151
rect 440 1131 460 1151
rect 480 1131 500 1151
rect 520 1131 540 1151
rect 560 1131 580 1151
rect 600 1131 620 1151
rect 640 1131 660 1151
rect 680 1131 700 1151
rect 720 1131 740 1151
rect 760 1131 780 1151
rect 800 1131 820 1151
rect 840 1131 860 1151
rect 880 1131 900 1151
rect 920 1131 940 1151
rect 960 1131 980 1151
rect 1000 1131 1020 1151
rect 1040 1131 1060 1151
rect 1080 1131 1100 1151
rect 1120 1131 1140 1151
rect 1160 1131 1180 1151
rect 1200 1131 1220 1151
rect 1240 1131 1260 1151
rect 1280 1131 1300 1151
rect 1320 1131 1340 1151
rect 1360 1131 1380 1151
rect 1400 1131 1420 1151
rect 1440 1131 1460 1151
rect 1480 1131 1500 1151
rect 1520 1131 1540 1151
rect 1560 1131 1580 1151
rect 1600 1131 1620 1151
rect 1640 1131 1660 1151
rect 1680 1131 1700 1151
rect 1720 1131 1740 1151
rect 1760 1131 1780 1151
rect 1800 1131 1820 1151
rect 1840 1131 1860 1151
rect 1880 1131 1900 1151
rect 1920 1131 1940 1151
rect 1960 1131 1980 1151
rect 2000 1131 2020 1151
rect 2040 1131 2060 1151
rect 2080 1131 2100 1151
rect 2120 1131 2140 1151
rect 2160 1131 2180 1151
rect 2200 1131 2220 1151
rect 2240 1131 2260 1151
rect 2280 1131 2300 1151
rect 2320 1131 2340 1151
rect 2360 1131 2380 1151
rect 2400 1131 2420 1151
rect 2440 1131 2460 1151
rect 2480 1131 2500 1151
rect 2520 1131 2540 1151
rect 2560 1131 2580 1151
rect 2600 1131 2620 1151
rect 2640 1131 2660 1151
rect 200 1049 220 1069
rect 240 1049 260 1069
rect 280 1049 300 1069
rect 320 1049 340 1069
rect 360 1049 380 1069
rect 400 1049 420 1069
rect 440 1049 460 1069
rect 480 1049 500 1069
rect 520 1049 540 1069
rect 560 1049 580 1069
rect 600 1049 620 1069
rect 640 1049 660 1069
rect 680 1049 700 1069
rect 720 1049 740 1069
rect 760 1049 780 1069
rect 800 1049 820 1069
rect 840 1049 860 1069
rect 880 1049 900 1069
rect 920 1049 940 1069
rect 960 1049 980 1069
rect 1000 1049 1020 1069
rect 1040 1049 1060 1069
rect 1080 1049 1100 1069
rect 1120 1049 1140 1069
rect 1160 1049 1180 1069
rect 1200 1049 1220 1069
rect 1240 1049 1260 1069
rect 1280 1049 1300 1069
rect 1320 1049 1340 1069
rect 1360 1049 1380 1069
rect 1400 1049 1420 1069
rect 1440 1049 1460 1069
rect 1480 1049 1500 1069
rect 1520 1049 1540 1069
rect 1560 1049 1580 1069
rect 1600 1049 1620 1069
rect 1640 1049 1660 1069
rect 1680 1049 1700 1069
rect 1720 1049 1740 1069
rect 1760 1049 1780 1069
rect 1800 1049 1820 1069
rect 1840 1049 1860 1069
rect 1880 1049 1900 1069
rect 1920 1049 1940 1069
rect 1960 1049 1980 1069
rect 2000 1049 2020 1069
rect 2040 1049 2060 1069
rect 2080 1049 2100 1069
rect 2120 1049 2140 1069
rect 2160 1049 2180 1069
rect 2200 1049 2220 1069
rect 2240 1049 2260 1069
rect 2280 1049 2300 1069
rect 2320 1049 2340 1069
rect 2360 1049 2380 1069
rect 2400 1049 2420 1069
rect 2440 1049 2460 1069
rect 2480 1049 2500 1069
rect 2520 1049 2540 1069
rect 2560 1049 2580 1069
rect 2600 1049 2620 1069
rect 2640 1049 2660 1069
rect 200 967 220 987
rect 240 967 260 987
rect 280 967 300 987
rect 320 967 340 987
rect 360 967 380 987
rect 400 967 420 987
rect 440 967 460 987
rect 480 967 500 987
rect 520 967 540 987
rect 560 967 580 987
rect 600 967 620 987
rect 640 967 660 987
rect 680 967 700 987
rect 720 967 740 987
rect 760 967 780 987
rect 800 967 820 987
rect 840 967 860 987
rect 880 967 900 987
rect 920 967 940 987
rect 960 967 980 987
rect 1000 967 1020 987
rect 1040 967 1060 987
rect 1080 967 1100 987
rect 1120 967 1140 987
rect 1160 967 1180 987
rect 1200 967 1220 987
rect 1240 967 1260 987
rect 1280 967 1300 987
rect 1320 967 1340 987
rect 1360 967 1380 987
rect 1400 967 1420 987
rect 1440 967 1460 987
rect 1480 967 1500 987
rect 1520 967 1540 987
rect 1560 967 1580 987
rect 1600 967 1620 987
rect 1640 967 1660 987
rect 1680 967 1700 987
rect 1720 967 1740 987
rect 1760 967 1780 987
rect 1800 967 1820 987
rect 1840 967 1860 987
rect 1880 967 1900 987
rect 1920 967 1940 987
rect 1960 967 1980 987
rect 2000 967 2020 987
rect 2040 967 2060 987
rect 2080 967 2100 987
rect 2120 967 2140 987
rect 2160 967 2180 987
rect 2200 967 2220 987
rect 2240 967 2260 987
rect 2280 967 2300 987
rect 2320 967 2340 987
rect 2360 967 2380 987
rect 2400 967 2420 987
rect 2440 967 2460 987
rect 2480 967 2500 987
rect 2520 967 2540 987
rect 2560 967 2580 987
rect 2600 967 2620 987
rect 2640 967 2660 987
rect 200 885 220 905
rect 240 885 260 905
rect 280 885 300 905
rect 320 885 340 905
rect 360 885 380 905
rect 400 885 420 905
rect 440 885 460 905
rect 480 885 500 905
rect 520 885 540 905
rect 560 885 580 905
rect 600 885 620 905
rect 640 885 660 905
rect 680 885 700 905
rect 720 885 740 905
rect 760 885 780 905
rect 800 885 820 905
rect 840 885 860 905
rect 880 885 900 905
rect 920 885 940 905
rect 960 885 980 905
rect 1000 885 1020 905
rect 1040 885 1060 905
rect 1080 885 1100 905
rect 1120 885 1140 905
rect 1160 885 1180 905
rect 1200 885 1220 905
rect 1240 885 1260 905
rect 1280 885 1300 905
rect 1320 885 1340 905
rect 1360 885 1380 905
rect 1400 885 1420 905
rect 1440 885 1460 905
rect 1480 885 1500 905
rect 1520 885 1540 905
rect 1560 885 1580 905
rect 1600 885 1620 905
rect 1640 885 1660 905
rect 1680 885 1700 905
rect 1720 885 1740 905
rect 1760 885 1780 905
rect 1800 885 1820 905
rect 1840 885 1860 905
rect 1880 885 1900 905
rect 1920 885 1940 905
rect 1960 885 1980 905
rect 2000 885 2020 905
rect 2040 885 2060 905
rect 2080 885 2100 905
rect 2120 885 2140 905
rect 2160 885 2180 905
rect 2200 885 2220 905
rect 2240 885 2260 905
rect 2280 885 2300 905
rect 2320 885 2340 905
rect 2360 885 2380 905
rect 2400 885 2420 905
rect 2440 885 2460 905
rect 2480 885 2500 905
rect 2520 885 2540 905
rect 2560 885 2580 905
rect 2600 885 2620 905
rect 2640 885 2660 905
rect 200 803 220 823
rect 240 803 260 823
rect 280 803 300 823
rect 320 803 340 823
rect 360 803 380 823
rect 400 803 420 823
rect 440 803 460 823
rect 480 803 500 823
rect 520 803 540 823
rect 560 803 580 823
rect 600 803 620 823
rect 640 803 660 823
rect 680 803 700 823
rect 720 803 740 823
rect 760 803 780 823
rect 800 803 820 823
rect 840 803 860 823
rect 880 803 900 823
rect 920 803 940 823
rect 960 803 980 823
rect 1000 803 1020 823
rect 1040 803 1060 823
rect 1080 803 1100 823
rect 1120 803 1140 823
rect 1160 803 1180 823
rect 1200 803 1220 823
rect 1240 803 1260 823
rect 1280 803 1300 823
rect 1320 803 1340 823
rect 1360 803 1380 823
rect 1400 803 1420 823
rect 1440 803 1460 823
rect 1480 803 1500 823
rect 1520 803 1540 823
rect 1560 803 1580 823
rect 1600 803 1620 823
rect 1640 803 1660 823
rect 1680 803 1700 823
rect 1720 803 1740 823
rect 1760 803 1780 823
rect 1800 803 1820 823
rect 1840 803 1860 823
rect 1880 803 1900 823
rect 1920 803 1940 823
rect 1960 803 1980 823
rect 2000 803 2020 823
rect 2040 803 2060 823
rect 2080 803 2100 823
rect 2120 803 2140 823
rect 2160 803 2180 823
rect 2200 803 2220 823
rect 2240 803 2260 823
rect 2280 803 2300 823
rect 2320 803 2340 823
rect 2360 803 2380 823
rect 2400 803 2420 823
rect 2440 803 2460 823
rect 2480 803 2500 823
rect 2520 803 2540 823
rect 2560 803 2580 823
rect 2600 803 2620 823
rect 2640 803 2660 823
rect 200 721 220 741
rect 240 721 260 741
rect 280 721 300 741
rect 320 721 340 741
rect 360 721 380 741
rect 400 721 420 741
rect 440 721 460 741
rect 480 721 500 741
rect 520 721 540 741
rect 560 721 580 741
rect 600 721 620 741
rect 640 721 660 741
rect 680 721 700 741
rect 720 721 740 741
rect 760 721 780 741
rect 800 721 820 741
rect 840 721 860 741
rect 880 721 900 741
rect 920 721 940 741
rect 960 721 980 741
rect 1000 721 1020 741
rect 1040 721 1060 741
rect 1080 721 1100 741
rect 1120 721 1140 741
rect 1160 721 1180 741
rect 1200 721 1220 741
rect 1240 721 1260 741
rect 1280 721 1300 741
rect 1320 721 1340 741
rect 1360 721 1380 741
rect 1400 721 1420 741
rect 1440 721 1460 741
rect 1480 721 1500 741
rect 1520 721 1540 741
rect 1560 721 1580 741
rect 1600 721 1620 741
rect 1640 721 1660 741
rect 1680 721 1700 741
rect 1720 721 1740 741
rect 1760 721 1780 741
rect 1800 721 1820 741
rect 1840 721 1860 741
rect 1880 721 1900 741
rect 1920 721 1940 741
rect 1960 721 1980 741
rect 2000 721 2020 741
rect 2040 721 2060 741
rect 2080 721 2100 741
rect 2120 721 2140 741
rect 2160 721 2180 741
rect 2200 721 2220 741
rect 2240 721 2260 741
rect 2280 721 2300 741
rect 2320 721 2340 741
rect 2360 721 2380 741
rect 2400 721 2420 741
rect 2440 721 2460 741
rect 2480 721 2500 741
rect 2520 721 2540 741
rect 2560 721 2580 741
rect 2600 721 2620 741
rect 2640 721 2660 741
rect 200 639 220 659
rect 240 639 260 659
rect 280 639 300 659
rect 320 639 340 659
rect 360 639 380 659
rect 400 639 420 659
rect 440 639 460 659
rect 480 639 500 659
rect 520 639 540 659
rect 560 639 580 659
rect 600 639 620 659
rect 640 639 660 659
rect 680 639 700 659
rect 720 639 740 659
rect 760 639 780 659
rect 800 639 820 659
rect 840 639 860 659
rect 880 639 900 659
rect 920 639 940 659
rect 960 639 980 659
rect 1000 639 1020 659
rect 1040 639 1060 659
rect 1080 639 1100 659
rect 1120 639 1140 659
rect 1160 639 1180 659
rect 1200 639 1220 659
rect 1240 639 1260 659
rect 1280 639 1300 659
rect 1320 639 1340 659
rect 1360 639 1380 659
rect 1400 639 1420 659
rect 1440 639 1460 659
rect 1480 639 1500 659
rect 1520 639 1540 659
rect 1560 639 1580 659
rect 1600 639 1620 659
rect 1640 639 1660 659
rect 1680 639 1700 659
rect 1720 639 1740 659
rect 1760 639 1780 659
rect 1800 639 1820 659
rect 1840 639 1860 659
rect 1880 639 1900 659
rect 1920 639 1940 659
rect 1960 639 1980 659
rect 2000 639 2020 659
rect 2040 639 2060 659
rect 2080 639 2100 659
rect 2120 639 2140 659
rect 2160 639 2180 659
rect 2200 639 2220 659
rect 2240 639 2260 659
rect 2280 639 2300 659
rect 2320 639 2340 659
rect 2360 639 2380 659
rect 2400 639 2420 659
rect 2440 639 2460 659
rect 2480 639 2500 659
rect 2520 639 2540 659
rect 2560 639 2580 659
rect 2600 639 2620 659
rect 2640 639 2660 659
rect 200 557 220 577
rect 240 557 260 577
rect 280 557 300 577
rect 320 557 340 577
rect 360 557 380 577
rect 400 557 420 577
rect 440 557 460 577
rect 480 557 500 577
rect 520 557 540 577
rect 560 557 580 577
rect 600 557 620 577
rect 640 557 660 577
rect 680 557 700 577
rect 720 557 740 577
rect 760 557 780 577
rect 800 557 820 577
rect 840 557 860 577
rect 880 557 900 577
rect 920 557 940 577
rect 960 557 980 577
rect 1000 557 1020 577
rect 1040 557 1060 577
rect 1080 557 1100 577
rect 1120 557 1140 577
rect 1160 557 1180 577
rect 1200 557 1220 577
rect 1240 557 1260 577
rect 1280 557 1300 577
rect 1320 557 1340 577
rect 1360 557 1380 577
rect 1400 557 1420 577
rect 1440 557 1460 577
rect 1480 557 1500 577
rect 1520 557 1540 577
rect 1560 557 1580 577
rect 1600 557 1620 577
rect 1640 557 1660 577
rect 1680 557 1700 577
rect 1720 557 1740 577
rect 1760 557 1780 577
rect 1800 557 1820 577
rect 1840 557 1860 577
rect 1880 557 1900 577
rect 1920 557 1940 577
rect 1960 557 1980 577
rect 2000 557 2020 577
rect 2040 557 2060 577
rect 2080 557 2100 577
rect 2120 557 2140 577
rect 2160 557 2180 577
rect 2200 557 2220 577
rect 2240 557 2260 577
rect 2280 557 2300 577
rect 2320 557 2340 577
rect 2360 557 2380 577
rect 2400 557 2420 577
rect 2440 557 2460 577
rect 2480 557 2500 577
rect 2520 557 2540 577
rect 2560 557 2580 577
rect 2600 557 2620 577
rect 2640 557 2660 577
rect 200 475 220 495
rect 240 475 260 495
rect 280 475 300 495
rect 320 475 340 495
rect 360 475 380 495
rect 400 475 420 495
rect 440 475 460 495
rect 480 475 500 495
rect 520 475 540 495
rect 560 475 580 495
rect 600 475 620 495
rect 640 475 660 495
rect 680 475 700 495
rect 720 475 740 495
rect 760 475 780 495
rect 800 475 820 495
rect 840 475 860 495
rect 880 475 900 495
rect 920 475 940 495
rect 960 475 980 495
rect 1000 475 1020 495
rect 1040 475 1060 495
rect 1080 475 1100 495
rect 1120 475 1140 495
rect 1160 475 1180 495
rect 1200 475 1220 495
rect 1240 475 1260 495
rect 1280 475 1300 495
rect 1320 475 1340 495
rect 1360 475 1380 495
rect 1400 475 1420 495
rect 1440 475 1460 495
rect 1480 475 1500 495
rect 1520 475 1540 495
rect 1560 475 1580 495
rect 1600 475 1620 495
rect 1640 475 1660 495
rect 1680 475 1700 495
rect 1720 475 1740 495
rect 1760 475 1780 495
rect 1800 475 1820 495
rect 1840 475 1860 495
rect 1880 475 1900 495
rect 1920 475 1940 495
rect 1960 475 1980 495
rect 2000 475 2020 495
rect 2040 475 2060 495
rect 2080 475 2100 495
rect 2120 475 2140 495
rect 2160 475 2180 495
rect 2200 475 2220 495
rect 2240 475 2260 495
rect 2280 475 2300 495
rect 2320 475 2340 495
rect 2360 475 2380 495
rect 2400 475 2420 495
rect 2440 475 2460 495
rect 2480 475 2500 495
rect 2520 475 2540 495
rect 2560 475 2580 495
rect 2600 475 2620 495
rect 2640 475 2660 495
rect 200 393 220 413
rect 240 393 260 413
rect 280 393 300 413
rect 320 393 340 413
rect 360 393 380 413
rect 400 393 420 413
rect 440 393 460 413
rect 480 393 500 413
rect 520 393 540 413
rect 560 393 580 413
rect 600 393 620 413
rect 640 393 660 413
rect 680 393 700 413
rect 720 393 740 413
rect 760 393 780 413
rect 800 393 820 413
rect 840 393 860 413
rect 880 393 900 413
rect 920 393 940 413
rect 960 393 980 413
rect 1000 393 1020 413
rect 1040 393 1060 413
rect 1080 393 1100 413
rect 1120 393 1140 413
rect 1160 393 1180 413
rect 1200 393 1220 413
rect 1240 393 1260 413
rect 1280 393 1300 413
rect 1320 393 1340 413
rect 1360 393 1380 413
rect 1400 393 1420 413
rect 1440 393 1460 413
rect 1480 393 1500 413
rect 1520 393 1540 413
rect 1560 393 1580 413
rect 1600 393 1620 413
rect 1640 393 1660 413
rect 1680 393 1700 413
rect 1720 393 1740 413
rect 1760 393 1780 413
rect 1800 393 1820 413
rect 1840 393 1860 413
rect 1880 393 1900 413
rect 1920 393 1940 413
rect 1960 393 1980 413
rect 2000 393 2020 413
rect 2040 393 2060 413
rect 2080 393 2100 413
rect 2120 393 2140 413
rect 2160 393 2180 413
rect 2200 393 2220 413
rect 2240 393 2260 413
rect 2280 393 2300 413
rect 2320 393 2340 413
rect 2360 393 2380 413
rect 2400 393 2420 413
rect 2440 393 2460 413
rect 2480 393 2500 413
rect 2520 393 2540 413
rect 2560 393 2580 413
rect 2600 393 2620 413
rect 2640 393 2660 413
rect 200 311 220 331
rect 240 311 260 331
rect 280 311 300 331
rect 320 311 340 331
rect 360 311 380 331
rect 400 311 420 331
rect 440 311 460 331
rect 480 311 500 331
rect 520 311 540 331
rect 560 311 580 331
rect 600 311 620 331
rect 640 311 660 331
rect 680 311 700 331
rect 720 311 740 331
rect 760 311 780 331
rect 800 311 820 331
rect 840 311 860 331
rect 880 311 900 331
rect 920 311 940 331
rect 960 311 980 331
rect 1000 311 1020 331
rect 1040 311 1060 331
rect 1080 311 1100 331
rect 1120 311 1140 331
rect 1160 311 1180 331
rect 1200 311 1220 331
rect 1240 311 1260 331
rect 1280 311 1300 331
rect 1320 311 1340 331
rect 1360 311 1380 331
rect 1400 311 1420 331
rect 1440 311 1460 331
rect 1480 311 1500 331
rect 1520 311 1540 331
rect 1560 311 1580 331
rect 1600 311 1620 331
rect 1640 311 1660 331
rect 1680 311 1700 331
rect 1720 311 1740 331
rect 1760 311 1780 331
rect 1800 311 1820 331
rect 1840 311 1860 331
rect 1880 311 1900 331
rect 1920 311 1940 331
rect 1960 311 1980 331
rect 2000 311 2020 331
rect 2040 311 2060 331
rect 2080 311 2100 331
rect 2120 311 2140 331
rect 2160 311 2180 331
rect 2200 311 2220 331
rect 2240 311 2260 331
rect 2280 311 2300 331
rect 2320 311 2340 331
rect 2360 311 2380 331
rect 2400 311 2420 331
rect 2440 311 2460 331
rect 2480 311 2500 331
rect 2520 311 2540 331
rect 2560 311 2580 331
rect 2600 311 2620 331
rect 2640 311 2660 331
rect 200 229 220 249
rect 240 229 260 249
rect 280 229 300 249
rect 320 229 340 249
rect 360 229 380 249
rect 400 229 420 249
rect 440 229 460 249
rect 480 229 500 249
rect 520 229 540 249
rect 560 229 580 249
rect 600 229 620 249
rect 640 229 660 249
rect 680 229 700 249
rect 720 229 740 249
rect 760 229 780 249
rect 800 229 820 249
rect 840 229 860 249
rect 880 229 900 249
rect 920 229 940 249
rect 960 229 980 249
rect 1000 229 1020 249
rect 1040 229 1060 249
rect 1080 229 1100 249
rect 1120 229 1140 249
rect 1160 229 1180 249
rect 1200 229 1220 249
rect 1240 229 1260 249
rect 1280 229 1300 249
rect 1320 229 1340 249
rect 1360 229 1380 249
rect 1400 229 1420 249
rect 1440 229 1460 249
rect 1480 229 1500 249
rect 1520 229 1540 249
rect 1560 229 1580 249
rect 1600 229 1620 249
rect 1640 229 1660 249
rect 1680 229 1700 249
rect 1720 229 1740 249
rect 1760 229 1780 249
rect 1800 229 1820 249
rect 1840 229 1860 249
rect 1880 229 1900 249
rect 1920 229 1940 249
rect 1960 229 1980 249
rect 2000 229 2020 249
rect 2040 229 2060 249
rect 2080 229 2100 249
rect 2120 229 2140 249
rect 2160 229 2180 249
rect 2200 229 2220 249
rect 2240 229 2260 249
rect 2280 229 2300 249
rect 2320 229 2340 249
rect 2360 229 2380 249
rect 2400 229 2420 249
rect 2440 229 2460 249
rect 2480 229 2500 249
rect 2520 229 2540 249
rect 2560 229 2580 249
rect 2600 229 2620 249
rect 2640 229 2660 249
rect 200 147 220 167
rect 240 147 260 167
rect 280 147 300 167
rect 320 147 340 167
rect 360 147 380 167
rect 400 147 420 167
rect 440 147 460 167
rect 480 147 500 167
rect 520 147 540 167
rect 560 147 580 167
rect 600 147 620 167
rect 640 147 660 167
rect 680 147 700 167
rect 720 147 740 167
rect 760 147 780 167
rect 800 147 820 167
rect 840 147 860 167
rect 880 147 900 167
rect 920 147 940 167
rect 960 147 980 167
rect 1000 147 1020 167
rect 1040 147 1060 167
rect 1080 147 1100 167
rect 1120 147 1140 167
rect 1160 147 1180 167
rect 1200 147 1220 167
rect 1240 147 1260 167
rect 1280 147 1300 167
rect 1320 147 1340 167
rect 1360 147 1380 167
rect 1400 147 1420 167
rect 1440 147 1460 167
rect 1480 147 1500 167
rect 1520 147 1540 167
rect 1560 147 1580 167
rect 1600 147 1620 167
rect 1640 147 1660 167
rect 1680 147 1700 167
rect 1720 147 1740 167
rect 1760 147 1780 167
rect 1800 147 1820 167
rect 1840 147 1860 167
rect 1880 147 1900 167
rect 1920 147 1940 167
rect 1960 147 1980 167
rect 2000 147 2020 167
rect 2040 147 2060 167
rect 2080 147 2100 167
rect 2120 147 2140 167
rect 2160 147 2180 167
rect 2200 147 2220 167
rect 2240 147 2260 167
rect 2280 147 2300 167
rect 2320 147 2340 167
rect 2360 147 2380 167
rect 2400 147 2420 167
rect 2440 147 2460 167
rect 2480 147 2500 167
rect 2520 147 2540 167
rect 2560 147 2580 167
rect 2600 147 2620 167
rect 2640 147 2660 167
rect 200 65 220 85
rect 240 65 260 85
rect 280 65 300 85
rect 320 65 340 85
rect 360 65 380 85
rect 400 65 420 85
rect 440 65 460 85
rect 480 65 500 85
rect 520 65 540 85
rect 560 65 580 85
rect 600 65 620 85
rect 640 65 660 85
rect 680 65 700 85
rect 720 65 740 85
rect 760 65 780 85
rect 800 65 820 85
rect 840 65 860 85
rect 880 65 900 85
rect 920 65 940 85
rect 960 65 980 85
rect 1000 65 1020 85
rect 1040 65 1060 85
rect 1080 65 1100 85
rect 1120 65 1140 85
rect 1160 65 1180 85
rect 1200 65 1220 85
rect 1240 65 1260 85
rect 1280 65 1300 85
rect 1320 65 1340 85
rect 1360 65 1380 85
rect 1400 65 1420 85
rect 1440 65 1460 85
rect 1480 65 1500 85
rect 1520 65 1540 85
rect 1560 65 1580 85
rect 1600 65 1620 85
rect 1640 65 1660 85
rect 1680 65 1700 85
rect 1720 65 1740 85
rect 1760 65 1780 85
rect 1800 65 1820 85
rect 1840 65 1860 85
rect 1880 65 1900 85
rect 1920 65 1940 85
rect 1960 65 1980 85
rect 2000 65 2020 85
rect 2040 65 2060 85
rect 2080 65 2100 85
rect 2120 65 2140 85
rect 2160 65 2180 85
rect 2200 65 2220 85
rect 2240 65 2260 85
rect 2280 65 2300 85
rect 2320 65 2340 85
rect 2360 65 2380 85
rect 2400 65 2420 85
rect 2440 65 2460 85
rect 2480 65 2500 85
rect 2520 65 2540 85
rect 2560 65 2580 85
rect 2600 65 2620 85
rect 2640 65 2660 85
rect 120 -285 140 -265
rect 160 -285 180 -265
rect 200 -285 220 -265
rect 240 -285 260 -265
rect 280 -285 300 -265
rect 320 -285 340 -265
rect 360 -285 380 -265
rect 400 -285 420 -265
rect 440 -285 460 -265
rect 480 -285 500 -265
rect 520 -285 540 -265
rect 560 -285 580 -265
rect 600 -285 620 -265
rect 640 -285 660 -265
rect 680 -285 700 -265
rect 720 -285 740 -265
rect 760 -285 780 -265
rect 800 -285 820 -265
rect 840 -285 860 -265
rect 880 -285 900 -265
rect 920 -285 940 -265
rect 960 -285 980 -265
rect 1000 -285 1020 -265
rect 1040 -285 1060 -265
rect 1080 -285 1100 -265
rect 1120 -285 1140 -265
rect 1160 -285 1180 -265
rect 1200 -285 1220 -265
rect 1240 -285 1260 -265
rect 1280 -285 1300 -265
rect 1320 -285 1340 -265
rect 1360 -285 1380 -265
rect 1400 -285 1420 -265
rect 1440 -285 1460 -265
rect 1480 -285 1500 -265
rect 1520 -285 1540 -265
rect 1560 -285 1580 -265
rect 1600 -285 1620 -265
rect 1640 -285 1660 -265
rect 1680 -285 1700 -265
rect 1720 -285 1740 -265
rect 1760 -285 1780 -265
rect 1800 -285 1820 -265
rect 1840 -285 1860 -265
rect 1880 -285 1900 -265
rect 1920 -285 1940 -265
rect 1960 -285 1980 -265
rect 2000 -285 2020 -265
rect 2040 -285 2060 -265
rect 2080 -285 2100 -265
rect 2120 -285 2140 -265
rect 2160 -285 2180 -265
rect 2200 -285 2220 -265
rect 2240 -285 2260 -265
rect 2280 -285 2300 -265
rect 2320 -285 2340 -265
rect 2360 -285 2380 -265
rect 2400 -285 2420 -265
rect 2440 -285 2460 -265
rect 2480 -285 2500 -265
rect 2520 -285 2540 -265
rect 2560 -285 2590 -265
rect 120 -380 140 -360
rect 160 -380 180 -360
rect 200 -380 220 -360
rect 240 -380 260 -360
rect 280 -380 300 -360
rect 320 -380 340 -360
rect 360 -380 380 -360
rect 400 -380 420 -360
rect 440 -380 460 -360
rect 480 -380 500 -360
rect 520 -380 540 -360
rect 560 -380 580 -360
rect 600 -380 620 -360
rect 640 -380 660 -360
rect 680 -380 700 -360
rect 720 -380 740 -360
rect 760 -380 780 -360
rect 800 -380 820 -360
rect 840 -380 860 -360
rect 880 -380 900 -360
rect 920 -380 940 -360
rect 960 -380 980 -360
rect 1000 -380 1020 -360
rect 1040 -380 1060 -360
rect 1080 -380 1100 -360
rect 1120 -380 1140 -360
rect 1160 -380 1180 -360
rect 1200 -380 1220 -360
rect 1240 -380 1260 -360
rect 1280 -380 1300 -360
rect 1320 -380 1340 -360
rect 1360 -380 1380 -360
rect 1400 -380 1420 -360
rect 1440 -380 1460 -360
rect 1480 -380 1500 -360
rect 1520 -380 1540 -360
rect 1560 -380 1580 -360
rect 1600 -380 1620 -360
rect 1640 -380 1660 -360
rect 1680 -380 1700 -360
rect 1720 -380 1740 -360
rect 1760 -380 1780 -360
rect 1800 -380 1820 -360
rect 1840 -380 1860 -360
rect 1880 -380 1900 -360
rect 1920 -380 1940 -360
rect 1960 -380 1980 -360
rect 2000 -380 2020 -360
rect 2040 -380 2060 -360
rect 2080 -380 2100 -360
rect 2120 -380 2140 -360
rect 2160 -380 2180 -360
rect 2200 -380 2220 -360
rect 2240 -380 2260 -360
rect 2280 -380 2300 -360
rect 2320 -380 2340 -360
rect 2360 -380 2380 -360
rect 2400 -380 2420 -360
rect 2440 -380 2460 -360
rect 2480 -380 2500 -360
rect 2520 -380 2540 -360
rect 2560 -380 2590 -360
rect 120 -475 140 -455
rect 160 -475 180 -455
rect 200 -475 220 -455
rect 240 -475 260 -455
rect 280 -475 300 -455
rect 320 -475 340 -455
rect 360 -475 380 -455
rect 400 -475 420 -455
rect 440 -475 460 -455
rect 480 -475 500 -455
rect 520 -475 540 -455
rect 560 -475 580 -455
rect 600 -475 620 -455
rect 640 -475 660 -455
rect 680 -475 700 -455
rect 720 -475 740 -455
rect 760 -475 780 -455
rect 800 -475 820 -455
rect 840 -475 860 -455
rect 880 -475 900 -455
rect 920 -475 940 -455
rect 960 -475 980 -455
rect 1000 -475 1020 -455
rect 1040 -475 1060 -455
rect 1080 -475 1100 -455
rect 1120 -475 1140 -455
rect 1160 -475 1180 -455
rect 1200 -475 1220 -455
rect 1240 -475 1260 -455
rect 1280 -475 1300 -455
rect 1320 -475 1340 -455
rect 1360 -475 1380 -455
rect 1400 -475 1420 -455
rect 1440 -475 1460 -455
rect 1480 -475 1500 -455
rect 1520 -475 1540 -455
rect 1560 -475 1580 -455
rect 1600 -475 1620 -455
rect 1640 -475 1660 -455
rect 1680 -475 1700 -455
rect 1720 -475 1740 -455
rect 1760 -475 1780 -455
rect 1800 -475 1820 -455
rect 1840 -475 1860 -455
rect 1880 -475 1900 -455
rect 1920 -475 1940 -455
rect 1960 -475 1980 -455
rect 2000 -475 2020 -455
rect 2040 -475 2060 -455
rect 2080 -475 2100 -455
rect 2120 -475 2140 -455
rect 2160 -475 2180 -455
rect 2200 -475 2220 -455
rect 2240 -475 2260 -455
rect 2280 -475 2300 -455
rect 2320 -475 2340 -455
rect 2360 -475 2380 -455
rect 2400 -475 2420 -455
rect 2440 -475 2460 -455
rect 2480 -475 2500 -455
rect 2520 -475 2540 -455
rect 2560 -475 2590 -455
rect 120 -570 140 -550
rect 160 -570 180 -550
rect 200 -570 220 -550
rect 240 -570 260 -550
rect 280 -570 300 -550
rect 320 -570 340 -550
rect 360 -570 380 -550
rect 400 -570 420 -550
rect 440 -570 460 -550
rect 480 -570 500 -550
rect 520 -570 540 -550
rect 560 -570 580 -550
rect 600 -570 620 -550
rect 640 -570 660 -550
rect 680 -570 700 -550
rect 720 -570 740 -550
rect 760 -570 780 -550
rect 800 -570 820 -550
rect 840 -570 860 -550
rect 880 -570 900 -550
rect 920 -570 940 -550
rect 960 -570 980 -550
rect 1000 -570 1020 -550
rect 1040 -570 1060 -550
rect 1080 -570 1100 -550
rect 1120 -570 1140 -550
rect 1160 -570 1180 -550
rect 1200 -570 1220 -550
rect 1240 -570 1260 -550
rect 1280 -570 1300 -550
rect 1320 -570 1340 -550
rect 1360 -570 1380 -550
rect 1400 -570 1420 -550
rect 1440 -570 1460 -550
rect 1480 -570 1500 -550
rect 1520 -570 1540 -550
rect 1560 -570 1580 -550
rect 1600 -570 1620 -550
rect 1640 -570 1660 -550
rect 1680 -570 1700 -550
rect 1720 -570 1740 -550
rect 1760 -570 1780 -550
rect 1800 -570 1820 -550
rect 1840 -570 1860 -550
rect 1880 -570 1900 -550
rect 1920 -570 1940 -550
rect 1960 -570 1980 -550
rect 2000 -570 2020 -550
rect 2040 -570 2060 -550
rect 2080 -570 2100 -550
rect 2120 -570 2140 -550
rect 2160 -570 2180 -550
rect 2200 -570 2220 -550
rect 2240 -570 2260 -550
rect 2280 -570 2300 -550
rect 2320 -570 2340 -550
rect 2360 -570 2380 -550
rect 2400 -570 2420 -550
rect 2440 -570 2460 -550
rect 2480 -570 2500 -550
rect 2520 -570 2540 -550
rect 2560 -570 2590 -550
rect 120 -665 140 -645
rect 160 -665 180 -645
rect 200 -665 220 -645
rect 240 -665 260 -645
rect 280 -665 300 -645
rect 320 -665 340 -645
rect 360 -665 380 -645
rect 400 -665 420 -645
rect 440 -665 460 -645
rect 480 -665 500 -645
rect 520 -665 540 -645
rect 560 -665 580 -645
rect 600 -665 620 -645
rect 640 -665 660 -645
rect 680 -665 700 -645
rect 720 -665 740 -645
rect 760 -665 780 -645
rect 800 -665 820 -645
rect 840 -665 860 -645
rect 880 -665 900 -645
rect 920 -665 940 -645
rect 960 -665 980 -645
rect 1000 -665 1020 -645
rect 1040 -665 1060 -645
rect 1080 -665 1100 -645
rect 1120 -665 1140 -645
rect 1160 -665 1180 -645
rect 1200 -665 1220 -645
rect 1240 -665 1260 -645
rect 1280 -665 1300 -645
rect 1320 -665 1340 -645
rect 1360 -665 1380 -645
rect 1400 -665 1420 -645
rect 1440 -665 1460 -645
rect 1480 -665 1500 -645
rect 1520 -665 1540 -645
rect 1560 -665 1580 -645
rect 1600 -665 1620 -645
rect 1640 -665 1660 -645
rect 1680 -665 1700 -645
rect 1720 -665 1740 -645
rect 1760 -665 1780 -645
rect 1800 -665 1820 -645
rect 1840 -665 1860 -645
rect 1880 -665 1900 -645
rect 1920 -665 1940 -645
rect 1960 -665 1980 -645
rect 2000 -665 2020 -645
rect 2040 -665 2060 -645
rect 2080 -665 2100 -645
rect 2120 -665 2140 -645
rect 2160 -665 2180 -645
rect 2200 -665 2220 -645
rect 2240 -665 2260 -645
rect 2280 -665 2300 -645
rect 2320 -665 2340 -645
rect 2360 -665 2380 -645
rect 2400 -665 2420 -645
rect 2440 -665 2460 -645
rect 2480 -665 2500 -645
rect 2520 -665 2540 -645
rect 2560 -665 2590 -645
rect 120 -760 140 -740
rect 160 -760 180 -740
rect 200 -760 220 -740
rect 240 -760 260 -740
rect 280 -760 300 -740
rect 320 -760 340 -740
rect 360 -760 380 -740
rect 400 -760 420 -740
rect 440 -760 460 -740
rect 480 -760 500 -740
rect 520 -760 540 -740
rect 560 -760 580 -740
rect 600 -760 620 -740
rect 640 -760 660 -740
rect 680 -760 700 -740
rect 720 -760 740 -740
rect 760 -760 780 -740
rect 800 -760 820 -740
rect 840 -760 860 -740
rect 880 -760 900 -740
rect 920 -760 940 -740
rect 960 -760 980 -740
rect 1000 -760 1020 -740
rect 1040 -760 1060 -740
rect 1080 -760 1100 -740
rect 1120 -760 1140 -740
rect 1160 -760 1180 -740
rect 1200 -760 1220 -740
rect 1240 -760 1260 -740
rect 1280 -760 1300 -740
rect 1320 -760 1340 -740
rect 1360 -760 1380 -740
rect 1400 -760 1420 -740
rect 1440 -760 1460 -740
rect 1480 -760 1500 -740
rect 1520 -760 1540 -740
rect 1560 -760 1580 -740
rect 1600 -760 1620 -740
rect 1640 -760 1660 -740
rect 1680 -760 1700 -740
rect 1720 -760 1740 -740
rect 1760 -760 1780 -740
rect 1800 -760 1820 -740
rect 1840 -760 1860 -740
rect 1880 -760 1900 -740
rect 1920 -760 1940 -740
rect 1960 -760 1980 -740
rect 2000 -760 2020 -740
rect 2040 -760 2060 -740
rect 2080 -760 2100 -740
rect 2120 -760 2140 -740
rect 2160 -760 2180 -740
rect 2200 -760 2220 -740
rect 2240 -760 2260 -740
rect 2280 -760 2300 -740
rect 2320 -760 2340 -740
rect 2360 -760 2380 -740
rect 2400 -760 2420 -740
rect 2440 -760 2460 -740
rect 2480 -760 2500 -740
rect 2520 -760 2540 -740
rect 2560 -760 2590 -740
rect 120 -855 140 -835
rect 160 -855 180 -835
rect 200 -855 220 -835
rect 240 -855 260 -835
rect 280 -855 300 -835
rect 320 -855 340 -835
rect 360 -855 380 -835
rect 400 -855 420 -835
rect 440 -855 460 -835
rect 480 -855 500 -835
rect 520 -855 540 -835
rect 560 -855 580 -835
rect 600 -855 620 -835
rect 640 -855 660 -835
rect 680 -855 700 -835
rect 720 -855 740 -835
rect 760 -855 780 -835
rect 800 -855 820 -835
rect 840 -855 860 -835
rect 880 -855 900 -835
rect 920 -855 940 -835
rect 960 -855 980 -835
rect 1000 -855 1020 -835
rect 1040 -855 1060 -835
rect 1080 -855 1100 -835
rect 1120 -855 1140 -835
rect 1160 -855 1180 -835
rect 1200 -855 1220 -835
rect 1240 -855 1260 -835
rect 1280 -855 1300 -835
rect 1320 -855 1340 -835
rect 1360 -855 1380 -835
rect 1400 -855 1420 -835
rect 1440 -855 1460 -835
rect 1480 -855 1500 -835
rect 1520 -855 1540 -835
rect 1560 -855 1580 -835
rect 1600 -855 1620 -835
rect 1640 -855 1660 -835
rect 1680 -855 1700 -835
rect 1720 -855 1740 -835
rect 1760 -855 1780 -835
rect 1800 -855 1820 -835
rect 1840 -855 1860 -835
rect 1880 -855 1900 -835
rect 1920 -855 1940 -835
rect 1960 -855 1980 -835
rect 2000 -855 2020 -835
rect 2040 -855 2060 -835
rect 2080 -855 2100 -835
rect 2120 -855 2140 -835
rect 2160 -855 2180 -835
rect 2200 -855 2220 -835
rect 2240 -855 2260 -835
rect 2280 -855 2300 -835
rect 2320 -855 2340 -835
rect 2360 -855 2380 -835
rect 2400 -855 2420 -835
rect 2440 -855 2460 -835
rect 2480 -855 2500 -835
rect 2520 -855 2540 -835
rect 2560 -855 2590 -835
rect 120 -950 140 -930
rect 160 -950 180 -930
rect 200 -950 220 -930
rect 240 -950 260 -930
rect 280 -950 300 -930
rect 320 -950 340 -930
rect 360 -950 380 -930
rect 400 -950 420 -930
rect 440 -950 460 -930
rect 480 -950 500 -930
rect 520 -950 540 -930
rect 560 -950 580 -930
rect 600 -950 620 -930
rect 640 -950 660 -930
rect 680 -950 700 -930
rect 720 -950 740 -930
rect 760 -950 780 -930
rect 800 -950 820 -930
rect 840 -950 860 -930
rect 880 -950 900 -930
rect 920 -950 940 -930
rect 960 -950 980 -930
rect 1000 -950 1020 -930
rect 1040 -950 1060 -930
rect 1080 -950 1100 -930
rect 1120 -950 1140 -930
rect 1160 -950 1180 -930
rect 1200 -950 1220 -930
rect 1240 -950 1260 -930
rect 1280 -950 1300 -930
rect 1320 -950 1340 -930
rect 1360 -950 1380 -930
rect 1400 -950 1420 -930
rect 1440 -950 1460 -930
rect 1480 -950 1500 -930
rect 1520 -950 1540 -930
rect 1560 -950 1580 -930
rect 1600 -950 1620 -930
rect 1640 -950 1660 -930
rect 1680 -950 1700 -930
rect 1720 -950 1740 -930
rect 1760 -950 1780 -930
rect 1800 -950 1820 -930
rect 1840 -950 1860 -930
rect 1880 -950 1900 -930
rect 1920 -950 1940 -930
rect 1960 -950 1980 -930
rect 2000 -950 2020 -930
rect 2040 -950 2060 -930
rect 2080 -950 2100 -930
rect 2120 -950 2140 -930
rect 2160 -950 2180 -930
rect 2200 -950 2220 -930
rect 2240 -950 2260 -930
rect 2280 -950 2300 -930
rect 2320 -950 2340 -930
rect 2360 -950 2380 -930
rect 2400 -950 2420 -930
rect 2440 -950 2460 -930
rect 2480 -950 2500 -930
rect 2520 -950 2540 -930
rect 2560 -950 2590 -930
rect 120 -1045 140 -1025
rect 160 -1045 180 -1025
rect 200 -1045 220 -1025
rect 240 -1045 260 -1025
rect 280 -1045 300 -1025
rect 320 -1045 340 -1025
rect 360 -1045 380 -1025
rect 400 -1045 420 -1025
rect 440 -1045 460 -1025
rect 480 -1045 500 -1025
rect 520 -1045 540 -1025
rect 560 -1045 580 -1025
rect 600 -1045 620 -1025
rect 640 -1045 660 -1025
rect 680 -1045 700 -1025
rect 720 -1045 740 -1025
rect 760 -1045 780 -1025
rect 800 -1045 820 -1025
rect 840 -1045 860 -1025
rect 880 -1045 900 -1025
rect 920 -1045 940 -1025
rect 960 -1045 980 -1025
rect 1000 -1045 1020 -1025
rect 1040 -1045 1060 -1025
rect 1080 -1045 1100 -1025
rect 1120 -1045 1140 -1025
rect 1160 -1045 1180 -1025
rect 1200 -1045 1220 -1025
rect 1240 -1045 1260 -1025
rect 1280 -1045 1300 -1025
rect 1320 -1045 1340 -1025
rect 1360 -1045 1380 -1025
rect 1400 -1045 1420 -1025
rect 1440 -1045 1460 -1025
rect 1480 -1045 1500 -1025
rect 1520 -1045 1540 -1025
rect 1560 -1045 1580 -1025
rect 1600 -1045 1620 -1025
rect 1640 -1045 1660 -1025
rect 1680 -1045 1700 -1025
rect 1720 -1045 1740 -1025
rect 1760 -1045 1780 -1025
rect 1800 -1045 1820 -1025
rect 1840 -1045 1860 -1025
rect 1880 -1045 1900 -1025
rect 1920 -1045 1940 -1025
rect 1960 -1045 1980 -1025
rect 2000 -1045 2020 -1025
rect 2040 -1045 2060 -1025
rect 2080 -1045 2100 -1025
rect 2120 -1045 2140 -1025
rect 2160 -1045 2180 -1025
rect 2200 -1045 2220 -1025
rect 2240 -1045 2260 -1025
rect 2280 -1045 2300 -1025
rect 2320 -1045 2340 -1025
rect 2360 -1045 2380 -1025
rect 2400 -1045 2420 -1025
rect 2440 -1045 2460 -1025
rect 2480 -1045 2500 -1025
rect 2520 -1045 2540 -1025
rect 2560 -1045 2590 -1025
rect 120 -1140 140 -1120
rect 160 -1140 180 -1120
rect 200 -1140 220 -1120
rect 240 -1140 260 -1120
rect 280 -1140 300 -1120
rect 320 -1140 340 -1120
rect 360 -1140 380 -1120
rect 400 -1140 420 -1120
rect 440 -1140 460 -1120
rect 480 -1140 500 -1120
rect 520 -1140 540 -1120
rect 560 -1140 580 -1120
rect 600 -1140 620 -1120
rect 640 -1140 660 -1120
rect 680 -1140 700 -1120
rect 720 -1140 740 -1120
rect 760 -1140 780 -1120
rect 800 -1140 820 -1120
rect 840 -1140 860 -1120
rect 880 -1140 900 -1120
rect 920 -1140 940 -1120
rect 960 -1140 980 -1120
rect 1000 -1140 1020 -1120
rect 1040 -1140 1060 -1120
rect 1080 -1140 1100 -1120
rect 1120 -1140 1140 -1120
rect 1160 -1140 1180 -1120
rect 1200 -1140 1220 -1120
rect 1240 -1140 1260 -1120
rect 1280 -1140 1300 -1120
rect 1320 -1140 1340 -1120
rect 1360 -1140 1380 -1120
rect 1400 -1140 1420 -1120
rect 1440 -1140 1460 -1120
rect 1480 -1140 1500 -1120
rect 1520 -1140 1540 -1120
rect 1560 -1140 1580 -1120
rect 1600 -1140 1620 -1120
rect 1640 -1140 1660 -1120
rect 1680 -1140 1700 -1120
rect 1720 -1140 1740 -1120
rect 1760 -1140 1780 -1120
rect 1800 -1140 1820 -1120
rect 1840 -1140 1860 -1120
rect 1880 -1140 1900 -1120
rect 1920 -1140 1940 -1120
rect 1960 -1140 1980 -1120
rect 2000 -1140 2020 -1120
rect 2040 -1140 2060 -1120
rect 2080 -1140 2100 -1120
rect 2120 -1140 2140 -1120
rect 2160 -1140 2180 -1120
rect 2200 -1140 2220 -1120
rect 2240 -1140 2260 -1120
rect 2280 -1140 2300 -1120
rect 2320 -1140 2340 -1120
rect 2360 -1140 2380 -1120
rect 2400 -1140 2420 -1120
rect 2440 -1140 2460 -1120
rect 2480 -1140 2500 -1120
rect 2520 -1140 2540 -1120
rect 2560 -1140 2590 -1120
rect 120 -1235 140 -1215
rect 160 -1235 180 -1215
rect 200 -1235 220 -1215
rect 240 -1235 260 -1215
rect 280 -1235 300 -1215
rect 320 -1235 340 -1215
rect 360 -1235 380 -1215
rect 400 -1235 420 -1215
rect 440 -1235 460 -1215
rect 480 -1235 500 -1215
rect 520 -1235 540 -1215
rect 560 -1235 580 -1215
rect 600 -1235 620 -1215
rect 640 -1235 660 -1215
rect 680 -1235 700 -1215
rect 720 -1235 740 -1215
rect 760 -1235 780 -1215
rect 800 -1235 820 -1215
rect 840 -1235 860 -1215
rect 880 -1235 900 -1215
rect 920 -1235 940 -1215
rect 960 -1235 980 -1215
rect 1000 -1235 1020 -1215
rect 1040 -1235 1060 -1215
rect 1080 -1235 1100 -1215
rect 1120 -1235 1140 -1215
rect 1160 -1235 1180 -1215
rect 1200 -1235 1220 -1215
rect 1240 -1235 1260 -1215
rect 1280 -1235 1300 -1215
rect 1320 -1235 1340 -1215
rect 1360 -1235 1380 -1215
rect 1400 -1235 1420 -1215
rect 1440 -1235 1460 -1215
rect 1480 -1235 1500 -1215
rect 1520 -1235 1540 -1215
rect 1560 -1235 1580 -1215
rect 1600 -1235 1620 -1215
rect 1640 -1235 1660 -1215
rect 1680 -1235 1700 -1215
rect 1720 -1235 1740 -1215
rect 1760 -1235 1780 -1215
rect 1800 -1235 1820 -1215
rect 1840 -1235 1860 -1215
rect 1880 -1235 1900 -1215
rect 1920 -1235 1940 -1215
rect 1960 -1235 1980 -1215
rect 2000 -1235 2020 -1215
rect 2040 -1235 2060 -1215
rect 2080 -1235 2100 -1215
rect 2120 -1235 2140 -1215
rect 2160 -1235 2180 -1215
rect 2200 -1235 2220 -1215
rect 2240 -1235 2260 -1215
rect 2280 -1235 2300 -1215
rect 2320 -1235 2340 -1215
rect 2360 -1235 2380 -1215
rect 2400 -1235 2420 -1215
rect 2440 -1235 2460 -1215
rect 2480 -1235 2500 -1215
rect 2520 -1235 2540 -1215
rect 2560 -1235 2590 -1215
rect 120 -1330 140 -1310
rect 160 -1330 180 -1310
rect 200 -1330 220 -1310
rect 240 -1330 260 -1310
rect 280 -1330 300 -1310
rect 320 -1330 340 -1310
rect 360 -1330 380 -1310
rect 400 -1330 420 -1310
rect 440 -1330 460 -1310
rect 480 -1330 500 -1310
rect 520 -1330 540 -1310
rect 560 -1330 580 -1310
rect 600 -1330 620 -1310
rect 640 -1330 660 -1310
rect 680 -1330 700 -1310
rect 720 -1330 740 -1310
rect 760 -1330 780 -1310
rect 800 -1330 820 -1310
rect 840 -1330 860 -1310
rect 880 -1330 900 -1310
rect 920 -1330 940 -1310
rect 960 -1330 980 -1310
rect 1000 -1330 1020 -1310
rect 1040 -1330 1060 -1310
rect 1080 -1330 1100 -1310
rect 1120 -1330 1140 -1310
rect 1160 -1330 1180 -1310
rect 1200 -1330 1220 -1310
rect 1240 -1330 1260 -1310
rect 1280 -1330 1300 -1310
rect 1320 -1330 1340 -1310
rect 1360 -1330 1380 -1310
rect 1400 -1330 1420 -1310
rect 1440 -1330 1460 -1310
rect 1480 -1330 1500 -1310
rect 1520 -1330 1540 -1310
rect 1560 -1330 1580 -1310
rect 1600 -1330 1620 -1310
rect 1640 -1330 1660 -1310
rect 1680 -1330 1700 -1310
rect 1720 -1330 1740 -1310
rect 1760 -1330 1780 -1310
rect 1800 -1330 1820 -1310
rect 1840 -1330 1860 -1310
rect 1880 -1330 1900 -1310
rect 1920 -1330 1940 -1310
rect 1960 -1330 1980 -1310
rect 2000 -1330 2020 -1310
rect 2040 -1330 2060 -1310
rect 2080 -1330 2100 -1310
rect 2120 -1330 2140 -1310
rect 2160 -1330 2180 -1310
rect 2200 -1330 2220 -1310
rect 2240 -1330 2260 -1310
rect 2280 -1330 2300 -1310
rect 2320 -1330 2340 -1310
rect 2360 -1330 2380 -1310
rect 2400 -1330 2420 -1310
rect 2440 -1330 2460 -1310
rect 2480 -1330 2500 -1310
rect 2520 -1330 2540 -1310
rect 2560 -1330 2590 -1310
rect 120 -1425 140 -1405
rect 160 -1425 180 -1405
rect 200 -1425 220 -1405
rect 240 -1425 260 -1405
rect 280 -1425 300 -1405
rect 320 -1425 340 -1405
rect 360 -1425 380 -1405
rect 400 -1425 420 -1405
rect 440 -1425 460 -1405
rect 480 -1425 500 -1405
rect 520 -1425 540 -1405
rect 560 -1425 580 -1405
rect 600 -1425 620 -1405
rect 640 -1425 660 -1405
rect 680 -1425 700 -1405
rect 720 -1425 740 -1405
rect 760 -1425 780 -1405
rect 800 -1425 820 -1405
rect 840 -1425 860 -1405
rect 880 -1425 900 -1405
rect 920 -1425 940 -1405
rect 960 -1425 980 -1405
rect 1000 -1425 1020 -1405
rect 1040 -1425 1060 -1405
rect 1080 -1425 1100 -1405
rect 1120 -1425 1140 -1405
rect 1160 -1425 1180 -1405
rect 1200 -1425 1220 -1405
rect 1240 -1425 1260 -1405
rect 1280 -1425 1300 -1405
rect 1320 -1425 1340 -1405
rect 1360 -1425 1380 -1405
rect 1400 -1425 1420 -1405
rect 1440 -1425 1460 -1405
rect 1480 -1425 1500 -1405
rect 1520 -1425 1540 -1405
rect 1560 -1425 1580 -1405
rect 1600 -1425 1620 -1405
rect 1640 -1425 1660 -1405
rect 1680 -1425 1700 -1405
rect 1720 -1425 1740 -1405
rect 1760 -1425 1780 -1405
rect 1800 -1425 1820 -1405
rect 1840 -1425 1860 -1405
rect 1880 -1425 1900 -1405
rect 1920 -1425 1940 -1405
rect 1960 -1425 1980 -1405
rect 2000 -1425 2020 -1405
rect 2040 -1425 2060 -1405
rect 2080 -1425 2100 -1405
rect 2120 -1425 2140 -1405
rect 2160 -1425 2180 -1405
rect 2200 -1425 2220 -1405
rect 2240 -1425 2260 -1405
rect 2280 -1425 2300 -1405
rect 2320 -1425 2340 -1405
rect 2360 -1425 2380 -1405
rect 2400 -1425 2420 -1405
rect 2440 -1425 2460 -1405
rect 2480 -1425 2500 -1405
rect 2520 -1425 2540 -1405
rect 2560 -1425 2590 -1405
rect 120 -1520 140 -1500
rect 160 -1520 180 -1500
rect 200 -1520 220 -1500
rect 240 -1520 260 -1500
rect 280 -1520 300 -1500
rect 320 -1520 340 -1500
rect 360 -1520 380 -1500
rect 400 -1520 420 -1500
rect 440 -1520 460 -1500
rect 480 -1520 500 -1500
rect 520 -1520 540 -1500
rect 560 -1520 580 -1500
rect 600 -1520 620 -1500
rect 640 -1520 660 -1500
rect 680 -1520 700 -1500
rect 720 -1520 740 -1500
rect 760 -1520 780 -1500
rect 800 -1520 820 -1500
rect 840 -1520 860 -1500
rect 880 -1520 900 -1500
rect 920 -1520 940 -1500
rect 960 -1520 980 -1500
rect 1000 -1520 1020 -1500
rect 1040 -1520 1060 -1500
rect 1080 -1520 1100 -1500
rect 1120 -1520 1140 -1500
rect 1160 -1520 1180 -1500
rect 1200 -1520 1220 -1500
rect 1240 -1520 1260 -1500
rect 1280 -1520 1300 -1500
rect 1320 -1520 1340 -1500
rect 1360 -1520 1380 -1500
rect 1400 -1520 1420 -1500
rect 1440 -1520 1460 -1500
rect 1480 -1520 1500 -1500
rect 1520 -1520 1540 -1500
rect 1560 -1520 1580 -1500
rect 1600 -1520 1620 -1500
rect 1640 -1520 1660 -1500
rect 1680 -1520 1700 -1500
rect 1720 -1520 1740 -1500
rect 1760 -1520 1780 -1500
rect 1800 -1520 1820 -1500
rect 1840 -1520 1860 -1500
rect 1880 -1520 1900 -1500
rect 1920 -1520 1940 -1500
rect 1960 -1520 1980 -1500
rect 2000 -1520 2020 -1500
rect 2040 -1520 2060 -1500
rect 2080 -1520 2100 -1500
rect 2120 -1520 2140 -1500
rect 2160 -1520 2180 -1500
rect 2200 -1520 2220 -1500
rect 2240 -1520 2260 -1500
rect 2280 -1520 2300 -1500
rect 2320 -1520 2340 -1500
rect 2360 -1520 2380 -1500
rect 2400 -1520 2420 -1500
rect 2440 -1520 2460 -1500
rect 2480 -1520 2500 -1500
rect 2520 -1520 2540 -1500
rect 2560 -1520 2590 -1500
rect 120 -1615 140 -1595
rect 160 -1615 180 -1595
rect 200 -1615 220 -1595
rect 240 -1615 260 -1595
rect 280 -1615 300 -1595
rect 320 -1615 340 -1595
rect 360 -1615 380 -1595
rect 400 -1615 420 -1595
rect 440 -1615 460 -1595
rect 480 -1615 500 -1595
rect 520 -1615 540 -1595
rect 560 -1615 580 -1595
rect 600 -1615 620 -1595
rect 640 -1615 660 -1595
rect 680 -1615 700 -1595
rect 720 -1615 740 -1595
rect 760 -1615 780 -1595
rect 800 -1615 820 -1595
rect 840 -1615 860 -1595
rect 880 -1615 900 -1595
rect 920 -1615 940 -1595
rect 960 -1615 980 -1595
rect 1000 -1615 1020 -1595
rect 1040 -1615 1060 -1595
rect 1080 -1615 1100 -1595
rect 1120 -1615 1140 -1595
rect 1160 -1615 1180 -1595
rect 1200 -1615 1220 -1595
rect 1240 -1615 1260 -1595
rect 1280 -1615 1300 -1595
rect 1320 -1615 1340 -1595
rect 1360 -1615 1380 -1595
rect 1400 -1615 1420 -1595
rect 1440 -1615 1460 -1595
rect 1480 -1615 1500 -1595
rect 1520 -1615 1540 -1595
rect 1560 -1615 1580 -1595
rect 1600 -1615 1620 -1595
rect 1640 -1615 1660 -1595
rect 1680 -1615 1700 -1595
rect 1720 -1615 1740 -1595
rect 1760 -1615 1780 -1595
rect 1800 -1615 1820 -1595
rect 1840 -1615 1860 -1595
rect 1880 -1615 1900 -1595
rect 1920 -1615 1940 -1595
rect 1960 -1615 1980 -1595
rect 2000 -1615 2020 -1595
rect 2040 -1615 2060 -1595
rect 2080 -1615 2100 -1595
rect 2120 -1615 2140 -1595
rect 2160 -1615 2180 -1595
rect 2200 -1615 2220 -1595
rect 2240 -1615 2260 -1595
rect 2280 -1615 2300 -1595
rect 2320 -1615 2340 -1595
rect 2360 -1615 2380 -1595
rect 2400 -1615 2420 -1595
rect 2440 -1615 2460 -1595
rect 2480 -1615 2500 -1595
rect 2520 -1615 2540 -1595
rect 2560 -1615 2590 -1595
rect 120 -1710 140 -1690
rect 160 -1710 180 -1690
rect 200 -1710 220 -1690
rect 240 -1710 260 -1690
rect 280 -1710 300 -1690
rect 320 -1710 340 -1690
rect 360 -1710 380 -1690
rect 400 -1710 420 -1690
rect 440 -1710 460 -1690
rect 480 -1710 500 -1690
rect 520 -1710 540 -1690
rect 560 -1710 580 -1690
rect 600 -1710 620 -1690
rect 640 -1710 660 -1690
rect 680 -1710 700 -1690
rect 720 -1710 740 -1690
rect 760 -1710 780 -1690
rect 800 -1710 820 -1690
rect 840 -1710 860 -1690
rect 880 -1710 900 -1690
rect 920 -1710 940 -1690
rect 960 -1710 980 -1690
rect 1000 -1710 1020 -1690
rect 1040 -1710 1060 -1690
rect 1080 -1710 1100 -1690
rect 1120 -1710 1140 -1690
rect 1160 -1710 1180 -1690
rect 1200 -1710 1220 -1690
rect 1240 -1710 1260 -1690
rect 1280 -1710 1300 -1690
rect 1320 -1710 1340 -1690
rect 1360 -1710 1380 -1690
rect 1400 -1710 1420 -1690
rect 1440 -1710 1460 -1690
rect 1480 -1710 1500 -1690
rect 1520 -1710 1540 -1690
rect 1560 -1710 1580 -1690
rect 1600 -1710 1620 -1690
rect 1640 -1710 1660 -1690
rect 1680 -1710 1700 -1690
rect 1720 -1710 1740 -1690
rect 1760 -1710 1780 -1690
rect 1800 -1710 1820 -1690
rect 1840 -1710 1860 -1690
rect 1880 -1710 1900 -1690
rect 1920 -1710 1940 -1690
rect 1960 -1710 1980 -1690
rect 2000 -1710 2020 -1690
rect 2040 -1710 2060 -1690
rect 2080 -1710 2100 -1690
rect 2120 -1710 2140 -1690
rect 2160 -1710 2180 -1690
rect 2200 -1710 2220 -1690
rect 2240 -1710 2260 -1690
rect 2280 -1710 2300 -1690
rect 2320 -1710 2340 -1690
rect 2360 -1710 2380 -1690
rect 2400 -1710 2420 -1690
rect 2440 -1710 2460 -1690
rect 2480 -1710 2500 -1690
rect 2520 -1710 2540 -1690
rect 2560 -1710 2590 -1690
rect 120 -1805 140 -1785
rect 160 -1805 180 -1785
rect 200 -1805 220 -1785
rect 240 -1805 260 -1785
rect 280 -1805 300 -1785
rect 320 -1805 340 -1785
rect 360 -1805 380 -1785
rect 400 -1805 420 -1785
rect 440 -1805 460 -1785
rect 480 -1805 500 -1785
rect 520 -1805 540 -1785
rect 560 -1805 580 -1785
rect 600 -1805 620 -1785
rect 640 -1805 660 -1785
rect 680 -1805 700 -1785
rect 720 -1805 740 -1785
rect 760 -1805 780 -1785
rect 800 -1805 820 -1785
rect 840 -1805 860 -1785
rect 880 -1805 900 -1785
rect 920 -1805 940 -1785
rect 960 -1805 980 -1785
rect 1000 -1805 1020 -1785
rect 1040 -1805 1060 -1785
rect 1080 -1805 1100 -1785
rect 1120 -1805 1140 -1785
rect 1160 -1805 1180 -1785
rect 1200 -1805 1220 -1785
rect 1240 -1805 1260 -1785
rect 1280 -1805 1300 -1785
rect 1320 -1805 1340 -1785
rect 1360 -1805 1380 -1785
rect 1400 -1805 1420 -1785
rect 1440 -1805 1460 -1785
rect 1480 -1805 1500 -1785
rect 1520 -1805 1540 -1785
rect 1560 -1805 1580 -1785
rect 1600 -1805 1620 -1785
rect 1640 -1805 1660 -1785
rect 1680 -1805 1700 -1785
rect 1720 -1805 1740 -1785
rect 1760 -1805 1780 -1785
rect 1800 -1805 1820 -1785
rect 1840 -1805 1860 -1785
rect 1880 -1805 1900 -1785
rect 1920 -1805 1940 -1785
rect 1960 -1805 1980 -1785
rect 2000 -1805 2020 -1785
rect 2040 -1805 2060 -1785
rect 2080 -1805 2100 -1785
rect 2120 -1805 2140 -1785
rect 2160 -1805 2180 -1785
rect 2200 -1805 2220 -1785
rect 2240 -1805 2260 -1785
rect 2280 -1805 2300 -1785
rect 2320 -1805 2340 -1785
rect 2360 -1805 2380 -1785
rect 2400 -1805 2420 -1785
rect 2440 -1805 2460 -1785
rect 2480 -1805 2500 -1785
rect 2520 -1805 2540 -1785
rect 2560 -1805 2590 -1785
rect 120 -1900 140 -1880
rect 160 -1900 180 -1880
rect 200 -1900 220 -1880
rect 240 -1900 260 -1880
rect 280 -1900 300 -1880
rect 320 -1900 340 -1880
rect 360 -1900 380 -1880
rect 400 -1900 420 -1880
rect 440 -1900 460 -1880
rect 480 -1900 500 -1880
rect 520 -1900 540 -1880
rect 560 -1900 580 -1880
rect 600 -1900 620 -1880
rect 640 -1900 660 -1880
rect 680 -1900 700 -1880
rect 720 -1900 740 -1880
rect 760 -1900 780 -1880
rect 800 -1900 820 -1880
rect 840 -1900 860 -1880
rect 880 -1900 900 -1880
rect 920 -1900 940 -1880
rect 960 -1900 980 -1880
rect 1000 -1900 1020 -1880
rect 1040 -1900 1060 -1880
rect 1080 -1900 1100 -1880
rect 1120 -1900 1140 -1880
rect 1160 -1900 1180 -1880
rect 1200 -1900 1220 -1880
rect 1240 -1900 1260 -1880
rect 1280 -1900 1300 -1880
rect 1320 -1900 1340 -1880
rect 1360 -1900 1380 -1880
rect 1400 -1900 1420 -1880
rect 1440 -1900 1460 -1880
rect 1480 -1900 1500 -1880
rect 1520 -1900 1540 -1880
rect 1560 -1900 1580 -1880
rect 1600 -1900 1620 -1880
rect 1640 -1900 1660 -1880
rect 1680 -1900 1700 -1880
rect 1720 -1900 1740 -1880
rect 1760 -1900 1780 -1880
rect 1800 -1900 1820 -1880
rect 1840 -1900 1860 -1880
rect 1880 -1900 1900 -1880
rect 1920 -1900 1940 -1880
rect 1960 -1900 1980 -1880
rect 2000 -1900 2020 -1880
rect 2040 -1900 2060 -1880
rect 2080 -1900 2100 -1880
rect 2120 -1900 2140 -1880
rect 2160 -1900 2180 -1880
rect 2200 -1900 2220 -1880
rect 2240 -1900 2260 -1880
rect 2280 -1900 2300 -1880
rect 2320 -1900 2340 -1880
rect 2360 -1900 2380 -1880
rect 2400 -1900 2420 -1880
rect 2440 -1900 2460 -1880
rect 2480 -1900 2500 -1880
rect 2520 -1900 2540 -1880
rect 2560 -1900 2590 -1880
rect 120 -1995 140 -1975
rect 160 -1995 180 -1975
rect 200 -1995 220 -1975
rect 240 -1995 260 -1975
rect 280 -1995 300 -1975
rect 320 -1995 340 -1975
rect 360 -1995 380 -1975
rect 400 -1995 420 -1975
rect 440 -1995 460 -1975
rect 480 -1995 500 -1975
rect 520 -1995 540 -1975
rect 560 -1995 580 -1975
rect 600 -1995 620 -1975
rect 640 -1995 660 -1975
rect 680 -1995 700 -1975
rect 720 -1995 740 -1975
rect 760 -1995 780 -1975
rect 800 -1995 820 -1975
rect 840 -1995 860 -1975
rect 880 -1995 900 -1975
rect 920 -1995 940 -1975
rect 960 -1995 980 -1975
rect 1000 -1995 1020 -1975
rect 1040 -1995 1060 -1975
rect 1080 -1995 1100 -1975
rect 1120 -1995 1140 -1975
rect 1160 -1995 1180 -1975
rect 1200 -1995 1220 -1975
rect 1240 -1995 1260 -1975
rect 1280 -1995 1300 -1975
rect 1320 -1995 1340 -1975
rect 1360 -1995 1380 -1975
rect 1400 -1995 1420 -1975
rect 1440 -1995 1460 -1975
rect 1480 -1995 1500 -1975
rect 1520 -1995 1540 -1975
rect 1560 -1995 1580 -1975
rect 1600 -1995 1620 -1975
rect 1640 -1995 1660 -1975
rect 1680 -1995 1700 -1975
rect 1720 -1995 1740 -1975
rect 1760 -1995 1780 -1975
rect 1800 -1995 1820 -1975
rect 1840 -1995 1860 -1975
rect 1880 -1995 1900 -1975
rect 1920 -1995 1940 -1975
rect 1960 -1995 1980 -1975
rect 2000 -1995 2020 -1975
rect 2040 -1995 2060 -1975
rect 2080 -1995 2100 -1975
rect 2120 -1995 2140 -1975
rect 2160 -1995 2180 -1975
rect 2200 -1995 2220 -1975
rect 2240 -1995 2260 -1975
rect 2280 -1995 2300 -1975
rect 2320 -1995 2340 -1975
rect 2360 -1995 2380 -1975
rect 2400 -1995 2420 -1975
rect 2440 -1995 2460 -1975
rect 2480 -1995 2500 -1975
rect 2520 -1995 2540 -1975
rect 2560 -1995 2590 -1975
rect 120 -2090 140 -2070
rect 160 -2090 180 -2070
rect 200 -2090 220 -2070
rect 240 -2090 260 -2070
rect 280 -2090 300 -2070
rect 320 -2090 340 -2070
rect 360 -2090 380 -2070
rect 400 -2090 420 -2070
rect 440 -2090 460 -2070
rect 480 -2090 500 -2070
rect 520 -2090 540 -2070
rect 560 -2090 580 -2070
rect 600 -2090 620 -2070
rect 640 -2090 660 -2070
rect 680 -2090 700 -2070
rect 720 -2090 740 -2070
rect 760 -2090 780 -2070
rect 800 -2090 820 -2070
rect 840 -2090 860 -2070
rect 880 -2090 900 -2070
rect 920 -2090 940 -2070
rect 960 -2090 980 -2070
rect 1000 -2090 1020 -2070
rect 1040 -2090 1060 -2070
rect 1080 -2090 1100 -2070
rect 1120 -2090 1140 -2070
rect 1160 -2090 1180 -2070
rect 1200 -2090 1220 -2070
rect 1240 -2090 1260 -2070
rect 1280 -2090 1300 -2070
rect 1320 -2090 1340 -2070
rect 1360 -2090 1380 -2070
rect 1400 -2090 1420 -2070
rect 1440 -2090 1460 -2070
rect 1480 -2090 1500 -2070
rect 1520 -2090 1540 -2070
rect 1560 -2090 1580 -2070
rect 1600 -2090 1620 -2070
rect 1640 -2090 1660 -2070
rect 1680 -2090 1700 -2070
rect 1720 -2090 1740 -2070
rect 1760 -2090 1780 -2070
rect 1800 -2090 1820 -2070
rect 1840 -2090 1860 -2070
rect 1880 -2090 1900 -2070
rect 1920 -2090 1940 -2070
rect 1960 -2090 1980 -2070
rect 2000 -2090 2020 -2070
rect 2040 -2090 2060 -2070
rect 2080 -2090 2100 -2070
rect 2120 -2090 2140 -2070
rect 2160 -2090 2180 -2070
rect 2200 -2090 2220 -2070
rect 2240 -2090 2260 -2070
rect 2280 -2090 2300 -2070
rect 2320 -2090 2340 -2070
rect 2360 -2090 2380 -2070
rect 2400 -2090 2420 -2070
rect 2440 -2090 2460 -2070
rect 2480 -2090 2500 -2070
rect 2520 -2090 2540 -2070
rect 2560 -2090 2590 -2070
rect 120 -2185 140 -2165
rect 160 -2185 180 -2165
rect 200 -2185 220 -2165
rect 240 -2185 260 -2165
rect 280 -2185 300 -2165
rect 320 -2185 340 -2165
rect 360 -2185 380 -2165
rect 400 -2185 420 -2165
rect 440 -2185 460 -2165
rect 480 -2185 500 -2165
rect 520 -2185 540 -2165
rect 560 -2185 580 -2165
rect 600 -2185 620 -2165
rect 640 -2185 660 -2165
rect 680 -2185 700 -2165
rect 720 -2185 740 -2165
rect 760 -2185 780 -2165
rect 800 -2185 820 -2165
rect 840 -2185 860 -2165
rect 880 -2185 900 -2165
rect 920 -2185 940 -2165
rect 960 -2185 980 -2165
rect 1000 -2185 1020 -2165
rect 1040 -2185 1060 -2165
rect 1080 -2185 1100 -2165
rect 1120 -2185 1140 -2165
rect 1160 -2185 1180 -2165
rect 1200 -2185 1220 -2165
rect 1240 -2185 1260 -2165
rect 1280 -2185 1300 -2165
rect 1320 -2185 1340 -2165
rect 1360 -2185 1380 -2165
rect 1400 -2185 1420 -2165
rect 1440 -2185 1460 -2165
rect 1480 -2185 1500 -2165
rect 1520 -2185 1540 -2165
rect 1560 -2185 1580 -2165
rect 1600 -2185 1620 -2165
rect 1640 -2185 1660 -2165
rect 1680 -2185 1700 -2165
rect 1720 -2185 1740 -2165
rect 1760 -2185 1780 -2165
rect 1800 -2185 1820 -2165
rect 1840 -2185 1860 -2165
rect 1880 -2185 1900 -2165
rect 1920 -2185 1940 -2165
rect 1960 -2185 1980 -2165
rect 2000 -2185 2020 -2165
rect 2040 -2185 2060 -2165
rect 2080 -2185 2100 -2165
rect 2120 -2185 2140 -2165
rect 2160 -2185 2180 -2165
rect 2200 -2185 2220 -2165
rect 2240 -2185 2260 -2165
rect 2280 -2185 2300 -2165
rect 2320 -2185 2340 -2165
rect 2360 -2185 2380 -2165
rect 2400 -2185 2420 -2165
rect 2440 -2185 2460 -2165
rect 2480 -2185 2500 -2165
rect 2520 -2185 2540 -2165
rect 2560 -2185 2590 -2165
rect 120 -2280 140 -2260
rect 160 -2280 180 -2260
rect 200 -2280 220 -2260
rect 240 -2280 260 -2260
rect 280 -2280 300 -2260
rect 320 -2280 340 -2260
rect 360 -2280 380 -2260
rect 400 -2280 420 -2260
rect 440 -2280 460 -2260
rect 480 -2280 500 -2260
rect 520 -2280 540 -2260
rect 560 -2280 580 -2260
rect 600 -2280 620 -2260
rect 640 -2280 660 -2260
rect 680 -2280 700 -2260
rect 720 -2280 740 -2260
rect 760 -2280 780 -2260
rect 800 -2280 820 -2260
rect 840 -2280 860 -2260
rect 880 -2280 900 -2260
rect 920 -2280 940 -2260
rect 960 -2280 980 -2260
rect 1000 -2280 1020 -2260
rect 1040 -2280 1060 -2260
rect 1080 -2280 1100 -2260
rect 1120 -2280 1140 -2260
rect 1160 -2280 1180 -2260
rect 1200 -2280 1220 -2260
rect 1240 -2280 1260 -2260
rect 1280 -2280 1300 -2260
rect 1320 -2280 1340 -2260
rect 1360 -2280 1380 -2260
rect 1400 -2280 1420 -2260
rect 1440 -2280 1460 -2260
rect 1480 -2280 1500 -2260
rect 1520 -2280 1540 -2260
rect 1560 -2280 1580 -2260
rect 1600 -2280 1620 -2260
rect 1640 -2280 1660 -2260
rect 1680 -2280 1700 -2260
rect 1720 -2280 1740 -2260
rect 1760 -2280 1780 -2260
rect 1800 -2280 1820 -2260
rect 1840 -2280 1860 -2260
rect 1880 -2280 1900 -2260
rect 1920 -2280 1940 -2260
rect 1960 -2280 1980 -2260
rect 2000 -2280 2020 -2260
rect 2040 -2280 2060 -2260
rect 2080 -2280 2100 -2260
rect 2120 -2280 2140 -2260
rect 2160 -2280 2180 -2260
rect 2200 -2280 2220 -2260
rect 2240 -2280 2260 -2260
rect 2280 -2280 2300 -2260
rect 2320 -2280 2340 -2260
rect 2360 -2280 2380 -2260
rect 2400 -2280 2420 -2260
rect 2440 -2280 2460 -2260
rect 2480 -2280 2500 -2260
rect 2520 -2280 2540 -2260
rect 2560 -2280 2590 -2260
rect 120 -2375 140 -2355
rect 160 -2375 180 -2355
rect 200 -2375 220 -2355
rect 240 -2375 260 -2355
rect 280 -2375 300 -2355
rect 320 -2375 340 -2355
rect 360 -2375 380 -2355
rect 400 -2375 420 -2355
rect 440 -2375 460 -2355
rect 480 -2375 500 -2355
rect 520 -2375 540 -2355
rect 560 -2375 580 -2355
rect 600 -2375 620 -2355
rect 640 -2375 660 -2355
rect 680 -2375 700 -2355
rect 720 -2375 740 -2355
rect 760 -2375 780 -2355
rect 800 -2375 820 -2355
rect 840 -2375 860 -2355
rect 880 -2375 900 -2355
rect 920 -2375 940 -2355
rect 960 -2375 980 -2355
rect 1000 -2375 1020 -2355
rect 1040 -2375 1060 -2355
rect 1080 -2375 1100 -2355
rect 1120 -2375 1140 -2355
rect 1160 -2375 1180 -2355
rect 1200 -2375 1220 -2355
rect 1240 -2375 1260 -2355
rect 1280 -2375 1300 -2355
rect 1320 -2375 1340 -2355
rect 1360 -2375 1380 -2355
rect 1400 -2375 1420 -2355
rect 1440 -2375 1460 -2355
rect 1480 -2375 1500 -2355
rect 1520 -2375 1540 -2355
rect 1560 -2375 1580 -2355
rect 1600 -2375 1620 -2355
rect 1640 -2375 1660 -2355
rect 1680 -2375 1700 -2355
rect 1720 -2375 1740 -2355
rect 1760 -2375 1780 -2355
rect 1800 -2375 1820 -2355
rect 1840 -2375 1860 -2355
rect 1880 -2375 1900 -2355
rect 1920 -2375 1940 -2355
rect 1960 -2375 1980 -2355
rect 2000 -2375 2020 -2355
rect 2040 -2375 2060 -2355
rect 2080 -2375 2100 -2355
rect 2120 -2375 2140 -2355
rect 2160 -2375 2180 -2355
rect 2200 -2375 2220 -2355
rect 2240 -2375 2260 -2355
rect 2280 -2375 2300 -2355
rect 2320 -2375 2340 -2355
rect 2360 -2375 2380 -2355
rect 2400 -2375 2420 -2355
rect 2440 -2375 2460 -2355
rect 2480 -2375 2500 -2355
rect 2520 -2375 2540 -2355
rect 2560 -2375 2590 -2355
rect 120 -2470 140 -2450
rect 160 -2470 180 -2450
rect 200 -2470 220 -2450
rect 240 -2470 260 -2450
rect 280 -2470 300 -2450
rect 320 -2470 340 -2450
rect 360 -2470 380 -2450
rect 400 -2470 420 -2450
rect 440 -2470 460 -2450
rect 480 -2470 500 -2450
rect 520 -2470 540 -2450
rect 560 -2470 580 -2450
rect 600 -2470 620 -2450
rect 640 -2470 660 -2450
rect 680 -2470 700 -2450
rect 720 -2470 740 -2450
rect 760 -2470 780 -2450
rect 800 -2470 820 -2450
rect 840 -2470 860 -2450
rect 880 -2470 900 -2450
rect 920 -2470 940 -2450
rect 960 -2470 980 -2450
rect 1000 -2470 1020 -2450
rect 1040 -2470 1060 -2450
rect 1080 -2470 1100 -2450
rect 1120 -2470 1140 -2450
rect 1160 -2470 1180 -2450
rect 1200 -2470 1220 -2450
rect 1240 -2470 1260 -2450
rect 1280 -2470 1300 -2450
rect 1320 -2470 1340 -2450
rect 1360 -2470 1380 -2450
rect 1400 -2470 1420 -2450
rect 1440 -2470 1460 -2450
rect 1480 -2470 1500 -2450
rect 1520 -2470 1540 -2450
rect 1560 -2470 1580 -2450
rect 1600 -2470 1620 -2450
rect 1640 -2470 1660 -2450
rect 1680 -2470 1700 -2450
rect 1720 -2470 1740 -2450
rect 1760 -2470 1780 -2450
rect 1800 -2470 1820 -2450
rect 1840 -2470 1860 -2450
rect 1880 -2470 1900 -2450
rect 1920 -2470 1940 -2450
rect 1960 -2470 1980 -2450
rect 2000 -2470 2020 -2450
rect 2040 -2470 2060 -2450
rect 2080 -2470 2100 -2450
rect 2120 -2470 2140 -2450
rect 2160 -2470 2180 -2450
rect 2200 -2470 2220 -2450
rect 2240 -2470 2260 -2450
rect 2280 -2470 2300 -2450
rect 2320 -2470 2340 -2450
rect 2360 -2470 2380 -2450
rect 2400 -2470 2420 -2450
rect 2440 -2470 2460 -2450
rect 2480 -2470 2500 -2450
rect 2520 -2470 2540 -2450
rect 2560 -2470 2590 -2450
rect 120 -2565 140 -2545
rect 160 -2565 180 -2545
rect 200 -2565 220 -2545
rect 240 -2565 260 -2545
rect 280 -2565 300 -2545
rect 320 -2565 340 -2545
rect 360 -2565 380 -2545
rect 400 -2565 420 -2545
rect 440 -2565 460 -2545
rect 480 -2565 500 -2545
rect 520 -2565 540 -2545
rect 560 -2565 580 -2545
rect 600 -2565 620 -2545
rect 640 -2565 660 -2545
rect 680 -2565 700 -2545
rect 720 -2565 740 -2545
rect 760 -2565 780 -2545
rect 800 -2565 820 -2545
rect 840 -2565 860 -2545
rect 880 -2565 900 -2545
rect 920 -2565 940 -2545
rect 960 -2565 980 -2545
rect 1000 -2565 1020 -2545
rect 1040 -2565 1060 -2545
rect 1080 -2565 1100 -2545
rect 1120 -2565 1140 -2545
rect 1160 -2565 1180 -2545
rect 1200 -2565 1220 -2545
rect 1240 -2565 1260 -2545
rect 1280 -2565 1300 -2545
rect 1320 -2565 1340 -2545
rect 1360 -2565 1380 -2545
rect 1400 -2565 1420 -2545
rect 1440 -2565 1460 -2545
rect 1480 -2565 1500 -2545
rect 1520 -2565 1540 -2545
rect 1560 -2565 1580 -2545
rect 1600 -2565 1620 -2545
rect 1640 -2565 1660 -2545
rect 1680 -2565 1700 -2545
rect 1720 -2565 1740 -2545
rect 1760 -2565 1780 -2545
rect 1800 -2565 1820 -2545
rect 1840 -2565 1860 -2545
rect 1880 -2565 1900 -2545
rect 1920 -2565 1940 -2545
rect 1960 -2565 1980 -2545
rect 2000 -2565 2020 -2545
rect 2040 -2565 2060 -2545
rect 2080 -2565 2100 -2545
rect 2120 -2565 2140 -2545
rect 2160 -2565 2180 -2545
rect 2200 -2565 2220 -2545
rect 2240 -2565 2260 -2545
rect 2280 -2565 2300 -2545
rect 2320 -2565 2340 -2545
rect 2360 -2565 2380 -2545
rect 2400 -2565 2420 -2545
rect 2440 -2565 2460 -2545
rect 2480 -2565 2500 -2545
rect 2520 -2565 2540 -2545
rect 2560 -2565 2590 -2545
rect 120 -2660 140 -2640
rect 160 -2660 180 -2640
rect 200 -2660 220 -2640
rect 240 -2660 260 -2640
rect 280 -2660 300 -2640
rect 320 -2660 340 -2640
rect 360 -2660 380 -2640
rect 400 -2660 420 -2640
rect 440 -2660 460 -2640
rect 480 -2660 500 -2640
rect 520 -2660 540 -2640
rect 560 -2660 580 -2640
rect 600 -2660 620 -2640
rect 640 -2660 660 -2640
rect 680 -2660 700 -2640
rect 720 -2660 740 -2640
rect 760 -2660 780 -2640
rect 800 -2660 820 -2640
rect 840 -2660 860 -2640
rect 880 -2660 900 -2640
rect 920 -2660 940 -2640
rect 960 -2660 980 -2640
rect 1000 -2660 1020 -2640
rect 1040 -2660 1060 -2640
rect 1080 -2660 1100 -2640
rect 1120 -2660 1140 -2640
rect 1160 -2660 1180 -2640
rect 1200 -2660 1220 -2640
rect 1240 -2660 1260 -2640
rect 1280 -2660 1300 -2640
rect 1320 -2660 1340 -2640
rect 1360 -2660 1380 -2640
rect 1400 -2660 1420 -2640
rect 1440 -2660 1460 -2640
rect 1480 -2660 1500 -2640
rect 1520 -2660 1540 -2640
rect 1560 -2660 1580 -2640
rect 1600 -2660 1620 -2640
rect 1640 -2660 1660 -2640
rect 1680 -2660 1700 -2640
rect 1720 -2660 1740 -2640
rect 1760 -2660 1780 -2640
rect 1800 -2660 1820 -2640
rect 1840 -2660 1860 -2640
rect 1880 -2660 1900 -2640
rect 1920 -2660 1940 -2640
rect 1960 -2660 1980 -2640
rect 2000 -2660 2020 -2640
rect 2040 -2660 2060 -2640
rect 2080 -2660 2100 -2640
rect 2120 -2660 2140 -2640
rect 2160 -2660 2180 -2640
rect 2200 -2660 2220 -2640
rect 2240 -2660 2260 -2640
rect 2280 -2660 2300 -2640
rect 2320 -2660 2340 -2640
rect 2360 -2660 2380 -2640
rect 2400 -2660 2420 -2640
rect 2440 -2660 2460 -2640
rect 2480 -2660 2500 -2640
rect 2520 -2660 2540 -2640
rect 2560 -2660 2590 -2640
rect 120 -2755 140 -2735
rect 160 -2755 180 -2735
rect 200 -2755 220 -2735
rect 240 -2755 260 -2735
rect 280 -2755 300 -2735
rect 320 -2755 340 -2735
rect 360 -2755 380 -2735
rect 400 -2755 420 -2735
rect 440 -2755 460 -2735
rect 480 -2755 500 -2735
rect 520 -2755 540 -2735
rect 560 -2755 580 -2735
rect 600 -2755 620 -2735
rect 640 -2755 660 -2735
rect 680 -2755 700 -2735
rect 720 -2755 740 -2735
rect 760 -2755 780 -2735
rect 800 -2755 820 -2735
rect 840 -2755 860 -2735
rect 880 -2755 900 -2735
rect 920 -2755 940 -2735
rect 960 -2755 980 -2735
rect 1000 -2755 1020 -2735
rect 1040 -2755 1060 -2735
rect 1080 -2755 1100 -2735
rect 1120 -2755 1140 -2735
rect 1160 -2755 1180 -2735
rect 1200 -2755 1220 -2735
rect 1240 -2755 1260 -2735
rect 1280 -2755 1300 -2735
rect 1320 -2755 1340 -2735
rect 1360 -2755 1380 -2735
rect 1400 -2755 1420 -2735
rect 1440 -2755 1460 -2735
rect 1480 -2755 1500 -2735
rect 1520 -2755 1540 -2735
rect 1560 -2755 1580 -2735
rect 1600 -2755 1620 -2735
rect 1640 -2755 1660 -2735
rect 1680 -2755 1700 -2735
rect 1720 -2755 1740 -2735
rect 1760 -2755 1780 -2735
rect 1800 -2755 1820 -2735
rect 1840 -2755 1860 -2735
rect 1880 -2755 1900 -2735
rect 1920 -2755 1940 -2735
rect 1960 -2755 1980 -2735
rect 2000 -2755 2020 -2735
rect 2040 -2755 2060 -2735
rect 2080 -2755 2100 -2735
rect 2120 -2755 2140 -2735
rect 2160 -2755 2180 -2735
rect 2200 -2755 2220 -2735
rect 2240 -2755 2260 -2735
rect 2280 -2755 2300 -2735
rect 2320 -2755 2340 -2735
rect 2360 -2755 2380 -2735
rect 2400 -2755 2420 -2735
rect 2440 -2755 2460 -2735
rect 2480 -2755 2500 -2735
rect 2520 -2755 2540 -2735
rect 2560 -2755 2590 -2735
<< psubdiff >>
rect 175 2260 2675 2270
rect 175 2240 200 2260
rect 220 2240 240 2260
rect 260 2240 280 2260
rect 300 2240 320 2260
rect 340 2240 360 2260
rect 380 2240 400 2260
rect 420 2240 440 2260
rect 460 2240 480 2260
rect 500 2240 520 2260
rect 540 2240 560 2260
rect 580 2240 600 2260
rect 620 2240 640 2260
rect 660 2240 680 2260
rect 700 2240 720 2260
rect 740 2240 760 2260
rect 780 2240 800 2260
rect 820 2240 840 2260
rect 860 2240 880 2260
rect 900 2240 920 2260
rect 940 2240 960 2260
rect 980 2240 1000 2260
rect 1020 2240 1040 2260
rect 1060 2240 1080 2260
rect 1100 2240 1120 2260
rect 1140 2240 1160 2260
rect 1180 2240 1200 2260
rect 1220 2240 1240 2260
rect 1260 2240 1280 2260
rect 1300 2240 1320 2260
rect 1340 2240 1360 2260
rect 1380 2240 1400 2260
rect 1420 2240 1440 2260
rect 1460 2240 1480 2260
rect 1500 2240 1520 2260
rect 1540 2240 1560 2260
rect 1580 2240 1600 2260
rect 1620 2240 1640 2260
rect 1660 2240 1680 2260
rect 1700 2240 1720 2260
rect 1740 2240 1760 2260
rect 1780 2240 1800 2260
rect 1820 2240 1840 2260
rect 1860 2240 1880 2260
rect 1900 2240 1920 2260
rect 1940 2240 1960 2260
rect 1980 2240 2000 2260
rect 2020 2240 2040 2260
rect 2060 2240 2080 2260
rect 2100 2240 2120 2260
rect 2140 2240 2160 2260
rect 2180 2240 2200 2260
rect 2220 2240 2240 2260
rect 2260 2240 2280 2260
rect 2300 2240 2320 2260
rect 2340 2240 2360 2260
rect 2380 2240 2400 2260
rect 2420 2240 2440 2260
rect 2460 2240 2480 2260
rect 2500 2240 2520 2260
rect 2540 2240 2560 2260
rect 2580 2240 2600 2260
rect 2620 2240 2640 2260
rect 2660 2240 2675 2260
rect 175 2230 2675 2240
rect 175 45 2675 55
rect 175 25 200 45
rect 220 25 240 45
rect 260 25 280 45
rect 300 25 320 45
rect 340 25 360 45
rect 380 25 400 45
rect 420 25 440 45
rect 460 25 480 45
rect 500 25 520 45
rect 540 25 560 45
rect 580 25 600 45
rect 620 25 640 45
rect 660 25 680 45
rect 700 25 720 45
rect 740 25 760 45
rect 780 25 800 45
rect 820 25 840 45
rect 860 25 880 45
rect 900 25 920 45
rect 940 25 960 45
rect 980 25 1000 45
rect 1020 25 1040 45
rect 1060 25 1080 45
rect 1100 25 1120 45
rect 1140 25 1160 45
rect 1180 25 1200 45
rect 1220 25 1240 45
rect 1260 25 1280 45
rect 1300 25 1320 45
rect 1340 25 1360 45
rect 1380 25 1400 45
rect 1420 25 1440 45
rect 1460 25 1480 45
rect 1500 25 1520 45
rect 1540 25 1560 45
rect 1580 25 1600 45
rect 1620 25 1640 45
rect 1660 25 1680 45
rect 1700 25 1720 45
rect 1740 25 1760 45
rect 1780 25 1800 45
rect 1820 25 1840 45
rect 1860 25 1880 45
rect 1900 25 1920 45
rect 1940 25 1960 45
rect 1980 25 2000 45
rect 2020 25 2040 45
rect 2060 25 2080 45
rect 2100 25 2120 45
rect 2140 25 2160 45
rect 2180 25 2200 45
rect 2220 25 2240 45
rect 2260 25 2280 45
rect 2300 25 2320 45
rect 2340 25 2360 45
rect 2380 25 2400 45
rect 2420 25 2440 45
rect 2460 25 2480 45
rect 2500 25 2520 45
rect 2540 25 2560 45
rect 2580 25 2600 45
rect 2620 25 2640 45
rect 2660 25 2675 45
rect 175 15 2675 25
rect 105 -225 2605 -215
rect 105 -245 120 -225
rect 140 -245 160 -225
rect 180 -245 200 -225
rect 220 -245 240 -225
rect 260 -245 280 -225
rect 300 -245 320 -225
rect 340 -245 360 -225
rect 380 -245 400 -225
rect 420 -245 440 -225
rect 460 -245 480 -225
rect 500 -245 520 -225
rect 540 -245 560 -225
rect 580 -245 600 -225
rect 620 -245 640 -225
rect 660 -245 680 -225
rect 700 -245 720 -225
rect 740 -245 760 -225
rect 780 -245 800 -225
rect 820 -245 840 -225
rect 860 -245 880 -225
rect 900 -245 920 -225
rect 940 -245 960 -225
rect 980 -245 1000 -225
rect 1020 -245 1040 -225
rect 1060 -245 1080 -225
rect 1100 -245 1120 -225
rect 1140 -245 1160 -225
rect 1180 -245 1200 -225
rect 1220 -245 1240 -225
rect 1260 -245 1280 -225
rect 1300 -245 1320 -225
rect 1340 -245 1360 -225
rect 1380 -245 1400 -225
rect 1420 -245 1440 -225
rect 1460 -245 1480 -225
rect 1500 -245 1520 -225
rect 1540 -245 1560 -225
rect 1580 -245 1600 -225
rect 1620 -245 1640 -225
rect 1660 -245 1680 -225
rect 1700 -245 1720 -225
rect 1740 -245 1760 -225
rect 1780 -245 1800 -225
rect 1820 -245 1840 -225
rect 1860 -245 1880 -225
rect 1900 -245 1920 -225
rect 1940 -245 1960 -225
rect 1980 -245 2000 -225
rect 2020 -245 2040 -225
rect 2060 -245 2080 -225
rect 2100 -245 2120 -225
rect 2140 -245 2160 -225
rect 2180 -245 2200 -225
rect 2220 -245 2240 -225
rect 2260 -245 2280 -225
rect 2300 -245 2320 -225
rect 2340 -245 2360 -225
rect 2380 -245 2400 -225
rect 2420 -245 2440 -225
rect 2460 -245 2480 -225
rect 2500 -245 2520 -225
rect 2540 -245 2560 -225
rect 2590 -245 2605 -225
rect 105 -255 2605 -245
rect 105 -2775 2605 -2765
rect 105 -2795 120 -2775
rect 140 -2795 160 -2775
rect 180 -2795 200 -2775
rect 220 -2795 240 -2775
rect 260 -2795 280 -2775
rect 300 -2795 320 -2775
rect 340 -2795 360 -2775
rect 380 -2795 400 -2775
rect 420 -2795 440 -2775
rect 460 -2795 480 -2775
rect 500 -2795 520 -2775
rect 540 -2795 560 -2775
rect 580 -2795 600 -2775
rect 620 -2795 640 -2775
rect 660 -2795 680 -2775
rect 700 -2795 720 -2775
rect 740 -2795 760 -2775
rect 780 -2795 800 -2775
rect 820 -2795 840 -2775
rect 860 -2795 880 -2775
rect 900 -2795 920 -2775
rect 940 -2795 960 -2775
rect 980 -2795 1000 -2775
rect 1020 -2795 1040 -2775
rect 1060 -2795 1080 -2775
rect 1100 -2795 1120 -2775
rect 1140 -2795 1160 -2775
rect 1180 -2795 1200 -2775
rect 1220 -2795 1240 -2775
rect 1260 -2795 1280 -2775
rect 1300 -2795 1320 -2775
rect 1340 -2795 1360 -2775
rect 1380 -2795 1400 -2775
rect 1420 -2795 1440 -2775
rect 1460 -2795 1480 -2775
rect 1500 -2795 1520 -2775
rect 1540 -2795 1560 -2775
rect 1580 -2795 1600 -2775
rect 1620 -2795 1640 -2775
rect 1660 -2795 1680 -2775
rect 1700 -2795 1720 -2775
rect 1740 -2795 1760 -2775
rect 1780 -2795 1800 -2775
rect 1820 -2795 1840 -2775
rect 1860 -2795 1880 -2775
rect 1900 -2795 1920 -2775
rect 1940 -2795 1960 -2775
rect 1980 -2795 2000 -2775
rect 2020 -2795 2040 -2775
rect 2060 -2795 2080 -2775
rect 2100 -2795 2120 -2775
rect 2140 -2795 2160 -2775
rect 2180 -2795 2200 -2775
rect 2220 -2795 2240 -2775
rect 2260 -2795 2280 -2775
rect 2300 -2795 2320 -2775
rect 2340 -2795 2360 -2775
rect 2380 -2795 2400 -2775
rect 2420 -2795 2440 -2775
rect 2460 -2795 2480 -2775
rect 2500 -2795 2520 -2775
rect 2540 -2795 2560 -2775
rect 2590 -2795 2605 -2775
rect 105 -2805 2605 -2795
<< nsubdiff >>
rect 1805 -35 1975 -20
rect 1805 -55 1820 -35
rect 1840 -55 1860 -35
rect 1880 -55 1900 -35
rect 1920 -55 1940 -35
rect 1960 -55 1975 -35
rect 1805 -70 1975 -55
<< psubdiffcont >>
rect 200 2240 220 2260
rect 240 2240 260 2260
rect 280 2240 300 2260
rect 320 2240 340 2260
rect 360 2240 380 2260
rect 400 2240 420 2260
rect 440 2240 460 2260
rect 480 2240 500 2260
rect 520 2240 540 2260
rect 560 2240 580 2260
rect 600 2240 620 2260
rect 640 2240 660 2260
rect 680 2240 700 2260
rect 720 2240 740 2260
rect 760 2240 780 2260
rect 800 2240 820 2260
rect 840 2240 860 2260
rect 880 2240 900 2260
rect 920 2240 940 2260
rect 960 2240 980 2260
rect 1000 2240 1020 2260
rect 1040 2240 1060 2260
rect 1080 2240 1100 2260
rect 1120 2240 1140 2260
rect 1160 2240 1180 2260
rect 1200 2240 1220 2260
rect 1240 2240 1260 2260
rect 1280 2240 1300 2260
rect 1320 2240 1340 2260
rect 1360 2240 1380 2260
rect 1400 2240 1420 2260
rect 1440 2240 1460 2260
rect 1480 2240 1500 2260
rect 1520 2240 1540 2260
rect 1560 2240 1580 2260
rect 1600 2240 1620 2260
rect 1640 2240 1660 2260
rect 1680 2240 1700 2260
rect 1720 2240 1740 2260
rect 1760 2240 1780 2260
rect 1800 2240 1820 2260
rect 1840 2240 1860 2260
rect 1880 2240 1900 2260
rect 1920 2240 1940 2260
rect 1960 2240 1980 2260
rect 2000 2240 2020 2260
rect 2040 2240 2060 2260
rect 2080 2240 2100 2260
rect 2120 2240 2140 2260
rect 2160 2240 2180 2260
rect 2200 2240 2220 2260
rect 2240 2240 2260 2260
rect 2280 2240 2300 2260
rect 2320 2240 2340 2260
rect 2360 2240 2380 2260
rect 2400 2240 2420 2260
rect 2440 2240 2460 2260
rect 2480 2240 2500 2260
rect 2520 2240 2540 2260
rect 2560 2240 2580 2260
rect 2600 2240 2620 2260
rect 2640 2240 2660 2260
rect 200 25 220 45
rect 240 25 260 45
rect 280 25 300 45
rect 320 25 340 45
rect 360 25 380 45
rect 400 25 420 45
rect 440 25 460 45
rect 480 25 500 45
rect 520 25 540 45
rect 560 25 580 45
rect 600 25 620 45
rect 640 25 660 45
rect 680 25 700 45
rect 720 25 740 45
rect 760 25 780 45
rect 800 25 820 45
rect 840 25 860 45
rect 880 25 900 45
rect 920 25 940 45
rect 960 25 980 45
rect 1000 25 1020 45
rect 1040 25 1060 45
rect 1080 25 1100 45
rect 1120 25 1140 45
rect 1160 25 1180 45
rect 1200 25 1220 45
rect 1240 25 1260 45
rect 1280 25 1300 45
rect 1320 25 1340 45
rect 1360 25 1380 45
rect 1400 25 1420 45
rect 1440 25 1460 45
rect 1480 25 1500 45
rect 1520 25 1540 45
rect 1560 25 1580 45
rect 1600 25 1620 45
rect 1640 25 1660 45
rect 1680 25 1700 45
rect 1720 25 1740 45
rect 1760 25 1780 45
rect 1800 25 1820 45
rect 1840 25 1860 45
rect 1880 25 1900 45
rect 1920 25 1940 45
rect 1960 25 1980 45
rect 2000 25 2020 45
rect 2040 25 2060 45
rect 2080 25 2100 45
rect 2120 25 2140 45
rect 2160 25 2180 45
rect 2200 25 2220 45
rect 2240 25 2260 45
rect 2280 25 2300 45
rect 2320 25 2340 45
rect 2360 25 2380 45
rect 2400 25 2420 45
rect 2440 25 2460 45
rect 2480 25 2500 45
rect 2520 25 2540 45
rect 2560 25 2580 45
rect 2600 25 2620 45
rect 2640 25 2660 45
rect 120 -245 140 -225
rect 160 -245 180 -225
rect 200 -245 220 -225
rect 240 -245 260 -225
rect 280 -245 300 -225
rect 320 -245 340 -225
rect 360 -245 380 -225
rect 400 -245 420 -225
rect 440 -245 460 -225
rect 480 -245 500 -225
rect 520 -245 540 -225
rect 560 -245 580 -225
rect 600 -245 620 -225
rect 640 -245 660 -225
rect 680 -245 700 -225
rect 720 -245 740 -225
rect 760 -245 780 -225
rect 800 -245 820 -225
rect 840 -245 860 -225
rect 880 -245 900 -225
rect 920 -245 940 -225
rect 960 -245 980 -225
rect 1000 -245 1020 -225
rect 1040 -245 1060 -225
rect 1080 -245 1100 -225
rect 1120 -245 1140 -225
rect 1160 -245 1180 -225
rect 1200 -245 1220 -225
rect 1240 -245 1260 -225
rect 1280 -245 1300 -225
rect 1320 -245 1340 -225
rect 1360 -245 1380 -225
rect 1400 -245 1420 -225
rect 1440 -245 1460 -225
rect 1480 -245 1500 -225
rect 1520 -245 1540 -225
rect 1560 -245 1580 -225
rect 1600 -245 1620 -225
rect 1640 -245 1660 -225
rect 1680 -245 1700 -225
rect 1720 -245 1740 -225
rect 1760 -245 1780 -225
rect 1800 -245 1820 -225
rect 1840 -245 1860 -225
rect 1880 -245 1900 -225
rect 1920 -245 1940 -225
rect 1960 -245 1980 -225
rect 2000 -245 2020 -225
rect 2040 -245 2060 -225
rect 2080 -245 2100 -225
rect 2120 -245 2140 -225
rect 2160 -245 2180 -225
rect 2200 -245 2220 -225
rect 2240 -245 2260 -225
rect 2280 -245 2300 -225
rect 2320 -245 2340 -225
rect 2360 -245 2380 -225
rect 2400 -245 2420 -225
rect 2440 -245 2460 -225
rect 2480 -245 2500 -225
rect 2520 -245 2540 -225
rect 2560 -245 2590 -225
rect 120 -2795 140 -2775
rect 160 -2795 180 -2775
rect 200 -2795 220 -2775
rect 240 -2795 260 -2775
rect 280 -2795 300 -2775
rect 320 -2795 340 -2775
rect 360 -2795 380 -2775
rect 400 -2795 420 -2775
rect 440 -2795 460 -2775
rect 480 -2795 500 -2775
rect 520 -2795 540 -2775
rect 560 -2795 580 -2775
rect 600 -2795 620 -2775
rect 640 -2795 660 -2775
rect 680 -2795 700 -2775
rect 720 -2795 740 -2775
rect 760 -2795 780 -2775
rect 800 -2795 820 -2775
rect 840 -2795 860 -2775
rect 880 -2795 900 -2775
rect 920 -2795 940 -2775
rect 960 -2795 980 -2775
rect 1000 -2795 1020 -2775
rect 1040 -2795 1060 -2775
rect 1080 -2795 1100 -2775
rect 1120 -2795 1140 -2775
rect 1160 -2795 1180 -2775
rect 1200 -2795 1220 -2775
rect 1240 -2795 1260 -2775
rect 1280 -2795 1300 -2775
rect 1320 -2795 1340 -2775
rect 1360 -2795 1380 -2775
rect 1400 -2795 1420 -2775
rect 1440 -2795 1460 -2775
rect 1480 -2795 1500 -2775
rect 1520 -2795 1540 -2775
rect 1560 -2795 1580 -2775
rect 1600 -2795 1620 -2775
rect 1640 -2795 1660 -2775
rect 1680 -2795 1700 -2775
rect 1720 -2795 1740 -2775
rect 1760 -2795 1780 -2775
rect 1800 -2795 1820 -2775
rect 1840 -2795 1860 -2775
rect 1880 -2795 1900 -2775
rect 1920 -2795 1940 -2775
rect 1960 -2795 1980 -2775
rect 2000 -2795 2020 -2775
rect 2040 -2795 2060 -2775
rect 2080 -2795 2100 -2775
rect 2120 -2795 2140 -2775
rect 2160 -2795 2180 -2775
rect 2200 -2795 2220 -2775
rect 2240 -2795 2260 -2775
rect 2280 -2795 2300 -2775
rect 2320 -2795 2340 -2775
rect 2360 -2795 2380 -2775
rect 2400 -2795 2420 -2775
rect 2440 -2795 2460 -2775
rect 2480 -2795 2500 -2775
rect 2520 -2795 2540 -2775
rect 2560 -2795 2590 -2775
<< nsubdiffcont >>
rect 1820 -55 1840 -35
rect 1860 -55 1880 -35
rect 1900 -55 1920 -35
rect 1940 -55 1960 -35
<< poly >>
rect 0 2182 165 2185
rect 0 2175 175 2182
rect 0 2155 10 2175
rect 30 2155 50 2175
rect 70 2155 90 2175
rect 110 2155 130 2175
rect 155 2155 175 2175
rect 0 2150 175 2155
rect 2675 2150 2690 2182
rect 0 2145 165 2150
rect 0 2100 165 2105
rect 0 2095 175 2100
rect 0 2075 10 2095
rect 30 2075 50 2095
rect 70 2075 90 2095
rect 110 2075 130 2095
rect 155 2075 175 2095
rect 0 2068 175 2075
rect 2675 2068 2690 2100
rect 0 2065 165 2068
rect 0 2018 165 2020
rect 0 2010 175 2018
rect 0 1990 10 2010
rect 30 1990 50 2010
rect 70 1990 90 2010
rect 110 1990 130 2010
rect 155 1990 175 2010
rect 0 1986 175 1990
rect 2675 1986 2690 2018
rect 0 1980 165 1986
rect 0 1936 165 1940
rect 0 1930 175 1936
rect 0 1910 10 1930
rect 30 1910 50 1930
rect 70 1910 90 1930
rect 110 1910 130 1930
rect 155 1910 175 1930
rect 0 1904 175 1910
rect 2675 1904 2690 1936
rect 0 1900 165 1904
rect 0 1854 165 1860
rect 0 1850 175 1854
rect 0 1830 10 1850
rect 30 1830 50 1850
rect 70 1830 90 1850
rect 110 1830 130 1850
rect 155 1830 175 1850
rect 0 1822 175 1830
rect 2675 1822 2690 1854
rect 0 1820 165 1822
rect 0 1772 165 1775
rect 0 1765 175 1772
rect 0 1745 10 1765
rect 30 1745 50 1765
rect 70 1745 90 1765
rect 110 1745 130 1765
rect 155 1745 175 1765
rect 0 1740 175 1745
rect 2675 1740 2690 1772
rect 0 1735 165 1740
rect 0 1690 165 1695
rect 0 1685 175 1690
rect 0 1665 10 1685
rect 30 1665 50 1685
rect 70 1665 90 1685
rect 110 1665 130 1685
rect 155 1665 175 1685
rect 0 1658 175 1665
rect 2675 1658 2690 1690
rect 0 1655 165 1658
rect 0 1608 165 1610
rect 0 1600 175 1608
rect 0 1580 10 1600
rect 30 1580 50 1600
rect 70 1580 90 1600
rect 110 1580 130 1600
rect 155 1580 175 1600
rect 0 1576 175 1580
rect 2675 1576 2690 1608
rect 0 1570 165 1576
rect 0 1526 165 1530
rect 0 1520 175 1526
rect 0 1500 10 1520
rect 30 1500 50 1520
rect 70 1500 90 1520
rect 110 1500 130 1520
rect 155 1500 175 1520
rect 0 1494 175 1500
rect 2675 1494 2690 1526
rect 0 1490 165 1494
rect 0 1444 165 1450
rect 0 1440 175 1444
rect 0 1420 10 1440
rect 30 1420 50 1440
rect 70 1420 90 1440
rect 110 1420 130 1440
rect 155 1420 175 1440
rect 0 1412 175 1420
rect 2675 1412 2690 1444
rect 0 1410 165 1412
rect 0 1362 165 1365
rect 0 1355 175 1362
rect 0 1335 10 1355
rect 30 1335 50 1355
rect 70 1335 90 1355
rect 110 1335 130 1355
rect 155 1335 175 1355
rect 0 1330 175 1335
rect 2675 1330 2690 1362
rect 0 1325 165 1330
rect 0 1280 165 1285
rect 0 1275 175 1280
rect 0 1255 10 1275
rect 30 1255 50 1275
rect 70 1255 90 1275
rect 110 1255 130 1275
rect 155 1255 175 1275
rect 0 1248 175 1255
rect 2675 1248 2690 1280
rect 0 1245 165 1248
rect 0 1198 165 1200
rect 0 1190 175 1198
rect 0 1170 10 1190
rect 30 1170 50 1190
rect 70 1170 90 1190
rect 110 1170 130 1190
rect 155 1170 175 1190
rect 0 1166 175 1170
rect 2675 1166 2690 1198
rect 0 1160 165 1166
rect 0 1116 165 1120
rect 0 1110 175 1116
rect 0 1090 10 1110
rect 30 1090 50 1110
rect 70 1090 90 1110
rect 110 1090 130 1110
rect 155 1090 175 1110
rect 0 1084 175 1090
rect 2675 1084 2690 1116
rect 0 1080 165 1084
rect 0 1034 165 1040
rect 0 1030 175 1034
rect 0 1010 10 1030
rect 30 1010 50 1030
rect 70 1010 90 1030
rect 110 1010 130 1030
rect 155 1010 175 1030
rect 0 1002 175 1010
rect 2675 1002 2690 1034
rect 0 1000 165 1002
rect 0 952 165 955
rect 0 945 175 952
rect 0 925 10 945
rect 30 925 50 945
rect 70 925 90 945
rect 110 925 130 945
rect 155 925 175 945
rect 0 920 175 925
rect 2675 920 2690 952
rect 0 915 165 920
rect 0 870 165 875
rect 0 865 175 870
rect 0 845 10 865
rect 30 845 50 865
rect 70 845 90 865
rect 110 845 130 865
rect 155 845 175 865
rect 0 838 175 845
rect 2675 838 2690 870
rect 0 835 165 838
rect 0 788 165 790
rect 0 780 175 788
rect 0 760 10 780
rect 30 760 50 780
rect 70 760 90 780
rect 110 760 130 780
rect 155 760 175 780
rect 0 756 175 760
rect 2675 756 2690 788
rect 0 750 165 756
rect 0 706 165 710
rect 0 700 175 706
rect 0 680 10 700
rect 30 680 50 700
rect 70 680 90 700
rect 110 680 130 700
rect 155 680 175 700
rect 0 674 175 680
rect 2675 674 2690 706
rect 0 670 165 674
rect 0 624 165 630
rect 0 620 175 624
rect 0 600 10 620
rect 30 600 50 620
rect 70 600 90 620
rect 110 600 130 620
rect 155 600 175 620
rect 0 592 175 600
rect 2675 592 2690 624
rect 0 590 165 592
rect 0 542 165 545
rect 0 535 175 542
rect 0 515 10 535
rect 30 515 50 535
rect 70 515 90 535
rect 110 515 130 535
rect 155 515 175 535
rect 0 510 175 515
rect 2675 510 2690 542
rect 0 505 165 510
rect 0 460 165 465
rect 0 455 175 460
rect 0 435 10 455
rect 30 435 50 455
rect 70 435 90 455
rect 110 435 130 455
rect 155 435 175 455
rect 0 428 175 435
rect 2675 428 2690 460
rect 0 425 165 428
rect 0 378 165 385
rect 0 375 175 378
rect 0 355 10 375
rect 30 355 50 375
rect 70 355 90 375
rect 110 355 130 375
rect 155 355 175 375
rect 0 346 175 355
rect 2675 346 2690 378
rect 0 345 165 346
rect 0 296 165 300
rect 0 290 175 296
rect 0 270 10 290
rect 30 270 50 290
rect 70 270 90 290
rect 110 270 130 290
rect 155 270 175 290
rect 0 264 175 270
rect 2675 264 2690 296
rect 0 260 165 264
rect 0 214 165 220
rect 0 210 175 214
rect 0 190 10 210
rect 30 190 50 210
rect 70 190 90 210
rect 110 190 130 210
rect 155 190 175 210
rect 0 182 175 190
rect 2675 182 2690 214
rect 0 180 165 182
rect 0 132 165 140
rect 0 130 175 132
rect 0 110 10 130
rect 30 110 50 130
rect 70 110 90 130
rect 110 110 130 130
rect 155 110 175 130
rect 0 100 175 110
rect 2675 100 2690 132
rect -70 -310 105 -300
rect -70 -335 -60 -310
rect -40 -335 -20 -310
rect 0 -335 20 -310
rect 40 -335 60 -310
rect 85 -335 105 -310
rect -70 -345 105 -335
rect 2605 -345 2620 -300
rect -70 -405 105 -395
rect -70 -430 -60 -405
rect -40 -430 -20 -405
rect 0 -430 20 -405
rect 40 -430 60 -405
rect 85 -430 105 -405
rect -70 -440 105 -430
rect 2605 -440 2620 -395
rect -70 -500 105 -490
rect -70 -525 -60 -500
rect -40 -525 -20 -500
rect 0 -525 20 -500
rect 40 -525 60 -500
rect 85 -525 105 -500
rect -70 -535 105 -525
rect 2605 -535 2620 -490
rect -70 -595 105 -585
rect -70 -620 -60 -595
rect -40 -620 -20 -595
rect 0 -620 20 -595
rect 40 -620 60 -595
rect 85 -620 105 -595
rect -70 -630 105 -620
rect 2605 -630 2620 -585
rect -70 -690 105 -680
rect -70 -715 -60 -690
rect -40 -715 -20 -690
rect 0 -715 20 -690
rect 40 -715 60 -690
rect 85 -715 105 -690
rect -70 -725 105 -715
rect 2605 -725 2620 -680
rect -70 -785 105 -775
rect -70 -810 -60 -785
rect -40 -810 -20 -785
rect 0 -810 20 -785
rect 40 -810 60 -785
rect 85 -810 105 -785
rect -70 -820 105 -810
rect 2605 -820 2620 -775
rect -70 -880 105 -870
rect -70 -905 -60 -880
rect -40 -905 -20 -880
rect 0 -905 20 -880
rect 40 -905 60 -880
rect 85 -905 105 -880
rect -70 -915 105 -905
rect 2605 -915 2620 -870
rect -70 -975 105 -965
rect -70 -1000 -60 -975
rect -40 -1000 -20 -975
rect 0 -1000 20 -975
rect 40 -1000 60 -975
rect 85 -1000 105 -975
rect -70 -1010 105 -1000
rect 2605 -1010 2620 -965
rect -70 -1070 105 -1060
rect -70 -1095 -60 -1070
rect -40 -1095 -20 -1070
rect 0 -1095 20 -1070
rect 40 -1095 60 -1070
rect 85 -1095 105 -1070
rect -70 -1105 105 -1095
rect 2605 -1105 2620 -1060
rect -70 -1165 105 -1155
rect -70 -1190 -60 -1165
rect -40 -1190 -20 -1165
rect 0 -1190 20 -1165
rect 40 -1190 60 -1165
rect 85 -1190 105 -1165
rect -70 -1200 105 -1190
rect 2605 -1200 2620 -1155
rect -70 -1260 105 -1250
rect -70 -1285 -60 -1260
rect -40 -1285 -20 -1260
rect 0 -1285 20 -1260
rect 40 -1285 60 -1260
rect 85 -1285 105 -1260
rect -70 -1295 105 -1285
rect 2605 -1295 2620 -1250
rect -70 -1355 105 -1345
rect -70 -1380 -60 -1355
rect -40 -1380 -20 -1355
rect 0 -1380 20 -1355
rect 40 -1380 60 -1355
rect 85 -1380 105 -1355
rect -70 -1390 105 -1380
rect 2605 -1390 2620 -1345
rect -70 -1450 105 -1440
rect -70 -1475 -60 -1450
rect -40 -1475 -20 -1450
rect 0 -1475 20 -1450
rect 40 -1475 60 -1450
rect 85 -1475 105 -1450
rect -70 -1485 105 -1475
rect 2605 -1485 2620 -1440
rect -70 -1545 105 -1535
rect -70 -1570 -60 -1545
rect -40 -1570 -20 -1545
rect 0 -1570 20 -1545
rect 40 -1570 60 -1545
rect 85 -1570 105 -1545
rect -70 -1580 105 -1570
rect 2605 -1580 2620 -1535
rect -70 -1640 105 -1630
rect -70 -1665 -60 -1640
rect -40 -1665 -20 -1640
rect 0 -1665 20 -1640
rect 40 -1665 60 -1640
rect 85 -1665 105 -1640
rect -70 -1675 105 -1665
rect 2605 -1675 2620 -1630
rect -70 -1735 105 -1725
rect -70 -1760 -60 -1735
rect -40 -1760 -20 -1735
rect 0 -1760 20 -1735
rect 40 -1760 60 -1735
rect 85 -1760 105 -1735
rect -70 -1770 105 -1760
rect 2605 -1770 2620 -1725
rect -70 -1830 105 -1820
rect -70 -1855 -60 -1830
rect -40 -1855 -20 -1830
rect 0 -1855 20 -1830
rect 40 -1855 60 -1830
rect 85 -1855 105 -1830
rect -70 -1865 105 -1855
rect 2605 -1865 2620 -1820
rect -70 -1925 105 -1915
rect -70 -1950 -60 -1925
rect -40 -1950 -20 -1925
rect 0 -1950 20 -1925
rect 40 -1950 60 -1925
rect 85 -1950 105 -1925
rect -70 -1960 105 -1950
rect 2605 -1960 2620 -1915
rect -70 -2020 105 -2010
rect -70 -2045 -60 -2020
rect -40 -2045 -20 -2020
rect 0 -2045 20 -2020
rect 40 -2045 60 -2020
rect 85 -2045 105 -2020
rect -70 -2055 105 -2045
rect 2605 -2055 2620 -2010
rect -70 -2115 105 -2105
rect -70 -2140 -60 -2115
rect -40 -2140 -20 -2115
rect 0 -2140 20 -2115
rect 40 -2140 60 -2115
rect 85 -2140 105 -2115
rect -70 -2150 105 -2140
rect 2605 -2150 2620 -2105
rect -70 -2210 105 -2200
rect -70 -2235 -60 -2210
rect -40 -2235 -20 -2210
rect 0 -2235 20 -2210
rect 40 -2235 60 -2210
rect 85 -2235 105 -2210
rect -70 -2245 105 -2235
rect 2605 -2245 2620 -2200
rect -70 -2305 105 -2295
rect -70 -2330 -60 -2305
rect -40 -2330 -20 -2305
rect 0 -2330 20 -2305
rect 40 -2330 60 -2305
rect 85 -2330 105 -2305
rect -70 -2340 105 -2330
rect 2605 -2340 2620 -2295
rect -70 -2400 105 -2390
rect -70 -2425 -60 -2400
rect -40 -2425 -20 -2400
rect 0 -2425 20 -2400
rect 40 -2425 60 -2400
rect 85 -2425 105 -2400
rect -70 -2435 105 -2425
rect 2605 -2435 2620 -2390
rect -70 -2495 105 -2485
rect -70 -2520 -60 -2495
rect -40 -2520 -20 -2495
rect 0 -2520 20 -2495
rect 40 -2520 60 -2495
rect 85 -2520 105 -2495
rect -70 -2530 105 -2520
rect 2605 -2530 2620 -2485
rect -70 -2590 105 -2580
rect -70 -2615 -60 -2590
rect -40 -2615 -20 -2590
rect 0 -2615 20 -2590
rect 40 -2615 60 -2590
rect 85 -2615 105 -2590
rect -70 -2625 105 -2615
rect 2605 -2625 2620 -2580
rect -70 -2685 105 -2675
rect -70 -2710 -60 -2685
rect -40 -2710 -20 -2685
rect 0 -2710 20 -2685
rect 40 -2710 60 -2685
rect 85 -2710 105 -2685
rect -70 -2720 105 -2710
rect 2605 -2720 2620 -2675
<< polycont >>
rect 10 2155 30 2175
rect 50 2155 70 2175
rect 90 2155 110 2175
rect 130 2155 155 2175
rect 10 2075 30 2095
rect 50 2075 70 2095
rect 90 2075 110 2095
rect 130 2075 155 2095
rect 10 1990 30 2010
rect 50 1990 70 2010
rect 90 1990 110 2010
rect 130 1990 155 2010
rect 10 1910 30 1930
rect 50 1910 70 1930
rect 90 1910 110 1930
rect 130 1910 155 1930
rect 10 1830 30 1850
rect 50 1830 70 1850
rect 90 1830 110 1850
rect 130 1830 155 1850
rect 10 1745 30 1765
rect 50 1745 70 1765
rect 90 1745 110 1765
rect 130 1745 155 1765
rect 10 1665 30 1685
rect 50 1665 70 1685
rect 90 1665 110 1685
rect 130 1665 155 1685
rect 10 1580 30 1600
rect 50 1580 70 1600
rect 90 1580 110 1600
rect 130 1580 155 1600
rect 10 1500 30 1520
rect 50 1500 70 1520
rect 90 1500 110 1520
rect 130 1500 155 1520
rect 10 1420 30 1440
rect 50 1420 70 1440
rect 90 1420 110 1440
rect 130 1420 155 1440
rect 10 1335 30 1355
rect 50 1335 70 1355
rect 90 1335 110 1355
rect 130 1335 155 1355
rect 10 1255 30 1275
rect 50 1255 70 1275
rect 90 1255 110 1275
rect 130 1255 155 1275
rect 10 1170 30 1190
rect 50 1170 70 1190
rect 90 1170 110 1190
rect 130 1170 155 1190
rect 10 1090 30 1110
rect 50 1090 70 1110
rect 90 1090 110 1110
rect 130 1090 155 1110
rect 10 1010 30 1030
rect 50 1010 70 1030
rect 90 1010 110 1030
rect 130 1010 155 1030
rect 10 925 30 945
rect 50 925 70 945
rect 90 925 110 945
rect 130 925 155 945
rect 10 845 30 865
rect 50 845 70 865
rect 90 845 110 865
rect 130 845 155 865
rect 10 760 30 780
rect 50 760 70 780
rect 90 760 110 780
rect 130 760 155 780
rect 10 680 30 700
rect 50 680 70 700
rect 90 680 110 700
rect 130 680 155 700
rect 10 600 30 620
rect 50 600 70 620
rect 90 600 110 620
rect 130 600 155 620
rect 10 515 30 535
rect 50 515 70 535
rect 90 515 110 535
rect 130 515 155 535
rect 10 435 30 455
rect 50 435 70 455
rect 90 435 110 455
rect 130 435 155 455
rect 10 355 30 375
rect 50 355 70 375
rect 90 355 110 375
rect 130 355 155 375
rect 10 270 30 290
rect 50 270 70 290
rect 90 270 110 290
rect 130 270 155 290
rect 10 190 30 210
rect 50 190 70 210
rect 90 190 110 210
rect 130 190 155 210
rect 10 110 30 130
rect 50 110 70 130
rect 90 110 110 130
rect 130 110 155 130
rect -60 -335 -40 -310
rect -20 -335 0 -310
rect 20 -335 40 -310
rect 60 -335 85 -310
rect -60 -430 -40 -405
rect -20 -430 0 -405
rect 20 -430 40 -405
rect 60 -430 85 -405
rect -60 -525 -40 -500
rect -20 -525 0 -500
rect 20 -525 40 -500
rect 60 -525 85 -500
rect -60 -620 -40 -595
rect -20 -620 0 -595
rect 20 -620 40 -595
rect 60 -620 85 -595
rect -60 -715 -40 -690
rect -20 -715 0 -690
rect 20 -715 40 -690
rect 60 -715 85 -690
rect -60 -810 -40 -785
rect -20 -810 0 -785
rect 20 -810 40 -785
rect 60 -810 85 -785
rect -60 -905 -40 -880
rect -20 -905 0 -880
rect 20 -905 40 -880
rect 60 -905 85 -880
rect -60 -1000 -40 -975
rect -20 -1000 0 -975
rect 20 -1000 40 -975
rect 60 -1000 85 -975
rect -60 -1095 -40 -1070
rect -20 -1095 0 -1070
rect 20 -1095 40 -1070
rect 60 -1095 85 -1070
rect -60 -1190 -40 -1165
rect -20 -1190 0 -1165
rect 20 -1190 40 -1165
rect 60 -1190 85 -1165
rect -60 -1285 -40 -1260
rect -20 -1285 0 -1260
rect 20 -1285 40 -1260
rect 60 -1285 85 -1260
rect -60 -1380 -40 -1355
rect -20 -1380 0 -1355
rect 20 -1380 40 -1355
rect 60 -1380 85 -1355
rect -60 -1475 -40 -1450
rect -20 -1475 0 -1450
rect 20 -1475 40 -1450
rect 60 -1475 85 -1450
rect -60 -1570 -40 -1545
rect -20 -1570 0 -1545
rect 20 -1570 40 -1545
rect 60 -1570 85 -1545
rect -60 -1665 -40 -1640
rect -20 -1665 0 -1640
rect 20 -1665 40 -1640
rect 60 -1665 85 -1640
rect -60 -1760 -40 -1735
rect -20 -1760 0 -1735
rect 20 -1760 40 -1735
rect 60 -1760 85 -1735
rect -60 -1855 -40 -1830
rect -20 -1855 0 -1830
rect 20 -1855 40 -1830
rect 60 -1855 85 -1830
rect -60 -1950 -40 -1925
rect -20 -1950 0 -1925
rect 20 -1950 40 -1925
rect 60 -1950 85 -1925
rect -60 -2045 -40 -2020
rect -20 -2045 0 -2020
rect 20 -2045 40 -2020
rect 60 -2045 85 -2020
rect -60 -2140 -40 -2115
rect -20 -2140 0 -2115
rect 20 -2140 40 -2115
rect 60 -2140 85 -2115
rect -60 -2235 -40 -2210
rect -20 -2235 0 -2210
rect 20 -2235 40 -2210
rect 60 -2235 85 -2210
rect -60 -2330 -40 -2305
rect -20 -2330 0 -2305
rect 20 -2330 40 -2305
rect 60 -2330 85 -2305
rect -60 -2425 -40 -2400
rect -20 -2425 0 -2400
rect 20 -2425 40 -2400
rect 60 -2425 85 -2400
rect -60 -2520 -40 -2495
rect -20 -2520 0 -2495
rect 20 -2520 40 -2495
rect 60 -2520 85 -2495
rect -60 -2615 -40 -2590
rect -20 -2615 0 -2590
rect 20 -2615 40 -2590
rect 60 -2615 85 -2590
rect -60 -2710 -40 -2685
rect -20 -2710 0 -2685
rect 20 -2710 40 -2685
rect 60 -2710 85 -2685
<< locali >>
rect 175 2260 2675 2270
rect 175 2240 200 2260
rect 220 2240 240 2260
rect 260 2240 280 2260
rect 300 2240 320 2260
rect 340 2240 360 2260
rect 380 2240 400 2260
rect 420 2240 440 2260
rect 460 2240 480 2260
rect 500 2240 520 2260
rect 540 2240 560 2260
rect 580 2240 600 2260
rect 620 2240 640 2260
rect 660 2240 680 2260
rect 700 2240 720 2260
rect 740 2240 760 2260
rect 780 2240 800 2260
rect 820 2240 840 2260
rect 860 2240 880 2260
rect 900 2240 920 2260
rect 940 2240 960 2260
rect 980 2240 1000 2260
rect 1020 2240 1040 2260
rect 1060 2240 1080 2260
rect 1100 2240 1120 2260
rect 1140 2240 1160 2260
rect 1180 2240 1200 2260
rect 1220 2240 1240 2260
rect 1260 2240 1280 2260
rect 1300 2240 1320 2260
rect 1340 2240 1360 2260
rect 1380 2240 1400 2260
rect 1420 2240 1440 2260
rect 1460 2240 1480 2260
rect 1500 2240 1520 2260
rect 1540 2240 1560 2260
rect 1580 2240 1600 2260
rect 1620 2240 1640 2260
rect 1660 2240 1680 2260
rect 1700 2240 1720 2260
rect 1740 2240 1760 2260
rect 1780 2240 1800 2260
rect 1820 2240 1840 2260
rect 1860 2240 1880 2260
rect 1900 2240 1920 2260
rect 1940 2240 1960 2260
rect 1980 2240 2000 2260
rect 2020 2240 2040 2260
rect 2060 2240 2080 2260
rect 2100 2240 2120 2260
rect 2140 2240 2160 2260
rect 2180 2240 2200 2260
rect 2220 2240 2240 2260
rect 2260 2240 2280 2260
rect 2300 2240 2320 2260
rect 2340 2240 2360 2260
rect 2380 2240 2400 2260
rect 2420 2240 2440 2260
rect 2460 2240 2480 2260
rect 2500 2240 2520 2260
rect 2540 2240 2560 2260
rect 2580 2240 2600 2260
rect 2620 2240 2640 2260
rect 2660 2240 2675 2260
rect 175 2217 2675 2240
rect 175 2197 200 2217
rect 220 2197 240 2217
rect 260 2197 280 2217
rect 300 2197 320 2217
rect 340 2197 360 2217
rect 380 2197 400 2217
rect 420 2197 440 2217
rect 460 2197 480 2217
rect 500 2197 520 2217
rect 540 2197 560 2217
rect 580 2197 600 2217
rect 620 2197 640 2217
rect 660 2197 680 2217
rect 700 2197 720 2217
rect 740 2197 760 2217
rect 780 2197 800 2217
rect 820 2197 840 2217
rect 860 2197 880 2217
rect 900 2197 920 2217
rect 940 2197 960 2217
rect 980 2197 1000 2217
rect 1020 2197 1040 2217
rect 1060 2197 1080 2217
rect 1100 2197 1120 2217
rect 1140 2197 1160 2217
rect 1180 2197 1200 2217
rect 1220 2197 1240 2217
rect 1260 2197 1280 2217
rect 1300 2197 1320 2217
rect 1340 2197 1360 2217
rect 1380 2197 1400 2217
rect 1420 2197 1440 2217
rect 1460 2197 1480 2217
rect 1500 2197 1520 2217
rect 1540 2197 1560 2217
rect 1580 2197 1600 2217
rect 1620 2197 1640 2217
rect 1660 2197 1680 2217
rect 1700 2197 1720 2217
rect 1740 2197 1760 2217
rect 1780 2197 1800 2217
rect 1820 2197 1840 2217
rect 1860 2197 1880 2217
rect 1900 2197 1920 2217
rect 1940 2197 1960 2217
rect 1980 2197 2000 2217
rect 2020 2197 2040 2217
rect 2060 2197 2080 2217
rect 2100 2197 2120 2217
rect 2140 2197 2160 2217
rect 2180 2197 2200 2217
rect 2220 2197 2240 2217
rect 2260 2197 2280 2217
rect 2300 2197 2320 2217
rect 2340 2197 2360 2217
rect 2380 2197 2400 2217
rect 2420 2197 2440 2217
rect 2460 2197 2480 2217
rect 2500 2197 2520 2217
rect 2540 2197 2560 2217
rect 2580 2197 2600 2217
rect 2620 2197 2640 2217
rect 2660 2197 2675 2217
rect 175 2187 2675 2197
rect 0 2175 155 2185
rect 0 2155 10 2175
rect 30 2155 50 2175
rect 70 2155 90 2175
rect 110 2155 130 2175
rect 0 2145 155 2155
rect 175 2135 2675 2145
rect 175 2115 200 2135
rect 220 2115 240 2135
rect 260 2115 280 2135
rect 300 2115 320 2135
rect 340 2115 360 2135
rect 380 2115 400 2135
rect 420 2115 440 2135
rect 460 2115 480 2135
rect 500 2115 520 2135
rect 540 2115 560 2135
rect 580 2115 600 2135
rect 620 2115 640 2135
rect 660 2115 680 2135
rect 700 2115 720 2135
rect 740 2115 760 2135
rect 780 2115 800 2135
rect 820 2115 840 2135
rect 860 2115 880 2135
rect 900 2115 920 2135
rect 940 2115 960 2135
rect 980 2115 1000 2135
rect 1020 2115 1040 2135
rect 1060 2115 1080 2135
rect 1100 2115 1120 2135
rect 1140 2115 1160 2135
rect 1180 2115 1200 2135
rect 1220 2115 1240 2135
rect 1260 2115 1280 2135
rect 1300 2115 1320 2135
rect 1340 2115 1360 2135
rect 1380 2115 1400 2135
rect 1420 2115 1440 2135
rect 1460 2115 1480 2135
rect 1500 2115 1520 2135
rect 1540 2115 1560 2135
rect 1580 2115 1600 2135
rect 1620 2115 1640 2135
rect 1660 2115 1680 2135
rect 1700 2115 1720 2135
rect 1740 2115 1760 2135
rect 1780 2115 1800 2135
rect 1820 2115 1840 2135
rect 1860 2115 1880 2135
rect 1900 2115 1920 2135
rect 1940 2115 1960 2135
rect 1980 2115 2000 2135
rect 2020 2115 2040 2135
rect 2060 2115 2080 2135
rect 2100 2115 2120 2135
rect 2140 2115 2160 2135
rect 2180 2115 2200 2135
rect 2220 2115 2240 2135
rect 2260 2115 2280 2135
rect 2300 2115 2320 2135
rect 2340 2115 2360 2135
rect 2380 2115 2400 2135
rect 2420 2115 2440 2135
rect 2460 2115 2480 2135
rect 2500 2115 2520 2135
rect 2540 2115 2560 2135
rect 2580 2115 2600 2135
rect 2620 2115 2640 2135
rect 2660 2115 2675 2135
rect 175 2105 2675 2115
rect 0 2095 155 2105
rect 0 2075 10 2095
rect 30 2075 50 2095
rect 70 2075 90 2095
rect 110 2075 130 2095
rect 0 2065 155 2075
rect 175 2053 2675 2063
rect 175 2033 200 2053
rect 220 2033 240 2053
rect 260 2033 280 2053
rect 300 2033 320 2053
rect 340 2033 360 2053
rect 380 2033 400 2053
rect 420 2033 440 2053
rect 460 2033 480 2053
rect 500 2033 520 2053
rect 540 2033 560 2053
rect 580 2033 600 2053
rect 620 2033 640 2053
rect 660 2033 680 2053
rect 700 2033 720 2053
rect 740 2033 760 2053
rect 780 2033 800 2053
rect 820 2033 840 2053
rect 860 2033 880 2053
rect 900 2033 920 2053
rect 940 2033 960 2053
rect 980 2033 1000 2053
rect 1020 2033 1040 2053
rect 1060 2033 1080 2053
rect 1100 2033 1120 2053
rect 1140 2033 1160 2053
rect 1180 2033 1200 2053
rect 1220 2033 1240 2053
rect 1260 2033 1280 2053
rect 1300 2033 1320 2053
rect 1340 2033 1360 2053
rect 1380 2033 1400 2053
rect 1420 2033 1440 2053
rect 1460 2033 1480 2053
rect 1500 2033 1520 2053
rect 1540 2033 1560 2053
rect 1580 2033 1600 2053
rect 1620 2033 1640 2053
rect 1660 2033 1680 2053
rect 1700 2033 1720 2053
rect 1740 2033 1760 2053
rect 1780 2033 1800 2053
rect 1820 2033 1840 2053
rect 1860 2033 1880 2053
rect 1900 2033 1920 2053
rect 1940 2033 1960 2053
rect 1980 2033 2000 2053
rect 2020 2033 2040 2053
rect 2060 2033 2080 2053
rect 2100 2033 2120 2053
rect 2140 2033 2160 2053
rect 2180 2033 2200 2053
rect 2220 2033 2240 2053
rect 2260 2033 2280 2053
rect 2300 2033 2320 2053
rect 2340 2033 2360 2053
rect 2380 2033 2400 2053
rect 2420 2033 2440 2053
rect 2460 2033 2480 2053
rect 2500 2033 2520 2053
rect 2540 2033 2560 2053
rect 2580 2033 2600 2053
rect 2620 2033 2640 2053
rect 2660 2033 2675 2053
rect 175 2023 2675 2033
rect 0 2010 155 2020
rect 0 1990 10 2010
rect 30 1990 50 2010
rect 70 1990 90 2010
rect 110 1990 130 2010
rect 0 1980 155 1990
rect 175 1971 2675 1981
rect 175 1951 200 1971
rect 220 1951 240 1971
rect 260 1951 280 1971
rect 300 1951 320 1971
rect 340 1951 360 1971
rect 380 1951 400 1971
rect 420 1951 440 1971
rect 460 1951 480 1971
rect 500 1951 520 1971
rect 540 1951 560 1971
rect 580 1951 600 1971
rect 620 1951 640 1971
rect 660 1951 680 1971
rect 700 1951 720 1971
rect 740 1951 760 1971
rect 780 1951 800 1971
rect 820 1951 840 1971
rect 860 1951 880 1971
rect 900 1951 920 1971
rect 940 1951 960 1971
rect 980 1951 1000 1971
rect 1020 1951 1040 1971
rect 1060 1951 1080 1971
rect 1100 1951 1120 1971
rect 1140 1951 1160 1971
rect 1180 1951 1200 1971
rect 1220 1951 1240 1971
rect 1260 1951 1280 1971
rect 1300 1951 1320 1971
rect 1340 1951 1360 1971
rect 1380 1951 1400 1971
rect 1420 1951 1440 1971
rect 1460 1951 1480 1971
rect 1500 1951 1520 1971
rect 1540 1951 1560 1971
rect 1580 1951 1600 1971
rect 1620 1951 1640 1971
rect 1660 1951 1680 1971
rect 1700 1951 1720 1971
rect 1740 1951 1760 1971
rect 1780 1951 1800 1971
rect 1820 1951 1840 1971
rect 1860 1951 1880 1971
rect 1900 1951 1920 1971
rect 1940 1951 1960 1971
rect 1980 1951 2000 1971
rect 2020 1951 2040 1971
rect 2060 1951 2080 1971
rect 2100 1951 2120 1971
rect 2140 1951 2160 1971
rect 2180 1951 2200 1971
rect 2220 1951 2240 1971
rect 2260 1951 2280 1971
rect 2300 1951 2320 1971
rect 2340 1951 2360 1971
rect 2380 1951 2400 1971
rect 2420 1951 2440 1971
rect 2460 1951 2480 1971
rect 2500 1951 2520 1971
rect 2540 1951 2560 1971
rect 2580 1951 2600 1971
rect 2620 1951 2640 1971
rect 2660 1951 2675 1971
rect 175 1941 2675 1951
rect 0 1930 155 1940
rect 0 1910 10 1930
rect 30 1910 50 1930
rect 70 1910 90 1930
rect 110 1910 130 1930
rect 0 1900 155 1910
rect 175 1889 2675 1899
rect 175 1869 200 1889
rect 220 1869 240 1889
rect 260 1869 280 1889
rect 300 1869 320 1889
rect 340 1869 360 1889
rect 380 1869 400 1889
rect 420 1869 440 1889
rect 460 1869 480 1889
rect 500 1869 520 1889
rect 540 1869 560 1889
rect 580 1869 600 1889
rect 620 1869 640 1889
rect 660 1869 680 1889
rect 700 1869 720 1889
rect 740 1869 760 1889
rect 780 1869 800 1889
rect 820 1869 840 1889
rect 860 1869 880 1889
rect 900 1869 920 1889
rect 940 1869 960 1889
rect 980 1869 1000 1889
rect 1020 1869 1040 1889
rect 1060 1869 1080 1889
rect 1100 1869 1120 1889
rect 1140 1869 1160 1889
rect 1180 1869 1200 1889
rect 1220 1869 1240 1889
rect 1260 1869 1280 1889
rect 1300 1869 1320 1889
rect 1340 1869 1360 1889
rect 1380 1869 1400 1889
rect 1420 1869 1440 1889
rect 1460 1869 1480 1889
rect 1500 1869 1520 1889
rect 1540 1869 1560 1889
rect 1580 1869 1600 1889
rect 1620 1869 1640 1889
rect 1660 1869 1680 1889
rect 1700 1869 1720 1889
rect 1740 1869 1760 1889
rect 1780 1869 1800 1889
rect 1820 1869 1840 1889
rect 1860 1869 1880 1889
rect 1900 1869 1920 1889
rect 1940 1869 1960 1889
rect 1980 1869 2000 1889
rect 2020 1869 2040 1889
rect 2060 1869 2080 1889
rect 2100 1869 2120 1889
rect 2140 1869 2160 1889
rect 2180 1869 2200 1889
rect 2220 1869 2240 1889
rect 2260 1869 2280 1889
rect 2300 1869 2320 1889
rect 2340 1869 2360 1889
rect 2380 1869 2400 1889
rect 2420 1869 2440 1889
rect 2460 1869 2480 1889
rect 2500 1869 2520 1889
rect 2540 1869 2560 1889
rect 2580 1869 2600 1889
rect 2620 1869 2640 1889
rect 2660 1869 2675 1889
rect 0 1850 155 1860
rect 175 1859 2675 1869
rect 0 1830 10 1850
rect 30 1830 50 1850
rect 70 1830 90 1850
rect 110 1830 130 1850
rect 0 1820 155 1830
rect 175 1807 2675 1817
rect 175 1787 200 1807
rect 220 1787 240 1807
rect 260 1787 280 1807
rect 300 1787 320 1807
rect 340 1787 360 1807
rect 380 1787 400 1807
rect 420 1787 440 1807
rect 460 1787 480 1807
rect 500 1787 520 1807
rect 540 1787 560 1807
rect 580 1787 600 1807
rect 620 1787 640 1807
rect 660 1787 680 1807
rect 700 1787 720 1807
rect 740 1787 760 1807
rect 780 1787 800 1807
rect 820 1787 840 1807
rect 860 1787 880 1807
rect 900 1787 920 1807
rect 940 1787 960 1807
rect 980 1787 1000 1807
rect 1020 1787 1040 1807
rect 1060 1787 1080 1807
rect 1100 1787 1120 1807
rect 1140 1787 1160 1807
rect 1180 1787 1200 1807
rect 1220 1787 1240 1807
rect 1260 1787 1280 1807
rect 1300 1787 1320 1807
rect 1340 1787 1360 1807
rect 1380 1787 1400 1807
rect 1420 1787 1440 1807
rect 1460 1787 1480 1807
rect 1500 1787 1520 1807
rect 1540 1787 1560 1807
rect 1580 1787 1600 1807
rect 1620 1787 1640 1807
rect 1660 1787 1680 1807
rect 1700 1787 1720 1807
rect 1740 1787 1760 1807
rect 1780 1787 1800 1807
rect 1820 1787 1840 1807
rect 1860 1787 1880 1807
rect 1900 1787 1920 1807
rect 1940 1787 1960 1807
rect 1980 1787 2000 1807
rect 2020 1787 2040 1807
rect 2060 1787 2080 1807
rect 2100 1787 2120 1807
rect 2140 1787 2160 1807
rect 2180 1787 2200 1807
rect 2220 1787 2240 1807
rect 2260 1787 2280 1807
rect 2300 1787 2320 1807
rect 2340 1787 2360 1807
rect 2380 1787 2400 1807
rect 2420 1787 2440 1807
rect 2460 1787 2480 1807
rect 2500 1787 2520 1807
rect 2540 1787 2560 1807
rect 2580 1787 2600 1807
rect 2620 1787 2640 1807
rect 2660 1787 2675 1807
rect 175 1777 2675 1787
rect 0 1765 155 1775
rect 0 1745 10 1765
rect 30 1745 50 1765
rect 70 1745 90 1765
rect 110 1745 130 1765
rect 0 1735 155 1745
rect 175 1725 2675 1735
rect 175 1705 200 1725
rect 220 1705 240 1725
rect 260 1705 280 1725
rect 300 1705 320 1725
rect 340 1705 360 1725
rect 380 1705 400 1725
rect 420 1705 440 1725
rect 460 1705 480 1725
rect 500 1705 520 1725
rect 540 1705 560 1725
rect 580 1705 600 1725
rect 620 1705 640 1725
rect 660 1705 680 1725
rect 700 1705 720 1725
rect 740 1705 760 1725
rect 780 1705 800 1725
rect 820 1705 840 1725
rect 860 1705 880 1725
rect 900 1705 920 1725
rect 940 1705 960 1725
rect 980 1705 1000 1725
rect 1020 1705 1040 1725
rect 1060 1705 1080 1725
rect 1100 1705 1120 1725
rect 1140 1705 1160 1725
rect 1180 1705 1200 1725
rect 1220 1705 1240 1725
rect 1260 1705 1280 1725
rect 1300 1705 1320 1725
rect 1340 1705 1360 1725
rect 1380 1705 1400 1725
rect 1420 1705 1440 1725
rect 1460 1705 1480 1725
rect 1500 1705 1520 1725
rect 1540 1705 1560 1725
rect 1580 1705 1600 1725
rect 1620 1705 1640 1725
rect 1660 1705 1680 1725
rect 1700 1705 1720 1725
rect 1740 1705 1760 1725
rect 1780 1705 1800 1725
rect 1820 1705 1840 1725
rect 1860 1705 1880 1725
rect 1900 1705 1920 1725
rect 1940 1705 1960 1725
rect 1980 1705 2000 1725
rect 2020 1705 2040 1725
rect 2060 1705 2080 1725
rect 2100 1705 2120 1725
rect 2140 1705 2160 1725
rect 2180 1705 2200 1725
rect 2220 1705 2240 1725
rect 2260 1705 2280 1725
rect 2300 1705 2320 1725
rect 2340 1705 2360 1725
rect 2380 1705 2400 1725
rect 2420 1705 2440 1725
rect 2460 1705 2480 1725
rect 2500 1705 2520 1725
rect 2540 1705 2560 1725
rect 2580 1705 2600 1725
rect 2620 1705 2640 1725
rect 2660 1705 2675 1725
rect 175 1695 2675 1705
rect 0 1685 155 1695
rect 0 1665 10 1685
rect 30 1665 50 1685
rect 70 1665 90 1685
rect 110 1665 130 1685
rect 0 1655 155 1665
rect 175 1643 2675 1653
rect 175 1623 200 1643
rect 220 1623 240 1643
rect 260 1623 280 1643
rect 300 1623 320 1643
rect 340 1623 360 1643
rect 380 1623 400 1643
rect 420 1623 440 1643
rect 460 1623 480 1643
rect 500 1623 520 1643
rect 540 1623 560 1643
rect 580 1623 600 1643
rect 620 1623 640 1643
rect 660 1623 680 1643
rect 700 1623 720 1643
rect 740 1623 760 1643
rect 780 1623 800 1643
rect 820 1623 840 1643
rect 860 1623 880 1643
rect 900 1623 920 1643
rect 940 1623 960 1643
rect 980 1623 1000 1643
rect 1020 1623 1040 1643
rect 1060 1623 1080 1643
rect 1100 1623 1120 1643
rect 1140 1623 1160 1643
rect 1180 1623 1200 1643
rect 1220 1623 1240 1643
rect 1260 1623 1280 1643
rect 1300 1623 1320 1643
rect 1340 1623 1360 1643
rect 1380 1623 1400 1643
rect 1420 1623 1440 1643
rect 1460 1623 1480 1643
rect 1500 1623 1520 1643
rect 1540 1623 1560 1643
rect 1580 1623 1600 1643
rect 1620 1623 1640 1643
rect 1660 1623 1680 1643
rect 1700 1623 1720 1643
rect 1740 1623 1760 1643
rect 1780 1623 1800 1643
rect 1820 1623 1840 1643
rect 1860 1623 1880 1643
rect 1900 1623 1920 1643
rect 1940 1623 1960 1643
rect 1980 1623 2000 1643
rect 2020 1623 2040 1643
rect 2060 1623 2080 1643
rect 2100 1623 2120 1643
rect 2140 1623 2160 1643
rect 2180 1623 2200 1643
rect 2220 1623 2240 1643
rect 2260 1623 2280 1643
rect 2300 1623 2320 1643
rect 2340 1623 2360 1643
rect 2380 1623 2400 1643
rect 2420 1623 2440 1643
rect 2460 1623 2480 1643
rect 2500 1623 2520 1643
rect 2540 1623 2560 1643
rect 2580 1623 2600 1643
rect 2620 1623 2640 1643
rect 2660 1623 2675 1643
rect 175 1613 2675 1623
rect 0 1600 155 1610
rect 0 1580 10 1600
rect 30 1580 50 1600
rect 70 1580 90 1600
rect 110 1580 130 1600
rect 0 1570 155 1580
rect 175 1561 2675 1571
rect 175 1541 200 1561
rect 220 1541 240 1561
rect 260 1541 280 1561
rect 300 1541 320 1561
rect 340 1541 360 1561
rect 380 1541 400 1561
rect 420 1541 440 1561
rect 460 1541 480 1561
rect 500 1541 520 1561
rect 540 1541 560 1561
rect 580 1541 600 1561
rect 620 1541 640 1561
rect 660 1541 680 1561
rect 700 1541 720 1561
rect 740 1541 760 1561
rect 780 1541 800 1561
rect 820 1541 840 1561
rect 860 1541 880 1561
rect 900 1541 920 1561
rect 940 1541 960 1561
rect 980 1541 1000 1561
rect 1020 1541 1040 1561
rect 1060 1541 1080 1561
rect 1100 1541 1120 1561
rect 1140 1541 1160 1561
rect 1180 1541 1200 1561
rect 1220 1541 1240 1561
rect 1260 1541 1280 1561
rect 1300 1541 1320 1561
rect 1340 1541 1360 1561
rect 1380 1541 1400 1561
rect 1420 1541 1440 1561
rect 1460 1541 1480 1561
rect 1500 1541 1520 1561
rect 1540 1541 1560 1561
rect 1580 1541 1600 1561
rect 1620 1541 1640 1561
rect 1660 1541 1680 1561
rect 1700 1541 1720 1561
rect 1740 1541 1760 1561
rect 1780 1541 1800 1561
rect 1820 1541 1840 1561
rect 1860 1541 1880 1561
rect 1900 1541 1920 1561
rect 1940 1541 1960 1561
rect 1980 1541 2000 1561
rect 2020 1541 2040 1561
rect 2060 1541 2080 1561
rect 2100 1541 2120 1561
rect 2140 1541 2160 1561
rect 2180 1541 2200 1561
rect 2220 1541 2240 1561
rect 2260 1541 2280 1561
rect 2300 1541 2320 1561
rect 2340 1541 2360 1561
rect 2380 1541 2400 1561
rect 2420 1541 2440 1561
rect 2460 1541 2480 1561
rect 2500 1541 2520 1561
rect 2540 1541 2560 1561
rect 2580 1541 2600 1561
rect 2620 1541 2640 1561
rect 2660 1541 2675 1561
rect 175 1531 2675 1541
rect 0 1520 155 1530
rect 0 1500 10 1520
rect 30 1500 50 1520
rect 70 1500 90 1520
rect 110 1500 130 1520
rect 0 1490 155 1500
rect 175 1479 2675 1489
rect 175 1459 200 1479
rect 220 1459 240 1479
rect 260 1459 280 1479
rect 300 1459 320 1479
rect 340 1459 360 1479
rect 380 1459 400 1479
rect 420 1459 440 1479
rect 460 1459 480 1479
rect 500 1459 520 1479
rect 540 1459 560 1479
rect 580 1459 600 1479
rect 620 1459 640 1479
rect 660 1459 680 1479
rect 700 1459 720 1479
rect 740 1459 760 1479
rect 780 1459 800 1479
rect 820 1459 840 1479
rect 860 1459 880 1479
rect 900 1459 920 1479
rect 940 1459 960 1479
rect 980 1459 1000 1479
rect 1020 1459 1040 1479
rect 1060 1459 1080 1479
rect 1100 1459 1120 1479
rect 1140 1459 1160 1479
rect 1180 1459 1200 1479
rect 1220 1459 1240 1479
rect 1260 1459 1280 1479
rect 1300 1459 1320 1479
rect 1340 1459 1360 1479
rect 1380 1459 1400 1479
rect 1420 1459 1440 1479
rect 1460 1459 1480 1479
rect 1500 1459 1520 1479
rect 1540 1459 1560 1479
rect 1580 1459 1600 1479
rect 1620 1459 1640 1479
rect 1660 1459 1680 1479
rect 1700 1459 1720 1479
rect 1740 1459 1760 1479
rect 1780 1459 1800 1479
rect 1820 1459 1840 1479
rect 1860 1459 1880 1479
rect 1900 1459 1920 1479
rect 1940 1459 1960 1479
rect 1980 1459 2000 1479
rect 2020 1459 2040 1479
rect 2060 1459 2080 1479
rect 2100 1459 2120 1479
rect 2140 1459 2160 1479
rect 2180 1459 2200 1479
rect 2220 1459 2240 1479
rect 2260 1459 2280 1479
rect 2300 1459 2320 1479
rect 2340 1459 2360 1479
rect 2380 1459 2400 1479
rect 2420 1459 2440 1479
rect 2460 1459 2480 1479
rect 2500 1459 2520 1479
rect 2540 1459 2560 1479
rect 2580 1459 2600 1479
rect 2620 1459 2640 1479
rect 2660 1459 2675 1479
rect 0 1440 155 1450
rect 175 1449 2675 1459
rect 0 1420 10 1440
rect 30 1420 50 1440
rect 70 1420 90 1440
rect 110 1420 130 1440
rect 0 1410 155 1420
rect 175 1397 2675 1407
rect 175 1377 200 1397
rect 220 1377 240 1397
rect 260 1377 280 1397
rect 300 1377 320 1397
rect 340 1377 360 1397
rect 380 1377 400 1397
rect 420 1377 440 1397
rect 460 1377 480 1397
rect 500 1377 520 1397
rect 540 1377 560 1397
rect 580 1377 600 1397
rect 620 1377 640 1397
rect 660 1377 680 1397
rect 700 1377 720 1397
rect 740 1377 760 1397
rect 780 1377 800 1397
rect 820 1377 840 1397
rect 860 1377 880 1397
rect 900 1377 920 1397
rect 940 1377 960 1397
rect 980 1377 1000 1397
rect 1020 1377 1040 1397
rect 1060 1377 1080 1397
rect 1100 1377 1120 1397
rect 1140 1377 1160 1397
rect 1180 1377 1200 1397
rect 1220 1377 1240 1397
rect 1260 1377 1280 1397
rect 1300 1377 1320 1397
rect 1340 1377 1360 1397
rect 1380 1377 1400 1397
rect 1420 1377 1440 1397
rect 1460 1377 1480 1397
rect 1500 1377 1520 1397
rect 1540 1377 1560 1397
rect 1580 1377 1600 1397
rect 1620 1377 1640 1397
rect 1660 1377 1680 1397
rect 1700 1377 1720 1397
rect 1740 1377 1760 1397
rect 1780 1377 1800 1397
rect 1820 1377 1840 1397
rect 1860 1377 1880 1397
rect 1900 1377 1920 1397
rect 1940 1377 1960 1397
rect 1980 1377 2000 1397
rect 2020 1377 2040 1397
rect 2060 1377 2080 1397
rect 2100 1377 2120 1397
rect 2140 1377 2160 1397
rect 2180 1377 2200 1397
rect 2220 1377 2240 1397
rect 2260 1377 2280 1397
rect 2300 1377 2320 1397
rect 2340 1377 2360 1397
rect 2380 1377 2400 1397
rect 2420 1377 2440 1397
rect 2460 1377 2480 1397
rect 2500 1377 2520 1397
rect 2540 1377 2560 1397
rect 2580 1377 2600 1397
rect 2620 1377 2640 1397
rect 2660 1377 2675 1397
rect 175 1367 2675 1377
rect 0 1355 155 1365
rect 0 1335 10 1355
rect 30 1335 50 1355
rect 70 1335 90 1355
rect 110 1335 130 1355
rect 0 1325 155 1335
rect 175 1315 2675 1325
rect 175 1295 200 1315
rect 220 1295 240 1315
rect 260 1295 280 1315
rect 300 1295 320 1315
rect 340 1295 360 1315
rect 380 1295 400 1315
rect 420 1295 440 1315
rect 460 1295 480 1315
rect 500 1295 520 1315
rect 540 1295 560 1315
rect 580 1295 600 1315
rect 620 1295 640 1315
rect 660 1295 680 1315
rect 700 1295 720 1315
rect 740 1295 760 1315
rect 780 1295 800 1315
rect 820 1295 840 1315
rect 860 1295 880 1315
rect 900 1295 920 1315
rect 940 1295 960 1315
rect 980 1295 1000 1315
rect 1020 1295 1040 1315
rect 1060 1295 1080 1315
rect 1100 1295 1120 1315
rect 1140 1295 1160 1315
rect 1180 1295 1200 1315
rect 1220 1295 1240 1315
rect 1260 1295 1280 1315
rect 1300 1295 1320 1315
rect 1340 1295 1360 1315
rect 1380 1295 1400 1315
rect 1420 1295 1440 1315
rect 1460 1295 1480 1315
rect 1500 1295 1520 1315
rect 1540 1295 1560 1315
rect 1580 1295 1600 1315
rect 1620 1295 1640 1315
rect 1660 1295 1680 1315
rect 1700 1295 1720 1315
rect 1740 1295 1760 1315
rect 1780 1295 1800 1315
rect 1820 1295 1840 1315
rect 1860 1295 1880 1315
rect 1900 1295 1920 1315
rect 1940 1295 1960 1315
rect 1980 1295 2000 1315
rect 2020 1295 2040 1315
rect 2060 1295 2080 1315
rect 2100 1295 2120 1315
rect 2140 1295 2160 1315
rect 2180 1295 2200 1315
rect 2220 1295 2240 1315
rect 2260 1295 2280 1315
rect 2300 1295 2320 1315
rect 2340 1295 2360 1315
rect 2380 1295 2400 1315
rect 2420 1295 2440 1315
rect 2460 1295 2480 1315
rect 2500 1295 2520 1315
rect 2540 1295 2560 1315
rect 2580 1295 2600 1315
rect 2620 1295 2640 1315
rect 2660 1295 2675 1315
rect 175 1285 2675 1295
rect 0 1275 155 1285
rect 0 1255 10 1275
rect 30 1255 50 1275
rect 70 1255 90 1275
rect 110 1255 130 1275
rect 0 1245 155 1255
rect 175 1233 2675 1243
rect 175 1213 200 1233
rect 220 1213 240 1233
rect 260 1213 280 1233
rect 300 1213 320 1233
rect 340 1213 360 1233
rect 380 1213 400 1233
rect 420 1213 440 1233
rect 460 1213 480 1233
rect 500 1213 520 1233
rect 540 1213 560 1233
rect 580 1213 600 1233
rect 620 1213 640 1233
rect 660 1213 680 1233
rect 700 1213 720 1233
rect 740 1213 760 1233
rect 780 1213 800 1233
rect 820 1213 840 1233
rect 860 1213 880 1233
rect 900 1213 920 1233
rect 940 1213 960 1233
rect 980 1213 1000 1233
rect 1020 1213 1040 1233
rect 1060 1213 1080 1233
rect 1100 1213 1120 1233
rect 1140 1213 1160 1233
rect 1180 1213 1200 1233
rect 1220 1213 1240 1233
rect 1260 1213 1280 1233
rect 1300 1213 1320 1233
rect 1340 1213 1360 1233
rect 1380 1213 1400 1233
rect 1420 1213 1440 1233
rect 1460 1213 1480 1233
rect 1500 1213 1520 1233
rect 1540 1213 1560 1233
rect 1580 1213 1600 1233
rect 1620 1213 1640 1233
rect 1660 1213 1680 1233
rect 1700 1213 1720 1233
rect 1740 1213 1760 1233
rect 1780 1213 1800 1233
rect 1820 1213 1840 1233
rect 1860 1213 1880 1233
rect 1900 1213 1920 1233
rect 1940 1213 1960 1233
rect 1980 1213 2000 1233
rect 2020 1213 2040 1233
rect 2060 1213 2080 1233
rect 2100 1213 2120 1233
rect 2140 1213 2160 1233
rect 2180 1213 2200 1233
rect 2220 1213 2240 1233
rect 2260 1213 2280 1233
rect 2300 1213 2320 1233
rect 2340 1213 2360 1233
rect 2380 1213 2400 1233
rect 2420 1213 2440 1233
rect 2460 1213 2480 1233
rect 2500 1213 2520 1233
rect 2540 1213 2560 1233
rect 2580 1213 2600 1233
rect 2620 1213 2640 1233
rect 2660 1213 2675 1233
rect 175 1203 2675 1213
rect 0 1190 155 1200
rect 0 1170 10 1190
rect 30 1170 50 1190
rect 70 1170 90 1190
rect 110 1170 130 1190
rect 0 1160 155 1170
rect 175 1151 2675 1161
rect 175 1131 200 1151
rect 220 1131 240 1151
rect 260 1131 280 1151
rect 300 1131 320 1151
rect 340 1131 360 1151
rect 380 1131 400 1151
rect 420 1131 440 1151
rect 460 1131 480 1151
rect 500 1131 520 1151
rect 540 1131 560 1151
rect 580 1131 600 1151
rect 620 1131 640 1151
rect 660 1131 680 1151
rect 700 1131 720 1151
rect 740 1131 760 1151
rect 780 1131 800 1151
rect 820 1131 840 1151
rect 860 1131 880 1151
rect 900 1131 920 1151
rect 940 1131 960 1151
rect 980 1131 1000 1151
rect 1020 1131 1040 1151
rect 1060 1131 1080 1151
rect 1100 1131 1120 1151
rect 1140 1131 1160 1151
rect 1180 1131 1200 1151
rect 1220 1131 1240 1151
rect 1260 1131 1280 1151
rect 1300 1131 1320 1151
rect 1340 1131 1360 1151
rect 1380 1131 1400 1151
rect 1420 1131 1440 1151
rect 1460 1131 1480 1151
rect 1500 1131 1520 1151
rect 1540 1131 1560 1151
rect 1580 1131 1600 1151
rect 1620 1131 1640 1151
rect 1660 1131 1680 1151
rect 1700 1131 1720 1151
rect 1740 1131 1760 1151
rect 1780 1131 1800 1151
rect 1820 1131 1840 1151
rect 1860 1131 1880 1151
rect 1900 1131 1920 1151
rect 1940 1131 1960 1151
rect 1980 1131 2000 1151
rect 2020 1131 2040 1151
rect 2060 1131 2080 1151
rect 2100 1131 2120 1151
rect 2140 1131 2160 1151
rect 2180 1131 2200 1151
rect 2220 1131 2240 1151
rect 2260 1131 2280 1151
rect 2300 1131 2320 1151
rect 2340 1131 2360 1151
rect 2380 1131 2400 1151
rect 2420 1131 2440 1151
rect 2460 1131 2480 1151
rect 2500 1131 2520 1151
rect 2540 1131 2560 1151
rect 2580 1131 2600 1151
rect 2620 1131 2640 1151
rect 2660 1131 2675 1151
rect 175 1121 2675 1131
rect 0 1110 155 1120
rect 0 1090 10 1110
rect 30 1090 50 1110
rect 70 1090 90 1110
rect 110 1090 130 1110
rect 0 1080 155 1090
rect 175 1069 2675 1079
rect 175 1049 200 1069
rect 220 1049 240 1069
rect 260 1049 280 1069
rect 300 1049 320 1069
rect 340 1049 360 1069
rect 380 1049 400 1069
rect 420 1049 440 1069
rect 460 1049 480 1069
rect 500 1049 520 1069
rect 540 1049 560 1069
rect 580 1049 600 1069
rect 620 1049 640 1069
rect 660 1049 680 1069
rect 700 1049 720 1069
rect 740 1049 760 1069
rect 780 1049 800 1069
rect 820 1049 840 1069
rect 860 1049 880 1069
rect 900 1049 920 1069
rect 940 1049 960 1069
rect 980 1049 1000 1069
rect 1020 1049 1040 1069
rect 1060 1049 1080 1069
rect 1100 1049 1120 1069
rect 1140 1049 1160 1069
rect 1180 1049 1200 1069
rect 1220 1049 1240 1069
rect 1260 1049 1280 1069
rect 1300 1049 1320 1069
rect 1340 1049 1360 1069
rect 1380 1049 1400 1069
rect 1420 1049 1440 1069
rect 1460 1049 1480 1069
rect 1500 1049 1520 1069
rect 1540 1049 1560 1069
rect 1580 1049 1600 1069
rect 1620 1049 1640 1069
rect 1660 1049 1680 1069
rect 1700 1049 1720 1069
rect 1740 1049 1760 1069
rect 1780 1049 1800 1069
rect 1820 1049 1840 1069
rect 1860 1049 1880 1069
rect 1900 1049 1920 1069
rect 1940 1049 1960 1069
rect 1980 1049 2000 1069
rect 2020 1049 2040 1069
rect 2060 1049 2080 1069
rect 2100 1049 2120 1069
rect 2140 1049 2160 1069
rect 2180 1049 2200 1069
rect 2220 1049 2240 1069
rect 2260 1049 2280 1069
rect 2300 1049 2320 1069
rect 2340 1049 2360 1069
rect 2380 1049 2400 1069
rect 2420 1049 2440 1069
rect 2460 1049 2480 1069
rect 2500 1049 2520 1069
rect 2540 1049 2560 1069
rect 2580 1049 2600 1069
rect 2620 1049 2640 1069
rect 2660 1049 2675 1069
rect 0 1030 155 1040
rect 175 1039 2675 1049
rect 0 1010 10 1030
rect 30 1010 50 1030
rect 70 1010 90 1030
rect 110 1010 130 1030
rect 0 1000 155 1010
rect 175 987 2675 997
rect 175 967 200 987
rect 220 967 240 987
rect 260 967 280 987
rect 300 967 320 987
rect 340 967 360 987
rect 380 967 400 987
rect 420 967 440 987
rect 460 967 480 987
rect 500 967 520 987
rect 540 967 560 987
rect 580 967 600 987
rect 620 967 640 987
rect 660 967 680 987
rect 700 967 720 987
rect 740 967 760 987
rect 780 967 800 987
rect 820 967 840 987
rect 860 967 880 987
rect 900 967 920 987
rect 940 967 960 987
rect 980 967 1000 987
rect 1020 967 1040 987
rect 1060 967 1080 987
rect 1100 967 1120 987
rect 1140 967 1160 987
rect 1180 967 1200 987
rect 1220 967 1240 987
rect 1260 967 1280 987
rect 1300 967 1320 987
rect 1340 967 1360 987
rect 1380 967 1400 987
rect 1420 967 1440 987
rect 1460 967 1480 987
rect 1500 967 1520 987
rect 1540 967 1560 987
rect 1580 967 1600 987
rect 1620 967 1640 987
rect 1660 967 1680 987
rect 1700 967 1720 987
rect 1740 967 1760 987
rect 1780 967 1800 987
rect 1820 967 1840 987
rect 1860 967 1880 987
rect 1900 967 1920 987
rect 1940 967 1960 987
rect 1980 967 2000 987
rect 2020 967 2040 987
rect 2060 967 2080 987
rect 2100 967 2120 987
rect 2140 967 2160 987
rect 2180 967 2200 987
rect 2220 967 2240 987
rect 2260 967 2280 987
rect 2300 967 2320 987
rect 2340 967 2360 987
rect 2380 967 2400 987
rect 2420 967 2440 987
rect 2460 967 2480 987
rect 2500 967 2520 987
rect 2540 967 2560 987
rect 2580 967 2600 987
rect 2620 967 2640 987
rect 2660 967 2675 987
rect 175 957 2675 967
rect 0 945 155 955
rect 0 925 10 945
rect 30 925 50 945
rect 70 925 90 945
rect 110 925 130 945
rect 0 915 155 925
rect 175 905 2675 915
rect 175 885 200 905
rect 220 885 240 905
rect 260 885 280 905
rect 300 885 320 905
rect 340 885 360 905
rect 380 885 400 905
rect 420 885 440 905
rect 460 885 480 905
rect 500 885 520 905
rect 540 885 560 905
rect 580 885 600 905
rect 620 885 640 905
rect 660 885 680 905
rect 700 885 720 905
rect 740 885 760 905
rect 780 885 800 905
rect 820 885 840 905
rect 860 885 880 905
rect 900 885 920 905
rect 940 885 960 905
rect 980 885 1000 905
rect 1020 885 1040 905
rect 1060 885 1080 905
rect 1100 885 1120 905
rect 1140 885 1160 905
rect 1180 885 1200 905
rect 1220 885 1240 905
rect 1260 885 1280 905
rect 1300 885 1320 905
rect 1340 885 1360 905
rect 1380 885 1400 905
rect 1420 885 1440 905
rect 1460 885 1480 905
rect 1500 885 1520 905
rect 1540 885 1560 905
rect 1580 885 1600 905
rect 1620 885 1640 905
rect 1660 885 1680 905
rect 1700 885 1720 905
rect 1740 885 1760 905
rect 1780 885 1800 905
rect 1820 885 1840 905
rect 1860 885 1880 905
rect 1900 885 1920 905
rect 1940 885 1960 905
rect 1980 885 2000 905
rect 2020 885 2040 905
rect 2060 885 2080 905
rect 2100 885 2120 905
rect 2140 885 2160 905
rect 2180 885 2200 905
rect 2220 885 2240 905
rect 2260 885 2280 905
rect 2300 885 2320 905
rect 2340 885 2360 905
rect 2380 885 2400 905
rect 2420 885 2440 905
rect 2460 885 2480 905
rect 2500 885 2520 905
rect 2540 885 2560 905
rect 2580 885 2600 905
rect 2620 885 2640 905
rect 2660 885 2675 905
rect 175 875 2675 885
rect 0 865 155 875
rect 0 845 10 865
rect 30 845 50 865
rect 70 845 90 865
rect 110 845 130 865
rect 0 835 155 845
rect 175 823 2675 833
rect 175 803 200 823
rect 220 803 240 823
rect 260 803 280 823
rect 300 803 320 823
rect 340 803 360 823
rect 380 803 400 823
rect 420 803 440 823
rect 460 803 480 823
rect 500 803 520 823
rect 540 803 560 823
rect 580 803 600 823
rect 620 803 640 823
rect 660 803 680 823
rect 700 803 720 823
rect 740 803 760 823
rect 780 803 800 823
rect 820 803 840 823
rect 860 803 880 823
rect 900 803 920 823
rect 940 803 960 823
rect 980 803 1000 823
rect 1020 803 1040 823
rect 1060 803 1080 823
rect 1100 803 1120 823
rect 1140 803 1160 823
rect 1180 803 1200 823
rect 1220 803 1240 823
rect 1260 803 1280 823
rect 1300 803 1320 823
rect 1340 803 1360 823
rect 1380 803 1400 823
rect 1420 803 1440 823
rect 1460 803 1480 823
rect 1500 803 1520 823
rect 1540 803 1560 823
rect 1580 803 1600 823
rect 1620 803 1640 823
rect 1660 803 1680 823
rect 1700 803 1720 823
rect 1740 803 1760 823
rect 1780 803 1800 823
rect 1820 803 1840 823
rect 1860 803 1880 823
rect 1900 803 1920 823
rect 1940 803 1960 823
rect 1980 803 2000 823
rect 2020 803 2040 823
rect 2060 803 2080 823
rect 2100 803 2120 823
rect 2140 803 2160 823
rect 2180 803 2200 823
rect 2220 803 2240 823
rect 2260 803 2280 823
rect 2300 803 2320 823
rect 2340 803 2360 823
rect 2380 803 2400 823
rect 2420 803 2440 823
rect 2460 803 2480 823
rect 2500 803 2520 823
rect 2540 803 2560 823
rect 2580 803 2600 823
rect 2620 803 2640 823
rect 2660 803 2675 823
rect 175 793 2675 803
rect 0 780 155 790
rect 0 760 10 780
rect 30 760 50 780
rect 70 760 90 780
rect 110 760 130 780
rect 0 750 155 760
rect 175 741 2675 751
rect 175 721 200 741
rect 220 721 240 741
rect 260 721 280 741
rect 300 721 320 741
rect 340 721 360 741
rect 380 721 400 741
rect 420 721 440 741
rect 460 721 480 741
rect 500 721 520 741
rect 540 721 560 741
rect 580 721 600 741
rect 620 721 640 741
rect 660 721 680 741
rect 700 721 720 741
rect 740 721 760 741
rect 780 721 800 741
rect 820 721 840 741
rect 860 721 880 741
rect 900 721 920 741
rect 940 721 960 741
rect 980 721 1000 741
rect 1020 721 1040 741
rect 1060 721 1080 741
rect 1100 721 1120 741
rect 1140 721 1160 741
rect 1180 721 1200 741
rect 1220 721 1240 741
rect 1260 721 1280 741
rect 1300 721 1320 741
rect 1340 721 1360 741
rect 1380 721 1400 741
rect 1420 721 1440 741
rect 1460 721 1480 741
rect 1500 721 1520 741
rect 1540 721 1560 741
rect 1580 721 1600 741
rect 1620 721 1640 741
rect 1660 721 1680 741
rect 1700 721 1720 741
rect 1740 721 1760 741
rect 1780 721 1800 741
rect 1820 721 1840 741
rect 1860 721 1880 741
rect 1900 721 1920 741
rect 1940 721 1960 741
rect 1980 721 2000 741
rect 2020 721 2040 741
rect 2060 721 2080 741
rect 2100 721 2120 741
rect 2140 721 2160 741
rect 2180 721 2200 741
rect 2220 721 2240 741
rect 2260 721 2280 741
rect 2300 721 2320 741
rect 2340 721 2360 741
rect 2380 721 2400 741
rect 2420 721 2440 741
rect 2460 721 2480 741
rect 2500 721 2520 741
rect 2540 721 2560 741
rect 2580 721 2600 741
rect 2620 721 2640 741
rect 2660 721 2675 741
rect 175 711 2675 721
rect 0 700 155 710
rect 0 680 10 700
rect 30 680 50 700
rect 70 680 90 700
rect 110 680 130 700
rect 0 670 155 680
rect 175 659 2675 669
rect 175 639 200 659
rect 220 639 240 659
rect 260 639 280 659
rect 300 639 320 659
rect 340 639 360 659
rect 380 639 400 659
rect 420 639 440 659
rect 460 639 480 659
rect 500 639 520 659
rect 540 639 560 659
rect 580 639 600 659
rect 620 639 640 659
rect 660 639 680 659
rect 700 639 720 659
rect 740 639 760 659
rect 780 639 800 659
rect 820 639 840 659
rect 860 639 880 659
rect 900 639 920 659
rect 940 639 960 659
rect 980 639 1000 659
rect 1020 639 1040 659
rect 1060 639 1080 659
rect 1100 639 1120 659
rect 1140 639 1160 659
rect 1180 639 1200 659
rect 1220 639 1240 659
rect 1260 639 1280 659
rect 1300 639 1320 659
rect 1340 639 1360 659
rect 1380 639 1400 659
rect 1420 639 1440 659
rect 1460 639 1480 659
rect 1500 639 1520 659
rect 1540 639 1560 659
rect 1580 639 1600 659
rect 1620 639 1640 659
rect 1660 639 1680 659
rect 1700 639 1720 659
rect 1740 639 1760 659
rect 1780 639 1800 659
rect 1820 639 1840 659
rect 1860 639 1880 659
rect 1900 639 1920 659
rect 1940 639 1960 659
rect 1980 639 2000 659
rect 2020 639 2040 659
rect 2060 639 2080 659
rect 2100 639 2120 659
rect 2140 639 2160 659
rect 2180 639 2200 659
rect 2220 639 2240 659
rect 2260 639 2280 659
rect 2300 639 2320 659
rect 2340 639 2360 659
rect 2380 639 2400 659
rect 2420 639 2440 659
rect 2460 639 2480 659
rect 2500 639 2520 659
rect 2540 639 2560 659
rect 2580 639 2600 659
rect 2620 639 2640 659
rect 2660 639 2675 659
rect 0 620 155 630
rect 175 629 2675 639
rect 0 600 10 620
rect 30 600 50 620
rect 70 600 90 620
rect 110 600 130 620
rect 0 590 155 600
rect 175 577 2675 587
rect 175 557 200 577
rect 220 557 240 577
rect 260 557 280 577
rect 300 557 320 577
rect 340 557 360 577
rect 380 557 400 577
rect 420 557 440 577
rect 460 557 480 577
rect 500 557 520 577
rect 540 557 560 577
rect 580 557 600 577
rect 620 557 640 577
rect 660 557 680 577
rect 700 557 720 577
rect 740 557 760 577
rect 780 557 800 577
rect 820 557 840 577
rect 860 557 880 577
rect 900 557 920 577
rect 940 557 960 577
rect 980 557 1000 577
rect 1020 557 1040 577
rect 1060 557 1080 577
rect 1100 557 1120 577
rect 1140 557 1160 577
rect 1180 557 1200 577
rect 1220 557 1240 577
rect 1260 557 1280 577
rect 1300 557 1320 577
rect 1340 557 1360 577
rect 1380 557 1400 577
rect 1420 557 1440 577
rect 1460 557 1480 577
rect 1500 557 1520 577
rect 1540 557 1560 577
rect 1580 557 1600 577
rect 1620 557 1640 577
rect 1660 557 1680 577
rect 1700 557 1720 577
rect 1740 557 1760 577
rect 1780 557 1800 577
rect 1820 557 1840 577
rect 1860 557 1880 577
rect 1900 557 1920 577
rect 1940 557 1960 577
rect 1980 557 2000 577
rect 2020 557 2040 577
rect 2060 557 2080 577
rect 2100 557 2120 577
rect 2140 557 2160 577
rect 2180 557 2200 577
rect 2220 557 2240 577
rect 2260 557 2280 577
rect 2300 557 2320 577
rect 2340 557 2360 577
rect 2380 557 2400 577
rect 2420 557 2440 577
rect 2460 557 2480 577
rect 2500 557 2520 577
rect 2540 557 2560 577
rect 2580 557 2600 577
rect 2620 557 2640 577
rect 2660 557 2675 577
rect 175 547 2675 557
rect 0 535 155 545
rect 0 515 10 535
rect 30 515 50 535
rect 70 515 90 535
rect 110 515 130 535
rect 0 505 155 515
rect 175 495 2675 505
rect 175 475 200 495
rect 220 475 240 495
rect 260 475 280 495
rect 300 475 320 495
rect 340 475 360 495
rect 380 475 400 495
rect 420 475 440 495
rect 460 475 480 495
rect 500 475 520 495
rect 540 475 560 495
rect 580 475 600 495
rect 620 475 640 495
rect 660 475 680 495
rect 700 475 720 495
rect 740 475 760 495
rect 780 475 800 495
rect 820 475 840 495
rect 860 475 880 495
rect 900 475 920 495
rect 940 475 960 495
rect 980 475 1000 495
rect 1020 475 1040 495
rect 1060 475 1080 495
rect 1100 475 1120 495
rect 1140 475 1160 495
rect 1180 475 1200 495
rect 1220 475 1240 495
rect 1260 475 1280 495
rect 1300 475 1320 495
rect 1340 475 1360 495
rect 1380 475 1400 495
rect 1420 475 1440 495
rect 1460 475 1480 495
rect 1500 475 1520 495
rect 1540 475 1560 495
rect 1580 475 1600 495
rect 1620 475 1640 495
rect 1660 475 1680 495
rect 1700 475 1720 495
rect 1740 475 1760 495
rect 1780 475 1800 495
rect 1820 475 1840 495
rect 1860 475 1880 495
rect 1900 475 1920 495
rect 1940 475 1960 495
rect 1980 475 2000 495
rect 2020 475 2040 495
rect 2060 475 2080 495
rect 2100 475 2120 495
rect 2140 475 2160 495
rect 2180 475 2200 495
rect 2220 475 2240 495
rect 2260 475 2280 495
rect 2300 475 2320 495
rect 2340 475 2360 495
rect 2380 475 2400 495
rect 2420 475 2440 495
rect 2460 475 2480 495
rect 2500 475 2520 495
rect 2540 475 2560 495
rect 2580 475 2600 495
rect 2620 475 2640 495
rect 2660 475 2675 495
rect 175 465 2675 475
rect 0 455 155 465
rect 0 435 10 455
rect 30 435 50 455
rect 70 435 90 455
rect 110 435 130 455
rect 0 425 155 435
rect 175 413 2675 423
rect 175 393 200 413
rect 220 393 240 413
rect 260 393 280 413
rect 300 393 320 413
rect 340 393 360 413
rect 380 393 400 413
rect 420 393 440 413
rect 460 393 480 413
rect 500 393 520 413
rect 540 393 560 413
rect 580 393 600 413
rect 620 393 640 413
rect 660 393 680 413
rect 700 393 720 413
rect 740 393 760 413
rect 780 393 800 413
rect 820 393 840 413
rect 860 393 880 413
rect 900 393 920 413
rect 940 393 960 413
rect 980 393 1000 413
rect 1020 393 1040 413
rect 1060 393 1080 413
rect 1100 393 1120 413
rect 1140 393 1160 413
rect 1180 393 1200 413
rect 1220 393 1240 413
rect 1260 393 1280 413
rect 1300 393 1320 413
rect 1340 393 1360 413
rect 1380 393 1400 413
rect 1420 393 1440 413
rect 1460 393 1480 413
rect 1500 393 1520 413
rect 1540 393 1560 413
rect 1580 393 1600 413
rect 1620 393 1640 413
rect 1660 393 1680 413
rect 1700 393 1720 413
rect 1740 393 1760 413
rect 1780 393 1800 413
rect 1820 393 1840 413
rect 1860 393 1880 413
rect 1900 393 1920 413
rect 1940 393 1960 413
rect 1980 393 2000 413
rect 2020 393 2040 413
rect 2060 393 2080 413
rect 2100 393 2120 413
rect 2140 393 2160 413
rect 2180 393 2200 413
rect 2220 393 2240 413
rect 2260 393 2280 413
rect 2300 393 2320 413
rect 2340 393 2360 413
rect 2380 393 2400 413
rect 2420 393 2440 413
rect 2460 393 2480 413
rect 2500 393 2520 413
rect 2540 393 2560 413
rect 2580 393 2600 413
rect 2620 393 2640 413
rect 2660 393 2675 413
rect 0 375 155 385
rect 175 383 2675 393
rect 0 355 10 375
rect 30 355 50 375
rect 70 355 90 375
rect 110 355 130 375
rect 0 345 155 355
rect 175 331 2675 341
rect 175 311 200 331
rect 220 311 240 331
rect 260 311 280 331
rect 300 311 320 331
rect 340 311 360 331
rect 380 311 400 331
rect 420 311 440 331
rect 460 311 480 331
rect 500 311 520 331
rect 540 311 560 331
rect 580 311 600 331
rect 620 311 640 331
rect 660 311 680 331
rect 700 311 720 331
rect 740 311 760 331
rect 780 311 800 331
rect 820 311 840 331
rect 860 311 880 331
rect 900 311 920 331
rect 940 311 960 331
rect 980 311 1000 331
rect 1020 311 1040 331
rect 1060 311 1080 331
rect 1100 311 1120 331
rect 1140 311 1160 331
rect 1180 311 1200 331
rect 1220 311 1240 331
rect 1260 311 1280 331
rect 1300 311 1320 331
rect 1340 311 1360 331
rect 1380 311 1400 331
rect 1420 311 1440 331
rect 1460 311 1480 331
rect 1500 311 1520 331
rect 1540 311 1560 331
rect 1580 311 1600 331
rect 1620 311 1640 331
rect 1660 311 1680 331
rect 1700 311 1720 331
rect 1740 311 1760 331
rect 1780 311 1800 331
rect 1820 311 1840 331
rect 1860 311 1880 331
rect 1900 311 1920 331
rect 1940 311 1960 331
rect 1980 311 2000 331
rect 2020 311 2040 331
rect 2060 311 2080 331
rect 2100 311 2120 331
rect 2140 311 2160 331
rect 2180 311 2200 331
rect 2220 311 2240 331
rect 2260 311 2280 331
rect 2300 311 2320 331
rect 2340 311 2360 331
rect 2380 311 2400 331
rect 2420 311 2440 331
rect 2460 311 2480 331
rect 2500 311 2520 331
rect 2540 311 2560 331
rect 2580 311 2600 331
rect 2620 311 2640 331
rect 2660 311 2675 331
rect 175 301 2675 311
rect 0 290 155 300
rect 0 270 10 290
rect 30 270 50 290
rect 70 270 90 290
rect 110 270 130 290
rect 0 260 155 270
rect 175 249 2675 259
rect 175 229 200 249
rect 220 229 240 249
rect 260 229 280 249
rect 300 229 320 249
rect 340 229 360 249
rect 380 229 400 249
rect 420 229 440 249
rect 460 229 480 249
rect 500 229 520 249
rect 540 229 560 249
rect 580 229 600 249
rect 620 229 640 249
rect 660 229 680 249
rect 700 229 720 249
rect 740 229 760 249
rect 780 229 800 249
rect 820 229 840 249
rect 860 229 880 249
rect 900 229 920 249
rect 940 229 960 249
rect 980 229 1000 249
rect 1020 229 1040 249
rect 1060 229 1080 249
rect 1100 229 1120 249
rect 1140 229 1160 249
rect 1180 229 1200 249
rect 1220 229 1240 249
rect 1260 229 1280 249
rect 1300 229 1320 249
rect 1340 229 1360 249
rect 1380 229 1400 249
rect 1420 229 1440 249
rect 1460 229 1480 249
rect 1500 229 1520 249
rect 1540 229 1560 249
rect 1580 229 1600 249
rect 1620 229 1640 249
rect 1660 229 1680 249
rect 1700 229 1720 249
rect 1740 229 1760 249
rect 1780 229 1800 249
rect 1820 229 1840 249
rect 1860 229 1880 249
rect 1900 229 1920 249
rect 1940 229 1960 249
rect 1980 229 2000 249
rect 2020 229 2040 249
rect 2060 229 2080 249
rect 2100 229 2120 249
rect 2140 229 2160 249
rect 2180 229 2200 249
rect 2220 229 2240 249
rect 2260 229 2280 249
rect 2300 229 2320 249
rect 2340 229 2360 249
rect 2380 229 2400 249
rect 2420 229 2440 249
rect 2460 229 2480 249
rect 2500 229 2520 249
rect 2540 229 2560 249
rect 2580 229 2600 249
rect 2620 229 2640 249
rect 2660 229 2675 249
rect 0 210 155 220
rect 175 219 2675 229
rect 0 190 10 210
rect 30 190 50 210
rect 70 190 90 210
rect 110 190 130 210
rect 0 180 155 190
rect 175 167 2675 177
rect 175 147 200 167
rect 220 147 240 167
rect 260 147 280 167
rect 300 147 320 167
rect 340 147 360 167
rect 380 147 400 167
rect 420 147 440 167
rect 460 147 480 167
rect 500 147 520 167
rect 540 147 560 167
rect 580 147 600 167
rect 620 147 640 167
rect 660 147 680 167
rect 700 147 720 167
rect 740 147 760 167
rect 780 147 800 167
rect 820 147 840 167
rect 860 147 880 167
rect 900 147 920 167
rect 940 147 960 167
rect 980 147 1000 167
rect 1020 147 1040 167
rect 1060 147 1080 167
rect 1100 147 1120 167
rect 1140 147 1160 167
rect 1180 147 1200 167
rect 1220 147 1240 167
rect 1260 147 1280 167
rect 1300 147 1320 167
rect 1340 147 1360 167
rect 1380 147 1400 167
rect 1420 147 1440 167
rect 1460 147 1480 167
rect 1500 147 1520 167
rect 1540 147 1560 167
rect 1580 147 1600 167
rect 1620 147 1640 167
rect 1660 147 1680 167
rect 1700 147 1720 167
rect 1740 147 1760 167
rect 1780 147 1800 167
rect 1820 147 1840 167
rect 1860 147 1880 167
rect 1900 147 1920 167
rect 1940 147 1960 167
rect 1980 147 2000 167
rect 2020 147 2040 167
rect 2060 147 2080 167
rect 2100 147 2120 167
rect 2140 147 2160 167
rect 2180 147 2200 167
rect 2220 147 2240 167
rect 2260 147 2280 167
rect 2300 147 2320 167
rect 2340 147 2360 167
rect 2380 147 2400 167
rect 2420 147 2440 167
rect 2460 147 2480 167
rect 2500 147 2520 167
rect 2540 147 2560 167
rect 2580 147 2600 167
rect 2620 147 2640 167
rect 2660 147 2675 167
rect 0 130 155 140
rect 175 137 2675 147
rect 0 110 10 130
rect 30 110 50 130
rect 70 110 90 130
rect 110 110 130 130
rect 0 100 155 110
rect 175 85 2675 95
rect 175 65 200 85
rect 220 65 240 85
rect 260 65 280 85
rect 300 65 320 85
rect 340 65 360 85
rect 380 65 400 85
rect 420 65 440 85
rect 460 65 480 85
rect 500 65 520 85
rect 540 65 560 85
rect 580 65 600 85
rect 620 65 640 85
rect 660 65 680 85
rect 700 65 720 85
rect 740 65 760 85
rect 780 65 800 85
rect 820 65 840 85
rect 860 65 880 85
rect 900 65 920 85
rect 940 65 960 85
rect 980 65 1000 85
rect 1020 65 1040 85
rect 1060 65 1080 85
rect 1100 65 1120 85
rect 1140 65 1160 85
rect 1180 65 1200 85
rect 1220 65 1240 85
rect 1260 65 1280 85
rect 1300 65 1320 85
rect 1340 65 1360 85
rect 1380 65 1400 85
rect 1420 65 1440 85
rect 1460 65 1480 85
rect 1500 65 1520 85
rect 1540 65 1560 85
rect 1580 65 1600 85
rect 1620 65 1640 85
rect 1660 65 1680 85
rect 1700 65 1720 85
rect 1740 65 1760 85
rect 1780 65 1800 85
rect 1820 65 1840 85
rect 1860 65 1880 85
rect 1900 65 1920 85
rect 1940 65 1960 85
rect 1980 65 2000 85
rect 2020 65 2040 85
rect 2060 65 2080 85
rect 2100 65 2120 85
rect 2140 65 2160 85
rect 2180 65 2200 85
rect 2220 65 2240 85
rect 2260 65 2280 85
rect 2300 65 2320 85
rect 2340 65 2360 85
rect 2380 65 2400 85
rect 2420 65 2440 85
rect 2460 65 2480 85
rect 2500 65 2520 85
rect 2540 65 2560 85
rect 2580 65 2600 85
rect 2620 65 2640 85
rect 2660 65 2675 85
rect 175 45 2675 65
rect 175 25 200 45
rect 220 25 240 45
rect 260 25 280 45
rect 300 25 320 45
rect 340 25 360 45
rect 380 25 400 45
rect 420 25 440 45
rect 460 25 480 45
rect 500 25 520 45
rect 540 25 560 45
rect 580 25 600 45
rect 620 25 640 45
rect 660 25 680 45
rect 700 25 720 45
rect 740 25 760 45
rect 780 25 800 45
rect 820 25 840 45
rect 860 25 880 45
rect 900 25 920 45
rect 940 25 960 45
rect 980 25 1000 45
rect 1020 25 1040 45
rect 1060 25 1080 45
rect 1100 25 1120 45
rect 1140 25 1160 45
rect 1180 25 1200 45
rect 1220 25 1240 45
rect 1260 25 1280 45
rect 1300 25 1320 45
rect 1340 25 1360 45
rect 1380 25 1400 45
rect 1420 25 1440 45
rect 1460 25 1480 45
rect 1500 25 1520 45
rect 1540 25 1560 45
rect 1580 25 1600 45
rect 1620 25 1640 45
rect 1660 25 1680 45
rect 1700 25 1720 45
rect 1740 25 1760 45
rect 1780 25 1800 45
rect 1820 25 1840 45
rect 1860 25 1880 45
rect 1900 25 1920 45
rect 1940 25 1960 45
rect 1980 25 2000 45
rect 2020 25 2040 45
rect 2060 25 2080 45
rect 2100 25 2120 45
rect 2140 25 2160 45
rect 2180 25 2200 45
rect 2220 25 2240 45
rect 2260 25 2280 45
rect 2300 25 2320 45
rect 2340 25 2360 45
rect 2380 25 2400 45
rect 2420 25 2440 45
rect 2460 25 2480 45
rect 2500 25 2520 45
rect 2540 25 2560 45
rect 2580 25 2600 45
rect 2620 25 2640 45
rect 2660 25 2675 45
rect 175 15 2675 25
rect 1805 -35 1975 -20
rect 1805 -55 1820 -35
rect 1840 -55 1860 -35
rect 1880 -55 1900 -35
rect 1920 -55 1940 -35
rect 1960 -55 1975 -35
rect 1805 -70 1975 -55
rect 105 -225 2605 -215
rect 105 -245 120 -225
rect 140 -245 160 -225
rect 180 -245 200 -225
rect 220 -245 240 -225
rect 260 -245 280 -225
rect 300 -245 320 -225
rect 340 -245 360 -225
rect 380 -245 400 -225
rect 420 -245 440 -225
rect 460 -245 480 -225
rect 500 -245 520 -225
rect 540 -245 560 -225
rect 580 -245 600 -225
rect 620 -245 640 -225
rect 660 -245 680 -225
rect 700 -245 720 -225
rect 740 -245 760 -225
rect 780 -245 800 -225
rect 820 -245 840 -225
rect 860 -245 880 -225
rect 900 -245 920 -225
rect 940 -245 960 -225
rect 980 -245 1000 -225
rect 1020 -245 1040 -225
rect 1060 -245 1080 -225
rect 1100 -245 1120 -225
rect 1140 -245 1160 -225
rect 1180 -245 1200 -225
rect 1220 -245 1240 -225
rect 1260 -245 1280 -225
rect 1300 -245 1320 -225
rect 1340 -245 1360 -225
rect 1380 -245 1400 -225
rect 1420 -245 1440 -225
rect 1460 -245 1480 -225
rect 1500 -245 1520 -225
rect 1540 -245 1560 -225
rect 1580 -245 1600 -225
rect 1620 -245 1640 -225
rect 1660 -245 1680 -225
rect 1700 -245 1720 -225
rect 1740 -245 1760 -225
rect 1780 -245 1800 -225
rect 1820 -245 1840 -225
rect 1860 -245 1880 -225
rect 1900 -245 1920 -225
rect 1940 -245 1960 -225
rect 1980 -245 2000 -225
rect 2020 -245 2040 -225
rect 2060 -245 2080 -225
rect 2100 -245 2120 -225
rect 2140 -245 2160 -225
rect 2180 -245 2200 -225
rect 2220 -245 2240 -225
rect 2260 -245 2280 -225
rect 2300 -245 2320 -225
rect 2340 -245 2360 -225
rect 2380 -245 2400 -225
rect 2420 -245 2440 -225
rect 2460 -245 2480 -225
rect 2500 -245 2520 -225
rect 2540 -245 2560 -225
rect 2590 -245 2605 -225
rect 105 -265 2605 -245
rect 105 -285 120 -265
rect 140 -285 160 -265
rect 180 -285 200 -265
rect 220 -285 240 -265
rect 260 -285 280 -265
rect 300 -285 320 -265
rect 340 -285 360 -265
rect 380 -285 400 -265
rect 420 -285 440 -265
rect 460 -285 480 -265
rect 500 -285 520 -265
rect 540 -285 560 -265
rect 580 -285 600 -265
rect 620 -285 640 -265
rect 660 -285 680 -265
rect 700 -285 720 -265
rect 740 -285 760 -265
rect 780 -285 800 -265
rect 820 -285 840 -265
rect 860 -285 880 -265
rect 900 -285 920 -265
rect 940 -285 960 -265
rect 980 -285 1000 -265
rect 1020 -285 1040 -265
rect 1060 -285 1080 -265
rect 1100 -285 1120 -265
rect 1140 -285 1160 -265
rect 1180 -285 1200 -265
rect 1220 -285 1240 -265
rect 1260 -285 1280 -265
rect 1300 -285 1320 -265
rect 1340 -285 1360 -265
rect 1380 -285 1400 -265
rect 1420 -285 1440 -265
rect 1460 -285 1480 -265
rect 1500 -285 1520 -265
rect 1540 -285 1560 -265
rect 1580 -285 1600 -265
rect 1620 -285 1640 -265
rect 1660 -285 1680 -265
rect 1700 -285 1720 -265
rect 1740 -285 1760 -265
rect 1780 -285 1800 -265
rect 1820 -285 1840 -265
rect 1860 -285 1880 -265
rect 1900 -285 1920 -265
rect 1940 -285 1960 -265
rect 1980 -285 2000 -265
rect 2020 -285 2040 -265
rect 2060 -285 2080 -265
rect 2100 -285 2120 -265
rect 2140 -285 2160 -265
rect 2180 -285 2200 -265
rect 2220 -285 2240 -265
rect 2260 -285 2280 -265
rect 2300 -285 2320 -265
rect 2340 -285 2360 -265
rect 2380 -285 2400 -265
rect 2420 -285 2440 -265
rect 2460 -285 2480 -265
rect 2500 -285 2520 -265
rect 2540 -285 2560 -265
rect 2590 -285 2605 -265
rect 105 -295 2605 -285
rect -70 -310 85 -300
rect -70 -335 -60 -310
rect -40 -335 -20 -310
rect 0 -335 20 -310
rect 40 -335 60 -310
rect -70 -345 85 -335
rect 105 -360 2605 -350
rect 105 -380 120 -360
rect 140 -380 160 -360
rect 180 -380 200 -360
rect 220 -380 240 -360
rect 260 -380 280 -360
rect 300 -380 320 -360
rect 340 -380 360 -360
rect 380 -380 400 -360
rect 420 -380 440 -360
rect 460 -380 480 -360
rect 500 -380 520 -360
rect 540 -380 560 -360
rect 580 -380 600 -360
rect 620 -380 640 -360
rect 660 -380 680 -360
rect 700 -380 720 -360
rect 740 -380 760 -360
rect 780 -380 800 -360
rect 820 -380 840 -360
rect 860 -380 880 -360
rect 900 -380 920 -360
rect 940 -380 960 -360
rect 980 -380 1000 -360
rect 1020 -380 1040 -360
rect 1060 -380 1080 -360
rect 1100 -380 1120 -360
rect 1140 -380 1160 -360
rect 1180 -380 1200 -360
rect 1220 -380 1240 -360
rect 1260 -380 1280 -360
rect 1300 -380 1320 -360
rect 1340 -380 1360 -360
rect 1380 -380 1400 -360
rect 1420 -380 1440 -360
rect 1460 -380 1480 -360
rect 1500 -380 1520 -360
rect 1540 -380 1560 -360
rect 1580 -380 1600 -360
rect 1620 -380 1640 -360
rect 1660 -380 1680 -360
rect 1700 -380 1720 -360
rect 1740 -380 1760 -360
rect 1780 -380 1800 -360
rect 1820 -380 1840 -360
rect 1860 -380 1880 -360
rect 1900 -380 1920 -360
rect 1940 -380 1960 -360
rect 1980 -380 2000 -360
rect 2020 -380 2040 -360
rect 2060 -380 2080 -360
rect 2100 -380 2120 -360
rect 2140 -380 2160 -360
rect 2180 -380 2200 -360
rect 2220 -380 2240 -360
rect 2260 -380 2280 -360
rect 2300 -380 2320 -360
rect 2340 -380 2360 -360
rect 2380 -380 2400 -360
rect 2420 -380 2440 -360
rect 2460 -380 2480 -360
rect 2500 -380 2520 -360
rect 2540 -380 2560 -360
rect 2590 -380 2605 -360
rect 105 -390 2605 -380
rect -70 -405 85 -395
rect -70 -430 -60 -405
rect -40 -430 -20 -405
rect 0 -430 20 -405
rect 40 -430 60 -405
rect -70 -440 85 -430
rect 105 -455 2605 -445
rect 105 -475 120 -455
rect 140 -475 160 -455
rect 180 -475 200 -455
rect 220 -475 240 -455
rect 260 -475 280 -455
rect 300 -475 320 -455
rect 340 -475 360 -455
rect 380 -475 400 -455
rect 420 -475 440 -455
rect 460 -475 480 -455
rect 500 -475 520 -455
rect 540 -475 560 -455
rect 580 -475 600 -455
rect 620 -475 640 -455
rect 660 -475 680 -455
rect 700 -475 720 -455
rect 740 -475 760 -455
rect 780 -475 800 -455
rect 820 -475 840 -455
rect 860 -475 880 -455
rect 900 -475 920 -455
rect 940 -475 960 -455
rect 980 -475 1000 -455
rect 1020 -475 1040 -455
rect 1060 -475 1080 -455
rect 1100 -475 1120 -455
rect 1140 -475 1160 -455
rect 1180 -475 1200 -455
rect 1220 -475 1240 -455
rect 1260 -475 1280 -455
rect 1300 -475 1320 -455
rect 1340 -475 1360 -455
rect 1380 -475 1400 -455
rect 1420 -475 1440 -455
rect 1460 -475 1480 -455
rect 1500 -475 1520 -455
rect 1540 -475 1560 -455
rect 1580 -475 1600 -455
rect 1620 -475 1640 -455
rect 1660 -475 1680 -455
rect 1700 -475 1720 -455
rect 1740 -475 1760 -455
rect 1780 -475 1800 -455
rect 1820 -475 1840 -455
rect 1860 -475 1880 -455
rect 1900 -475 1920 -455
rect 1940 -475 1960 -455
rect 1980 -475 2000 -455
rect 2020 -475 2040 -455
rect 2060 -475 2080 -455
rect 2100 -475 2120 -455
rect 2140 -475 2160 -455
rect 2180 -475 2200 -455
rect 2220 -475 2240 -455
rect 2260 -475 2280 -455
rect 2300 -475 2320 -455
rect 2340 -475 2360 -455
rect 2380 -475 2400 -455
rect 2420 -475 2440 -455
rect 2460 -475 2480 -455
rect 2500 -475 2520 -455
rect 2540 -475 2560 -455
rect 2590 -475 2605 -455
rect 105 -485 2605 -475
rect -70 -500 85 -490
rect -70 -525 -60 -500
rect -40 -525 -20 -500
rect 0 -525 20 -500
rect 40 -525 60 -500
rect -70 -535 85 -525
rect 105 -550 2605 -540
rect 105 -570 120 -550
rect 140 -570 160 -550
rect 180 -570 200 -550
rect 220 -570 240 -550
rect 260 -570 280 -550
rect 300 -570 320 -550
rect 340 -570 360 -550
rect 380 -570 400 -550
rect 420 -570 440 -550
rect 460 -570 480 -550
rect 500 -570 520 -550
rect 540 -570 560 -550
rect 580 -570 600 -550
rect 620 -570 640 -550
rect 660 -570 680 -550
rect 700 -570 720 -550
rect 740 -570 760 -550
rect 780 -570 800 -550
rect 820 -570 840 -550
rect 860 -570 880 -550
rect 900 -570 920 -550
rect 940 -570 960 -550
rect 980 -570 1000 -550
rect 1020 -570 1040 -550
rect 1060 -570 1080 -550
rect 1100 -570 1120 -550
rect 1140 -570 1160 -550
rect 1180 -570 1200 -550
rect 1220 -570 1240 -550
rect 1260 -570 1280 -550
rect 1300 -570 1320 -550
rect 1340 -570 1360 -550
rect 1380 -570 1400 -550
rect 1420 -570 1440 -550
rect 1460 -570 1480 -550
rect 1500 -570 1520 -550
rect 1540 -570 1560 -550
rect 1580 -570 1600 -550
rect 1620 -570 1640 -550
rect 1660 -570 1680 -550
rect 1700 -570 1720 -550
rect 1740 -570 1760 -550
rect 1780 -570 1800 -550
rect 1820 -570 1840 -550
rect 1860 -570 1880 -550
rect 1900 -570 1920 -550
rect 1940 -570 1960 -550
rect 1980 -570 2000 -550
rect 2020 -570 2040 -550
rect 2060 -570 2080 -550
rect 2100 -570 2120 -550
rect 2140 -570 2160 -550
rect 2180 -570 2200 -550
rect 2220 -570 2240 -550
rect 2260 -570 2280 -550
rect 2300 -570 2320 -550
rect 2340 -570 2360 -550
rect 2380 -570 2400 -550
rect 2420 -570 2440 -550
rect 2460 -570 2480 -550
rect 2500 -570 2520 -550
rect 2540 -570 2560 -550
rect 2590 -570 2605 -550
rect 105 -580 2605 -570
rect -70 -595 85 -585
rect -70 -620 -60 -595
rect -40 -620 -20 -595
rect 0 -620 20 -595
rect 40 -620 60 -595
rect -70 -630 85 -620
rect 105 -645 2605 -635
rect 105 -665 120 -645
rect 140 -665 160 -645
rect 180 -665 200 -645
rect 220 -665 240 -645
rect 260 -665 280 -645
rect 300 -665 320 -645
rect 340 -665 360 -645
rect 380 -665 400 -645
rect 420 -665 440 -645
rect 460 -665 480 -645
rect 500 -665 520 -645
rect 540 -665 560 -645
rect 580 -665 600 -645
rect 620 -665 640 -645
rect 660 -665 680 -645
rect 700 -665 720 -645
rect 740 -665 760 -645
rect 780 -665 800 -645
rect 820 -665 840 -645
rect 860 -665 880 -645
rect 900 -665 920 -645
rect 940 -665 960 -645
rect 980 -665 1000 -645
rect 1020 -665 1040 -645
rect 1060 -665 1080 -645
rect 1100 -665 1120 -645
rect 1140 -665 1160 -645
rect 1180 -665 1200 -645
rect 1220 -665 1240 -645
rect 1260 -665 1280 -645
rect 1300 -665 1320 -645
rect 1340 -665 1360 -645
rect 1380 -665 1400 -645
rect 1420 -665 1440 -645
rect 1460 -665 1480 -645
rect 1500 -665 1520 -645
rect 1540 -665 1560 -645
rect 1580 -665 1600 -645
rect 1620 -665 1640 -645
rect 1660 -665 1680 -645
rect 1700 -665 1720 -645
rect 1740 -665 1760 -645
rect 1780 -665 1800 -645
rect 1820 -665 1840 -645
rect 1860 -665 1880 -645
rect 1900 -665 1920 -645
rect 1940 -665 1960 -645
rect 1980 -665 2000 -645
rect 2020 -665 2040 -645
rect 2060 -665 2080 -645
rect 2100 -665 2120 -645
rect 2140 -665 2160 -645
rect 2180 -665 2200 -645
rect 2220 -665 2240 -645
rect 2260 -665 2280 -645
rect 2300 -665 2320 -645
rect 2340 -665 2360 -645
rect 2380 -665 2400 -645
rect 2420 -665 2440 -645
rect 2460 -665 2480 -645
rect 2500 -665 2520 -645
rect 2540 -665 2560 -645
rect 2590 -665 2605 -645
rect 105 -675 2605 -665
rect -70 -690 85 -680
rect -70 -715 -60 -690
rect -40 -715 -20 -690
rect 0 -715 20 -690
rect 40 -715 60 -690
rect -70 -725 85 -715
rect 105 -740 2605 -730
rect 105 -760 120 -740
rect 140 -760 160 -740
rect 180 -760 200 -740
rect 220 -760 240 -740
rect 260 -760 280 -740
rect 300 -760 320 -740
rect 340 -760 360 -740
rect 380 -760 400 -740
rect 420 -760 440 -740
rect 460 -760 480 -740
rect 500 -760 520 -740
rect 540 -760 560 -740
rect 580 -760 600 -740
rect 620 -760 640 -740
rect 660 -760 680 -740
rect 700 -760 720 -740
rect 740 -760 760 -740
rect 780 -760 800 -740
rect 820 -760 840 -740
rect 860 -760 880 -740
rect 900 -760 920 -740
rect 940 -760 960 -740
rect 980 -760 1000 -740
rect 1020 -760 1040 -740
rect 1060 -760 1080 -740
rect 1100 -760 1120 -740
rect 1140 -760 1160 -740
rect 1180 -760 1200 -740
rect 1220 -760 1240 -740
rect 1260 -760 1280 -740
rect 1300 -760 1320 -740
rect 1340 -760 1360 -740
rect 1380 -760 1400 -740
rect 1420 -760 1440 -740
rect 1460 -760 1480 -740
rect 1500 -760 1520 -740
rect 1540 -760 1560 -740
rect 1580 -760 1600 -740
rect 1620 -760 1640 -740
rect 1660 -760 1680 -740
rect 1700 -760 1720 -740
rect 1740 -760 1760 -740
rect 1780 -760 1800 -740
rect 1820 -760 1840 -740
rect 1860 -760 1880 -740
rect 1900 -760 1920 -740
rect 1940 -760 1960 -740
rect 1980 -760 2000 -740
rect 2020 -760 2040 -740
rect 2060 -760 2080 -740
rect 2100 -760 2120 -740
rect 2140 -760 2160 -740
rect 2180 -760 2200 -740
rect 2220 -760 2240 -740
rect 2260 -760 2280 -740
rect 2300 -760 2320 -740
rect 2340 -760 2360 -740
rect 2380 -760 2400 -740
rect 2420 -760 2440 -740
rect 2460 -760 2480 -740
rect 2500 -760 2520 -740
rect 2540 -760 2560 -740
rect 2590 -760 2605 -740
rect 105 -770 2605 -760
rect -70 -785 85 -775
rect -70 -810 -60 -785
rect -40 -810 -20 -785
rect 0 -810 20 -785
rect 40 -810 60 -785
rect -70 -820 85 -810
rect 105 -835 2605 -825
rect 105 -855 120 -835
rect 140 -855 160 -835
rect 180 -855 200 -835
rect 220 -855 240 -835
rect 260 -855 280 -835
rect 300 -855 320 -835
rect 340 -855 360 -835
rect 380 -855 400 -835
rect 420 -855 440 -835
rect 460 -855 480 -835
rect 500 -855 520 -835
rect 540 -855 560 -835
rect 580 -855 600 -835
rect 620 -855 640 -835
rect 660 -855 680 -835
rect 700 -855 720 -835
rect 740 -855 760 -835
rect 780 -855 800 -835
rect 820 -855 840 -835
rect 860 -855 880 -835
rect 900 -855 920 -835
rect 940 -855 960 -835
rect 980 -855 1000 -835
rect 1020 -855 1040 -835
rect 1060 -855 1080 -835
rect 1100 -855 1120 -835
rect 1140 -855 1160 -835
rect 1180 -855 1200 -835
rect 1220 -855 1240 -835
rect 1260 -855 1280 -835
rect 1300 -855 1320 -835
rect 1340 -855 1360 -835
rect 1380 -855 1400 -835
rect 1420 -855 1440 -835
rect 1460 -855 1480 -835
rect 1500 -855 1520 -835
rect 1540 -855 1560 -835
rect 1580 -855 1600 -835
rect 1620 -855 1640 -835
rect 1660 -855 1680 -835
rect 1700 -855 1720 -835
rect 1740 -855 1760 -835
rect 1780 -855 1800 -835
rect 1820 -855 1840 -835
rect 1860 -855 1880 -835
rect 1900 -855 1920 -835
rect 1940 -855 1960 -835
rect 1980 -855 2000 -835
rect 2020 -855 2040 -835
rect 2060 -855 2080 -835
rect 2100 -855 2120 -835
rect 2140 -855 2160 -835
rect 2180 -855 2200 -835
rect 2220 -855 2240 -835
rect 2260 -855 2280 -835
rect 2300 -855 2320 -835
rect 2340 -855 2360 -835
rect 2380 -855 2400 -835
rect 2420 -855 2440 -835
rect 2460 -855 2480 -835
rect 2500 -855 2520 -835
rect 2540 -855 2560 -835
rect 2590 -855 2605 -835
rect 105 -865 2605 -855
rect -70 -880 85 -870
rect -70 -905 -60 -880
rect -40 -905 -20 -880
rect 0 -905 20 -880
rect 40 -905 60 -880
rect -70 -915 85 -905
rect 105 -930 2605 -920
rect 105 -950 120 -930
rect 140 -950 160 -930
rect 180 -950 200 -930
rect 220 -950 240 -930
rect 260 -950 280 -930
rect 300 -950 320 -930
rect 340 -950 360 -930
rect 380 -950 400 -930
rect 420 -950 440 -930
rect 460 -950 480 -930
rect 500 -950 520 -930
rect 540 -950 560 -930
rect 580 -950 600 -930
rect 620 -950 640 -930
rect 660 -950 680 -930
rect 700 -950 720 -930
rect 740 -950 760 -930
rect 780 -950 800 -930
rect 820 -950 840 -930
rect 860 -950 880 -930
rect 900 -950 920 -930
rect 940 -950 960 -930
rect 980 -950 1000 -930
rect 1020 -950 1040 -930
rect 1060 -950 1080 -930
rect 1100 -950 1120 -930
rect 1140 -950 1160 -930
rect 1180 -950 1200 -930
rect 1220 -950 1240 -930
rect 1260 -950 1280 -930
rect 1300 -950 1320 -930
rect 1340 -950 1360 -930
rect 1380 -950 1400 -930
rect 1420 -950 1440 -930
rect 1460 -950 1480 -930
rect 1500 -950 1520 -930
rect 1540 -950 1560 -930
rect 1580 -950 1600 -930
rect 1620 -950 1640 -930
rect 1660 -950 1680 -930
rect 1700 -950 1720 -930
rect 1740 -950 1760 -930
rect 1780 -950 1800 -930
rect 1820 -950 1840 -930
rect 1860 -950 1880 -930
rect 1900 -950 1920 -930
rect 1940 -950 1960 -930
rect 1980 -950 2000 -930
rect 2020 -950 2040 -930
rect 2060 -950 2080 -930
rect 2100 -950 2120 -930
rect 2140 -950 2160 -930
rect 2180 -950 2200 -930
rect 2220 -950 2240 -930
rect 2260 -950 2280 -930
rect 2300 -950 2320 -930
rect 2340 -950 2360 -930
rect 2380 -950 2400 -930
rect 2420 -950 2440 -930
rect 2460 -950 2480 -930
rect 2500 -950 2520 -930
rect 2540 -950 2560 -930
rect 2590 -950 2605 -930
rect 105 -960 2605 -950
rect -70 -975 85 -965
rect -70 -1000 -60 -975
rect -40 -1000 -20 -975
rect 0 -1000 20 -975
rect 40 -1000 60 -975
rect -70 -1010 85 -1000
rect 105 -1025 2605 -1015
rect 105 -1045 120 -1025
rect 140 -1045 160 -1025
rect 180 -1045 200 -1025
rect 220 -1045 240 -1025
rect 260 -1045 280 -1025
rect 300 -1045 320 -1025
rect 340 -1045 360 -1025
rect 380 -1045 400 -1025
rect 420 -1045 440 -1025
rect 460 -1045 480 -1025
rect 500 -1045 520 -1025
rect 540 -1045 560 -1025
rect 580 -1045 600 -1025
rect 620 -1045 640 -1025
rect 660 -1045 680 -1025
rect 700 -1045 720 -1025
rect 740 -1045 760 -1025
rect 780 -1045 800 -1025
rect 820 -1045 840 -1025
rect 860 -1045 880 -1025
rect 900 -1045 920 -1025
rect 940 -1045 960 -1025
rect 980 -1045 1000 -1025
rect 1020 -1045 1040 -1025
rect 1060 -1045 1080 -1025
rect 1100 -1045 1120 -1025
rect 1140 -1045 1160 -1025
rect 1180 -1045 1200 -1025
rect 1220 -1045 1240 -1025
rect 1260 -1045 1280 -1025
rect 1300 -1045 1320 -1025
rect 1340 -1045 1360 -1025
rect 1380 -1045 1400 -1025
rect 1420 -1045 1440 -1025
rect 1460 -1045 1480 -1025
rect 1500 -1045 1520 -1025
rect 1540 -1045 1560 -1025
rect 1580 -1045 1600 -1025
rect 1620 -1045 1640 -1025
rect 1660 -1045 1680 -1025
rect 1700 -1045 1720 -1025
rect 1740 -1045 1760 -1025
rect 1780 -1045 1800 -1025
rect 1820 -1045 1840 -1025
rect 1860 -1045 1880 -1025
rect 1900 -1045 1920 -1025
rect 1940 -1045 1960 -1025
rect 1980 -1045 2000 -1025
rect 2020 -1045 2040 -1025
rect 2060 -1045 2080 -1025
rect 2100 -1045 2120 -1025
rect 2140 -1045 2160 -1025
rect 2180 -1045 2200 -1025
rect 2220 -1045 2240 -1025
rect 2260 -1045 2280 -1025
rect 2300 -1045 2320 -1025
rect 2340 -1045 2360 -1025
rect 2380 -1045 2400 -1025
rect 2420 -1045 2440 -1025
rect 2460 -1045 2480 -1025
rect 2500 -1045 2520 -1025
rect 2540 -1045 2560 -1025
rect 2590 -1045 2605 -1025
rect 105 -1055 2605 -1045
rect -70 -1070 85 -1060
rect -70 -1095 -60 -1070
rect -40 -1095 -20 -1070
rect 0 -1095 20 -1070
rect 40 -1095 60 -1070
rect -70 -1105 85 -1095
rect 105 -1120 2605 -1110
rect 105 -1140 120 -1120
rect 140 -1140 160 -1120
rect 180 -1140 200 -1120
rect 220 -1140 240 -1120
rect 260 -1140 280 -1120
rect 300 -1140 320 -1120
rect 340 -1140 360 -1120
rect 380 -1140 400 -1120
rect 420 -1140 440 -1120
rect 460 -1140 480 -1120
rect 500 -1140 520 -1120
rect 540 -1140 560 -1120
rect 580 -1140 600 -1120
rect 620 -1140 640 -1120
rect 660 -1140 680 -1120
rect 700 -1140 720 -1120
rect 740 -1140 760 -1120
rect 780 -1140 800 -1120
rect 820 -1140 840 -1120
rect 860 -1140 880 -1120
rect 900 -1140 920 -1120
rect 940 -1140 960 -1120
rect 980 -1140 1000 -1120
rect 1020 -1140 1040 -1120
rect 1060 -1140 1080 -1120
rect 1100 -1140 1120 -1120
rect 1140 -1140 1160 -1120
rect 1180 -1140 1200 -1120
rect 1220 -1140 1240 -1120
rect 1260 -1140 1280 -1120
rect 1300 -1140 1320 -1120
rect 1340 -1140 1360 -1120
rect 1380 -1140 1400 -1120
rect 1420 -1140 1440 -1120
rect 1460 -1140 1480 -1120
rect 1500 -1140 1520 -1120
rect 1540 -1140 1560 -1120
rect 1580 -1140 1600 -1120
rect 1620 -1140 1640 -1120
rect 1660 -1140 1680 -1120
rect 1700 -1140 1720 -1120
rect 1740 -1140 1760 -1120
rect 1780 -1140 1800 -1120
rect 1820 -1140 1840 -1120
rect 1860 -1140 1880 -1120
rect 1900 -1140 1920 -1120
rect 1940 -1140 1960 -1120
rect 1980 -1140 2000 -1120
rect 2020 -1140 2040 -1120
rect 2060 -1140 2080 -1120
rect 2100 -1140 2120 -1120
rect 2140 -1140 2160 -1120
rect 2180 -1140 2200 -1120
rect 2220 -1140 2240 -1120
rect 2260 -1140 2280 -1120
rect 2300 -1140 2320 -1120
rect 2340 -1140 2360 -1120
rect 2380 -1140 2400 -1120
rect 2420 -1140 2440 -1120
rect 2460 -1140 2480 -1120
rect 2500 -1140 2520 -1120
rect 2540 -1140 2560 -1120
rect 2590 -1140 2605 -1120
rect 105 -1150 2605 -1140
rect -70 -1165 85 -1155
rect -70 -1190 -60 -1165
rect -40 -1190 -20 -1165
rect 0 -1190 20 -1165
rect 40 -1190 60 -1165
rect -70 -1200 85 -1190
rect 105 -1215 2605 -1205
rect 105 -1235 120 -1215
rect 140 -1235 160 -1215
rect 180 -1235 200 -1215
rect 220 -1235 240 -1215
rect 260 -1235 280 -1215
rect 300 -1235 320 -1215
rect 340 -1235 360 -1215
rect 380 -1235 400 -1215
rect 420 -1235 440 -1215
rect 460 -1235 480 -1215
rect 500 -1235 520 -1215
rect 540 -1235 560 -1215
rect 580 -1235 600 -1215
rect 620 -1235 640 -1215
rect 660 -1235 680 -1215
rect 700 -1235 720 -1215
rect 740 -1235 760 -1215
rect 780 -1235 800 -1215
rect 820 -1235 840 -1215
rect 860 -1235 880 -1215
rect 900 -1235 920 -1215
rect 940 -1235 960 -1215
rect 980 -1235 1000 -1215
rect 1020 -1235 1040 -1215
rect 1060 -1235 1080 -1215
rect 1100 -1235 1120 -1215
rect 1140 -1235 1160 -1215
rect 1180 -1235 1200 -1215
rect 1220 -1235 1240 -1215
rect 1260 -1235 1280 -1215
rect 1300 -1235 1320 -1215
rect 1340 -1235 1360 -1215
rect 1380 -1235 1400 -1215
rect 1420 -1235 1440 -1215
rect 1460 -1235 1480 -1215
rect 1500 -1235 1520 -1215
rect 1540 -1235 1560 -1215
rect 1580 -1235 1600 -1215
rect 1620 -1235 1640 -1215
rect 1660 -1235 1680 -1215
rect 1700 -1235 1720 -1215
rect 1740 -1235 1760 -1215
rect 1780 -1235 1800 -1215
rect 1820 -1235 1840 -1215
rect 1860 -1235 1880 -1215
rect 1900 -1235 1920 -1215
rect 1940 -1235 1960 -1215
rect 1980 -1235 2000 -1215
rect 2020 -1235 2040 -1215
rect 2060 -1235 2080 -1215
rect 2100 -1235 2120 -1215
rect 2140 -1235 2160 -1215
rect 2180 -1235 2200 -1215
rect 2220 -1235 2240 -1215
rect 2260 -1235 2280 -1215
rect 2300 -1235 2320 -1215
rect 2340 -1235 2360 -1215
rect 2380 -1235 2400 -1215
rect 2420 -1235 2440 -1215
rect 2460 -1235 2480 -1215
rect 2500 -1235 2520 -1215
rect 2540 -1235 2560 -1215
rect 2590 -1235 2605 -1215
rect 105 -1245 2605 -1235
rect -70 -1260 85 -1250
rect -70 -1285 -60 -1260
rect -40 -1285 -20 -1260
rect 0 -1285 20 -1260
rect 40 -1285 60 -1260
rect -70 -1295 85 -1285
rect 105 -1310 2605 -1300
rect 105 -1330 120 -1310
rect 140 -1330 160 -1310
rect 180 -1330 200 -1310
rect 220 -1330 240 -1310
rect 260 -1330 280 -1310
rect 300 -1330 320 -1310
rect 340 -1330 360 -1310
rect 380 -1330 400 -1310
rect 420 -1330 440 -1310
rect 460 -1330 480 -1310
rect 500 -1330 520 -1310
rect 540 -1330 560 -1310
rect 580 -1330 600 -1310
rect 620 -1330 640 -1310
rect 660 -1330 680 -1310
rect 700 -1330 720 -1310
rect 740 -1330 760 -1310
rect 780 -1330 800 -1310
rect 820 -1330 840 -1310
rect 860 -1330 880 -1310
rect 900 -1330 920 -1310
rect 940 -1330 960 -1310
rect 980 -1330 1000 -1310
rect 1020 -1330 1040 -1310
rect 1060 -1330 1080 -1310
rect 1100 -1330 1120 -1310
rect 1140 -1330 1160 -1310
rect 1180 -1330 1200 -1310
rect 1220 -1330 1240 -1310
rect 1260 -1330 1280 -1310
rect 1300 -1330 1320 -1310
rect 1340 -1330 1360 -1310
rect 1380 -1330 1400 -1310
rect 1420 -1330 1440 -1310
rect 1460 -1330 1480 -1310
rect 1500 -1330 1520 -1310
rect 1540 -1330 1560 -1310
rect 1580 -1330 1600 -1310
rect 1620 -1330 1640 -1310
rect 1660 -1330 1680 -1310
rect 1700 -1330 1720 -1310
rect 1740 -1330 1760 -1310
rect 1780 -1330 1800 -1310
rect 1820 -1330 1840 -1310
rect 1860 -1330 1880 -1310
rect 1900 -1330 1920 -1310
rect 1940 -1330 1960 -1310
rect 1980 -1330 2000 -1310
rect 2020 -1330 2040 -1310
rect 2060 -1330 2080 -1310
rect 2100 -1330 2120 -1310
rect 2140 -1330 2160 -1310
rect 2180 -1330 2200 -1310
rect 2220 -1330 2240 -1310
rect 2260 -1330 2280 -1310
rect 2300 -1330 2320 -1310
rect 2340 -1330 2360 -1310
rect 2380 -1330 2400 -1310
rect 2420 -1330 2440 -1310
rect 2460 -1330 2480 -1310
rect 2500 -1330 2520 -1310
rect 2540 -1330 2560 -1310
rect 2590 -1330 2605 -1310
rect 105 -1340 2605 -1330
rect -70 -1355 85 -1345
rect -70 -1380 -60 -1355
rect -40 -1380 -20 -1355
rect 0 -1380 20 -1355
rect 40 -1380 60 -1355
rect -70 -1390 85 -1380
rect 105 -1405 2605 -1395
rect 105 -1425 120 -1405
rect 140 -1425 160 -1405
rect 180 -1425 200 -1405
rect 220 -1425 240 -1405
rect 260 -1425 280 -1405
rect 300 -1425 320 -1405
rect 340 -1425 360 -1405
rect 380 -1425 400 -1405
rect 420 -1425 440 -1405
rect 460 -1425 480 -1405
rect 500 -1425 520 -1405
rect 540 -1425 560 -1405
rect 580 -1425 600 -1405
rect 620 -1425 640 -1405
rect 660 -1425 680 -1405
rect 700 -1425 720 -1405
rect 740 -1425 760 -1405
rect 780 -1425 800 -1405
rect 820 -1425 840 -1405
rect 860 -1425 880 -1405
rect 900 -1425 920 -1405
rect 940 -1425 960 -1405
rect 980 -1425 1000 -1405
rect 1020 -1425 1040 -1405
rect 1060 -1425 1080 -1405
rect 1100 -1425 1120 -1405
rect 1140 -1425 1160 -1405
rect 1180 -1425 1200 -1405
rect 1220 -1425 1240 -1405
rect 1260 -1425 1280 -1405
rect 1300 -1425 1320 -1405
rect 1340 -1425 1360 -1405
rect 1380 -1425 1400 -1405
rect 1420 -1425 1440 -1405
rect 1460 -1425 1480 -1405
rect 1500 -1425 1520 -1405
rect 1540 -1425 1560 -1405
rect 1580 -1425 1600 -1405
rect 1620 -1425 1640 -1405
rect 1660 -1425 1680 -1405
rect 1700 -1425 1720 -1405
rect 1740 -1425 1760 -1405
rect 1780 -1425 1800 -1405
rect 1820 -1425 1840 -1405
rect 1860 -1425 1880 -1405
rect 1900 -1425 1920 -1405
rect 1940 -1425 1960 -1405
rect 1980 -1425 2000 -1405
rect 2020 -1425 2040 -1405
rect 2060 -1425 2080 -1405
rect 2100 -1425 2120 -1405
rect 2140 -1425 2160 -1405
rect 2180 -1425 2200 -1405
rect 2220 -1425 2240 -1405
rect 2260 -1425 2280 -1405
rect 2300 -1425 2320 -1405
rect 2340 -1425 2360 -1405
rect 2380 -1425 2400 -1405
rect 2420 -1425 2440 -1405
rect 2460 -1425 2480 -1405
rect 2500 -1425 2520 -1405
rect 2540 -1425 2560 -1405
rect 2590 -1425 2605 -1405
rect 105 -1435 2605 -1425
rect -70 -1450 85 -1440
rect -70 -1475 -60 -1450
rect -40 -1475 -20 -1450
rect 0 -1475 20 -1450
rect 40 -1475 60 -1450
rect -70 -1485 85 -1475
rect 105 -1500 2605 -1490
rect 105 -1520 120 -1500
rect 140 -1520 160 -1500
rect 180 -1520 200 -1500
rect 220 -1520 240 -1500
rect 260 -1520 280 -1500
rect 300 -1520 320 -1500
rect 340 -1520 360 -1500
rect 380 -1520 400 -1500
rect 420 -1520 440 -1500
rect 460 -1520 480 -1500
rect 500 -1520 520 -1500
rect 540 -1520 560 -1500
rect 580 -1520 600 -1500
rect 620 -1520 640 -1500
rect 660 -1520 680 -1500
rect 700 -1520 720 -1500
rect 740 -1520 760 -1500
rect 780 -1520 800 -1500
rect 820 -1520 840 -1500
rect 860 -1520 880 -1500
rect 900 -1520 920 -1500
rect 940 -1520 960 -1500
rect 980 -1520 1000 -1500
rect 1020 -1520 1040 -1500
rect 1060 -1520 1080 -1500
rect 1100 -1520 1120 -1500
rect 1140 -1520 1160 -1500
rect 1180 -1520 1200 -1500
rect 1220 -1520 1240 -1500
rect 1260 -1520 1280 -1500
rect 1300 -1520 1320 -1500
rect 1340 -1520 1360 -1500
rect 1380 -1520 1400 -1500
rect 1420 -1520 1440 -1500
rect 1460 -1520 1480 -1500
rect 1500 -1520 1520 -1500
rect 1540 -1520 1560 -1500
rect 1580 -1520 1600 -1500
rect 1620 -1520 1640 -1500
rect 1660 -1520 1680 -1500
rect 1700 -1520 1720 -1500
rect 1740 -1520 1760 -1500
rect 1780 -1520 1800 -1500
rect 1820 -1520 1840 -1500
rect 1860 -1520 1880 -1500
rect 1900 -1520 1920 -1500
rect 1940 -1520 1960 -1500
rect 1980 -1520 2000 -1500
rect 2020 -1520 2040 -1500
rect 2060 -1520 2080 -1500
rect 2100 -1520 2120 -1500
rect 2140 -1520 2160 -1500
rect 2180 -1520 2200 -1500
rect 2220 -1520 2240 -1500
rect 2260 -1520 2280 -1500
rect 2300 -1520 2320 -1500
rect 2340 -1520 2360 -1500
rect 2380 -1520 2400 -1500
rect 2420 -1520 2440 -1500
rect 2460 -1520 2480 -1500
rect 2500 -1520 2520 -1500
rect 2540 -1520 2560 -1500
rect 2590 -1520 2605 -1500
rect 105 -1530 2605 -1520
rect -70 -1545 85 -1535
rect -70 -1570 -60 -1545
rect -40 -1570 -20 -1545
rect 0 -1570 20 -1545
rect 40 -1570 60 -1545
rect -70 -1580 85 -1570
rect 105 -1595 2605 -1585
rect 105 -1615 120 -1595
rect 140 -1615 160 -1595
rect 180 -1615 200 -1595
rect 220 -1615 240 -1595
rect 260 -1615 280 -1595
rect 300 -1615 320 -1595
rect 340 -1615 360 -1595
rect 380 -1615 400 -1595
rect 420 -1615 440 -1595
rect 460 -1615 480 -1595
rect 500 -1615 520 -1595
rect 540 -1615 560 -1595
rect 580 -1615 600 -1595
rect 620 -1615 640 -1595
rect 660 -1615 680 -1595
rect 700 -1615 720 -1595
rect 740 -1615 760 -1595
rect 780 -1615 800 -1595
rect 820 -1615 840 -1595
rect 860 -1615 880 -1595
rect 900 -1615 920 -1595
rect 940 -1615 960 -1595
rect 980 -1615 1000 -1595
rect 1020 -1615 1040 -1595
rect 1060 -1615 1080 -1595
rect 1100 -1615 1120 -1595
rect 1140 -1615 1160 -1595
rect 1180 -1615 1200 -1595
rect 1220 -1615 1240 -1595
rect 1260 -1615 1280 -1595
rect 1300 -1615 1320 -1595
rect 1340 -1615 1360 -1595
rect 1380 -1615 1400 -1595
rect 1420 -1615 1440 -1595
rect 1460 -1615 1480 -1595
rect 1500 -1615 1520 -1595
rect 1540 -1615 1560 -1595
rect 1580 -1615 1600 -1595
rect 1620 -1615 1640 -1595
rect 1660 -1615 1680 -1595
rect 1700 -1615 1720 -1595
rect 1740 -1615 1760 -1595
rect 1780 -1615 1800 -1595
rect 1820 -1615 1840 -1595
rect 1860 -1615 1880 -1595
rect 1900 -1615 1920 -1595
rect 1940 -1615 1960 -1595
rect 1980 -1615 2000 -1595
rect 2020 -1615 2040 -1595
rect 2060 -1615 2080 -1595
rect 2100 -1615 2120 -1595
rect 2140 -1615 2160 -1595
rect 2180 -1615 2200 -1595
rect 2220 -1615 2240 -1595
rect 2260 -1615 2280 -1595
rect 2300 -1615 2320 -1595
rect 2340 -1615 2360 -1595
rect 2380 -1615 2400 -1595
rect 2420 -1615 2440 -1595
rect 2460 -1615 2480 -1595
rect 2500 -1615 2520 -1595
rect 2540 -1615 2560 -1595
rect 2590 -1615 2605 -1595
rect 105 -1625 2605 -1615
rect -70 -1640 85 -1630
rect -70 -1665 -60 -1640
rect -40 -1665 -20 -1640
rect 0 -1665 20 -1640
rect 40 -1665 60 -1640
rect -70 -1675 85 -1665
rect 105 -1690 2605 -1680
rect 105 -1710 120 -1690
rect 140 -1710 160 -1690
rect 180 -1710 200 -1690
rect 220 -1710 240 -1690
rect 260 -1710 280 -1690
rect 300 -1710 320 -1690
rect 340 -1710 360 -1690
rect 380 -1710 400 -1690
rect 420 -1710 440 -1690
rect 460 -1710 480 -1690
rect 500 -1710 520 -1690
rect 540 -1710 560 -1690
rect 580 -1710 600 -1690
rect 620 -1710 640 -1690
rect 660 -1710 680 -1690
rect 700 -1710 720 -1690
rect 740 -1710 760 -1690
rect 780 -1710 800 -1690
rect 820 -1710 840 -1690
rect 860 -1710 880 -1690
rect 900 -1710 920 -1690
rect 940 -1710 960 -1690
rect 980 -1710 1000 -1690
rect 1020 -1710 1040 -1690
rect 1060 -1710 1080 -1690
rect 1100 -1710 1120 -1690
rect 1140 -1710 1160 -1690
rect 1180 -1710 1200 -1690
rect 1220 -1710 1240 -1690
rect 1260 -1710 1280 -1690
rect 1300 -1710 1320 -1690
rect 1340 -1710 1360 -1690
rect 1380 -1710 1400 -1690
rect 1420 -1710 1440 -1690
rect 1460 -1710 1480 -1690
rect 1500 -1710 1520 -1690
rect 1540 -1710 1560 -1690
rect 1580 -1710 1600 -1690
rect 1620 -1710 1640 -1690
rect 1660 -1710 1680 -1690
rect 1700 -1710 1720 -1690
rect 1740 -1710 1760 -1690
rect 1780 -1710 1800 -1690
rect 1820 -1710 1840 -1690
rect 1860 -1710 1880 -1690
rect 1900 -1710 1920 -1690
rect 1940 -1710 1960 -1690
rect 1980 -1710 2000 -1690
rect 2020 -1710 2040 -1690
rect 2060 -1710 2080 -1690
rect 2100 -1710 2120 -1690
rect 2140 -1710 2160 -1690
rect 2180 -1710 2200 -1690
rect 2220 -1710 2240 -1690
rect 2260 -1710 2280 -1690
rect 2300 -1710 2320 -1690
rect 2340 -1710 2360 -1690
rect 2380 -1710 2400 -1690
rect 2420 -1710 2440 -1690
rect 2460 -1710 2480 -1690
rect 2500 -1710 2520 -1690
rect 2540 -1710 2560 -1690
rect 2590 -1710 2605 -1690
rect 105 -1720 2605 -1710
rect -70 -1735 85 -1725
rect -70 -1760 -60 -1735
rect -40 -1760 -20 -1735
rect 0 -1760 20 -1735
rect 40 -1760 60 -1735
rect -70 -1770 85 -1760
rect 105 -1785 2605 -1775
rect 105 -1805 120 -1785
rect 140 -1805 160 -1785
rect 180 -1805 200 -1785
rect 220 -1805 240 -1785
rect 260 -1805 280 -1785
rect 300 -1805 320 -1785
rect 340 -1805 360 -1785
rect 380 -1805 400 -1785
rect 420 -1805 440 -1785
rect 460 -1805 480 -1785
rect 500 -1805 520 -1785
rect 540 -1805 560 -1785
rect 580 -1805 600 -1785
rect 620 -1805 640 -1785
rect 660 -1805 680 -1785
rect 700 -1805 720 -1785
rect 740 -1805 760 -1785
rect 780 -1805 800 -1785
rect 820 -1805 840 -1785
rect 860 -1805 880 -1785
rect 900 -1805 920 -1785
rect 940 -1805 960 -1785
rect 980 -1805 1000 -1785
rect 1020 -1805 1040 -1785
rect 1060 -1805 1080 -1785
rect 1100 -1805 1120 -1785
rect 1140 -1805 1160 -1785
rect 1180 -1805 1200 -1785
rect 1220 -1805 1240 -1785
rect 1260 -1805 1280 -1785
rect 1300 -1805 1320 -1785
rect 1340 -1805 1360 -1785
rect 1380 -1805 1400 -1785
rect 1420 -1805 1440 -1785
rect 1460 -1805 1480 -1785
rect 1500 -1805 1520 -1785
rect 1540 -1805 1560 -1785
rect 1580 -1805 1600 -1785
rect 1620 -1805 1640 -1785
rect 1660 -1805 1680 -1785
rect 1700 -1805 1720 -1785
rect 1740 -1805 1760 -1785
rect 1780 -1805 1800 -1785
rect 1820 -1805 1840 -1785
rect 1860 -1805 1880 -1785
rect 1900 -1805 1920 -1785
rect 1940 -1805 1960 -1785
rect 1980 -1805 2000 -1785
rect 2020 -1805 2040 -1785
rect 2060 -1805 2080 -1785
rect 2100 -1805 2120 -1785
rect 2140 -1805 2160 -1785
rect 2180 -1805 2200 -1785
rect 2220 -1805 2240 -1785
rect 2260 -1805 2280 -1785
rect 2300 -1805 2320 -1785
rect 2340 -1805 2360 -1785
rect 2380 -1805 2400 -1785
rect 2420 -1805 2440 -1785
rect 2460 -1805 2480 -1785
rect 2500 -1805 2520 -1785
rect 2540 -1805 2560 -1785
rect 2590 -1805 2605 -1785
rect 105 -1815 2605 -1805
rect -70 -1830 85 -1820
rect -70 -1855 -60 -1830
rect -40 -1855 -20 -1830
rect 0 -1855 20 -1830
rect 40 -1855 60 -1830
rect -70 -1865 85 -1855
rect 105 -1880 2605 -1870
rect 105 -1900 120 -1880
rect 140 -1900 160 -1880
rect 180 -1900 200 -1880
rect 220 -1900 240 -1880
rect 260 -1900 280 -1880
rect 300 -1900 320 -1880
rect 340 -1900 360 -1880
rect 380 -1900 400 -1880
rect 420 -1900 440 -1880
rect 460 -1900 480 -1880
rect 500 -1900 520 -1880
rect 540 -1900 560 -1880
rect 580 -1900 600 -1880
rect 620 -1900 640 -1880
rect 660 -1900 680 -1880
rect 700 -1900 720 -1880
rect 740 -1900 760 -1880
rect 780 -1900 800 -1880
rect 820 -1900 840 -1880
rect 860 -1900 880 -1880
rect 900 -1900 920 -1880
rect 940 -1900 960 -1880
rect 980 -1900 1000 -1880
rect 1020 -1900 1040 -1880
rect 1060 -1900 1080 -1880
rect 1100 -1900 1120 -1880
rect 1140 -1900 1160 -1880
rect 1180 -1900 1200 -1880
rect 1220 -1900 1240 -1880
rect 1260 -1900 1280 -1880
rect 1300 -1900 1320 -1880
rect 1340 -1900 1360 -1880
rect 1380 -1900 1400 -1880
rect 1420 -1900 1440 -1880
rect 1460 -1900 1480 -1880
rect 1500 -1900 1520 -1880
rect 1540 -1900 1560 -1880
rect 1580 -1900 1600 -1880
rect 1620 -1900 1640 -1880
rect 1660 -1900 1680 -1880
rect 1700 -1900 1720 -1880
rect 1740 -1900 1760 -1880
rect 1780 -1900 1800 -1880
rect 1820 -1900 1840 -1880
rect 1860 -1900 1880 -1880
rect 1900 -1900 1920 -1880
rect 1940 -1900 1960 -1880
rect 1980 -1900 2000 -1880
rect 2020 -1900 2040 -1880
rect 2060 -1900 2080 -1880
rect 2100 -1900 2120 -1880
rect 2140 -1900 2160 -1880
rect 2180 -1900 2200 -1880
rect 2220 -1900 2240 -1880
rect 2260 -1900 2280 -1880
rect 2300 -1900 2320 -1880
rect 2340 -1900 2360 -1880
rect 2380 -1900 2400 -1880
rect 2420 -1900 2440 -1880
rect 2460 -1900 2480 -1880
rect 2500 -1900 2520 -1880
rect 2540 -1900 2560 -1880
rect 2590 -1900 2605 -1880
rect 105 -1910 2605 -1900
rect -70 -1925 85 -1915
rect -70 -1950 -60 -1925
rect -40 -1950 -20 -1925
rect 0 -1950 20 -1925
rect 40 -1950 60 -1925
rect -70 -1960 85 -1950
rect 105 -1975 2605 -1965
rect 105 -1995 120 -1975
rect 140 -1995 160 -1975
rect 180 -1995 200 -1975
rect 220 -1995 240 -1975
rect 260 -1995 280 -1975
rect 300 -1995 320 -1975
rect 340 -1995 360 -1975
rect 380 -1995 400 -1975
rect 420 -1995 440 -1975
rect 460 -1995 480 -1975
rect 500 -1995 520 -1975
rect 540 -1995 560 -1975
rect 580 -1995 600 -1975
rect 620 -1995 640 -1975
rect 660 -1995 680 -1975
rect 700 -1995 720 -1975
rect 740 -1995 760 -1975
rect 780 -1995 800 -1975
rect 820 -1995 840 -1975
rect 860 -1995 880 -1975
rect 900 -1995 920 -1975
rect 940 -1995 960 -1975
rect 980 -1995 1000 -1975
rect 1020 -1995 1040 -1975
rect 1060 -1995 1080 -1975
rect 1100 -1995 1120 -1975
rect 1140 -1995 1160 -1975
rect 1180 -1995 1200 -1975
rect 1220 -1995 1240 -1975
rect 1260 -1995 1280 -1975
rect 1300 -1995 1320 -1975
rect 1340 -1995 1360 -1975
rect 1380 -1995 1400 -1975
rect 1420 -1995 1440 -1975
rect 1460 -1995 1480 -1975
rect 1500 -1995 1520 -1975
rect 1540 -1995 1560 -1975
rect 1580 -1995 1600 -1975
rect 1620 -1995 1640 -1975
rect 1660 -1995 1680 -1975
rect 1700 -1995 1720 -1975
rect 1740 -1995 1760 -1975
rect 1780 -1995 1800 -1975
rect 1820 -1995 1840 -1975
rect 1860 -1995 1880 -1975
rect 1900 -1995 1920 -1975
rect 1940 -1995 1960 -1975
rect 1980 -1995 2000 -1975
rect 2020 -1995 2040 -1975
rect 2060 -1995 2080 -1975
rect 2100 -1995 2120 -1975
rect 2140 -1995 2160 -1975
rect 2180 -1995 2200 -1975
rect 2220 -1995 2240 -1975
rect 2260 -1995 2280 -1975
rect 2300 -1995 2320 -1975
rect 2340 -1995 2360 -1975
rect 2380 -1995 2400 -1975
rect 2420 -1995 2440 -1975
rect 2460 -1995 2480 -1975
rect 2500 -1995 2520 -1975
rect 2540 -1995 2560 -1975
rect 2590 -1995 2605 -1975
rect 105 -2005 2605 -1995
rect -70 -2020 85 -2010
rect -70 -2045 -60 -2020
rect -40 -2045 -20 -2020
rect 0 -2045 20 -2020
rect 40 -2045 60 -2020
rect -70 -2055 85 -2045
rect 105 -2070 2605 -2060
rect 105 -2090 120 -2070
rect 140 -2090 160 -2070
rect 180 -2090 200 -2070
rect 220 -2090 240 -2070
rect 260 -2090 280 -2070
rect 300 -2090 320 -2070
rect 340 -2090 360 -2070
rect 380 -2090 400 -2070
rect 420 -2090 440 -2070
rect 460 -2090 480 -2070
rect 500 -2090 520 -2070
rect 540 -2090 560 -2070
rect 580 -2090 600 -2070
rect 620 -2090 640 -2070
rect 660 -2090 680 -2070
rect 700 -2090 720 -2070
rect 740 -2090 760 -2070
rect 780 -2090 800 -2070
rect 820 -2090 840 -2070
rect 860 -2090 880 -2070
rect 900 -2090 920 -2070
rect 940 -2090 960 -2070
rect 980 -2090 1000 -2070
rect 1020 -2090 1040 -2070
rect 1060 -2090 1080 -2070
rect 1100 -2090 1120 -2070
rect 1140 -2090 1160 -2070
rect 1180 -2090 1200 -2070
rect 1220 -2090 1240 -2070
rect 1260 -2090 1280 -2070
rect 1300 -2090 1320 -2070
rect 1340 -2090 1360 -2070
rect 1380 -2090 1400 -2070
rect 1420 -2090 1440 -2070
rect 1460 -2090 1480 -2070
rect 1500 -2090 1520 -2070
rect 1540 -2090 1560 -2070
rect 1580 -2090 1600 -2070
rect 1620 -2090 1640 -2070
rect 1660 -2090 1680 -2070
rect 1700 -2090 1720 -2070
rect 1740 -2090 1760 -2070
rect 1780 -2090 1800 -2070
rect 1820 -2090 1840 -2070
rect 1860 -2090 1880 -2070
rect 1900 -2090 1920 -2070
rect 1940 -2090 1960 -2070
rect 1980 -2090 2000 -2070
rect 2020 -2090 2040 -2070
rect 2060 -2090 2080 -2070
rect 2100 -2090 2120 -2070
rect 2140 -2090 2160 -2070
rect 2180 -2090 2200 -2070
rect 2220 -2090 2240 -2070
rect 2260 -2090 2280 -2070
rect 2300 -2090 2320 -2070
rect 2340 -2090 2360 -2070
rect 2380 -2090 2400 -2070
rect 2420 -2090 2440 -2070
rect 2460 -2090 2480 -2070
rect 2500 -2090 2520 -2070
rect 2540 -2090 2560 -2070
rect 2590 -2090 2605 -2070
rect 105 -2100 2605 -2090
rect -70 -2115 85 -2105
rect -70 -2140 -60 -2115
rect -40 -2140 -20 -2115
rect 0 -2140 20 -2115
rect 40 -2140 60 -2115
rect -70 -2150 85 -2140
rect 105 -2165 2605 -2155
rect 105 -2185 120 -2165
rect 140 -2185 160 -2165
rect 180 -2185 200 -2165
rect 220 -2185 240 -2165
rect 260 -2185 280 -2165
rect 300 -2185 320 -2165
rect 340 -2185 360 -2165
rect 380 -2185 400 -2165
rect 420 -2185 440 -2165
rect 460 -2185 480 -2165
rect 500 -2185 520 -2165
rect 540 -2185 560 -2165
rect 580 -2185 600 -2165
rect 620 -2185 640 -2165
rect 660 -2185 680 -2165
rect 700 -2185 720 -2165
rect 740 -2185 760 -2165
rect 780 -2185 800 -2165
rect 820 -2185 840 -2165
rect 860 -2185 880 -2165
rect 900 -2185 920 -2165
rect 940 -2185 960 -2165
rect 980 -2185 1000 -2165
rect 1020 -2185 1040 -2165
rect 1060 -2185 1080 -2165
rect 1100 -2185 1120 -2165
rect 1140 -2185 1160 -2165
rect 1180 -2185 1200 -2165
rect 1220 -2185 1240 -2165
rect 1260 -2185 1280 -2165
rect 1300 -2185 1320 -2165
rect 1340 -2185 1360 -2165
rect 1380 -2185 1400 -2165
rect 1420 -2185 1440 -2165
rect 1460 -2185 1480 -2165
rect 1500 -2185 1520 -2165
rect 1540 -2185 1560 -2165
rect 1580 -2185 1600 -2165
rect 1620 -2185 1640 -2165
rect 1660 -2185 1680 -2165
rect 1700 -2185 1720 -2165
rect 1740 -2185 1760 -2165
rect 1780 -2185 1800 -2165
rect 1820 -2185 1840 -2165
rect 1860 -2185 1880 -2165
rect 1900 -2185 1920 -2165
rect 1940 -2185 1960 -2165
rect 1980 -2185 2000 -2165
rect 2020 -2185 2040 -2165
rect 2060 -2185 2080 -2165
rect 2100 -2185 2120 -2165
rect 2140 -2185 2160 -2165
rect 2180 -2185 2200 -2165
rect 2220 -2185 2240 -2165
rect 2260 -2185 2280 -2165
rect 2300 -2185 2320 -2165
rect 2340 -2185 2360 -2165
rect 2380 -2185 2400 -2165
rect 2420 -2185 2440 -2165
rect 2460 -2185 2480 -2165
rect 2500 -2185 2520 -2165
rect 2540 -2185 2560 -2165
rect 2590 -2185 2605 -2165
rect 105 -2195 2605 -2185
rect -70 -2210 85 -2200
rect -70 -2235 -60 -2210
rect -40 -2235 -20 -2210
rect 0 -2235 20 -2210
rect 40 -2235 60 -2210
rect -70 -2245 85 -2235
rect 105 -2260 2605 -2250
rect 105 -2280 120 -2260
rect 140 -2280 160 -2260
rect 180 -2280 200 -2260
rect 220 -2280 240 -2260
rect 260 -2280 280 -2260
rect 300 -2280 320 -2260
rect 340 -2280 360 -2260
rect 380 -2280 400 -2260
rect 420 -2280 440 -2260
rect 460 -2280 480 -2260
rect 500 -2280 520 -2260
rect 540 -2280 560 -2260
rect 580 -2280 600 -2260
rect 620 -2280 640 -2260
rect 660 -2280 680 -2260
rect 700 -2280 720 -2260
rect 740 -2280 760 -2260
rect 780 -2280 800 -2260
rect 820 -2280 840 -2260
rect 860 -2280 880 -2260
rect 900 -2280 920 -2260
rect 940 -2280 960 -2260
rect 980 -2280 1000 -2260
rect 1020 -2280 1040 -2260
rect 1060 -2280 1080 -2260
rect 1100 -2280 1120 -2260
rect 1140 -2280 1160 -2260
rect 1180 -2280 1200 -2260
rect 1220 -2280 1240 -2260
rect 1260 -2280 1280 -2260
rect 1300 -2280 1320 -2260
rect 1340 -2280 1360 -2260
rect 1380 -2280 1400 -2260
rect 1420 -2280 1440 -2260
rect 1460 -2280 1480 -2260
rect 1500 -2280 1520 -2260
rect 1540 -2280 1560 -2260
rect 1580 -2280 1600 -2260
rect 1620 -2280 1640 -2260
rect 1660 -2280 1680 -2260
rect 1700 -2280 1720 -2260
rect 1740 -2280 1760 -2260
rect 1780 -2280 1800 -2260
rect 1820 -2280 1840 -2260
rect 1860 -2280 1880 -2260
rect 1900 -2280 1920 -2260
rect 1940 -2280 1960 -2260
rect 1980 -2280 2000 -2260
rect 2020 -2280 2040 -2260
rect 2060 -2280 2080 -2260
rect 2100 -2280 2120 -2260
rect 2140 -2280 2160 -2260
rect 2180 -2280 2200 -2260
rect 2220 -2280 2240 -2260
rect 2260 -2280 2280 -2260
rect 2300 -2280 2320 -2260
rect 2340 -2280 2360 -2260
rect 2380 -2280 2400 -2260
rect 2420 -2280 2440 -2260
rect 2460 -2280 2480 -2260
rect 2500 -2280 2520 -2260
rect 2540 -2280 2560 -2260
rect 2590 -2280 2605 -2260
rect 105 -2290 2605 -2280
rect -70 -2305 85 -2295
rect -70 -2330 -60 -2305
rect -40 -2330 -20 -2305
rect 0 -2330 20 -2305
rect 40 -2330 60 -2305
rect -70 -2340 85 -2330
rect 105 -2355 2605 -2345
rect 105 -2375 120 -2355
rect 140 -2375 160 -2355
rect 180 -2375 200 -2355
rect 220 -2375 240 -2355
rect 260 -2375 280 -2355
rect 300 -2375 320 -2355
rect 340 -2375 360 -2355
rect 380 -2375 400 -2355
rect 420 -2375 440 -2355
rect 460 -2375 480 -2355
rect 500 -2375 520 -2355
rect 540 -2375 560 -2355
rect 580 -2375 600 -2355
rect 620 -2375 640 -2355
rect 660 -2375 680 -2355
rect 700 -2375 720 -2355
rect 740 -2375 760 -2355
rect 780 -2375 800 -2355
rect 820 -2375 840 -2355
rect 860 -2375 880 -2355
rect 900 -2375 920 -2355
rect 940 -2375 960 -2355
rect 980 -2375 1000 -2355
rect 1020 -2375 1040 -2355
rect 1060 -2375 1080 -2355
rect 1100 -2375 1120 -2355
rect 1140 -2375 1160 -2355
rect 1180 -2375 1200 -2355
rect 1220 -2375 1240 -2355
rect 1260 -2375 1280 -2355
rect 1300 -2375 1320 -2355
rect 1340 -2375 1360 -2355
rect 1380 -2375 1400 -2355
rect 1420 -2375 1440 -2355
rect 1460 -2375 1480 -2355
rect 1500 -2375 1520 -2355
rect 1540 -2375 1560 -2355
rect 1580 -2375 1600 -2355
rect 1620 -2375 1640 -2355
rect 1660 -2375 1680 -2355
rect 1700 -2375 1720 -2355
rect 1740 -2375 1760 -2355
rect 1780 -2375 1800 -2355
rect 1820 -2375 1840 -2355
rect 1860 -2375 1880 -2355
rect 1900 -2375 1920 -2355
rect 1940 -2375 1960 -2355
rect 1980 -2375 2000 -2355
rect 2020 -2375 2040 -2355
rect 2060 -2375 2080 -2355
rect 2100 -2375 2120 -2355
rect 2140 -2375 2160 -2355
rect 2180 -2375 2200 -2355
rect 2220 -2375 2240 -2355
rect 2260 -2375 2280 -2355
rect 2300 -2375 2320 -2355
rect 2340 -2375 2360 -2355
rect 2380 -2375 2400 -2355
rect 2420 -2375 2440 -2355
rect 2460 -2375 2480 -2355
rect 2500 -2375 2520 -2355
rect 2540 -2375 2560 -2355
rect 2590 -2375 2605 -2355
rect 105 -2385 2605 -2375
rect -70 -2400 85 -2390
rect -70 -2425 -60 -2400
rect -40 -2425 -20 -2400
rect 0 -2425 20 -2400
rect 40 -2425 60 -2400
rect -70 -2435 85 -2425
rect 105 -2450 2605 -2440
rect 105 -2470 120 -2450
rect 140 -2470 160 -2450
rect 180 -2470 200 -2450
rect 220 -2470 240 -2450
rect 260 -2470 280 -2450
rect 300 -2470 320 -2450
rect 340 -2470 360 -2450
rect 380 -2470 400 -2450
rect 420 -2470 440 -2450
rect 460 -2470 480 -2450
rect 500 -2470 520 -2450
rect 540 -2470 560 -2450
rect 580 -2470 600 -2450
rect 620 -2470 640 -2450
rect 660 -2470 680 -2450
rect 700 -2470 720 -2450
rect 740 -2470 760 -2450
rect 780 -2470 800 -2450
rect 820 -2470 840 -2450
rect 860 -2470 880 -2450
rect 900 -2470 920 -2450
rect 940 -2470 960 -2450
rect 980 -2470 1000 -2450
rect 1020 -2470 1040 -2450
rect 1060 -2470 1080 -2450
rect 1100 -2470 1120 -2450
rect 1140 -2470 1160 -2450
rect 1180 -2470 1200 -2450
rect 1220 -2470 1240 -2450
rect 1260 -2470 1280 -2450
rect 1300 -2470 1320 -2450
rect 1340 -2470 1360 -2450
rect 1380 -2470 1400 -2450
rect 1420 -2470 1440 -2450
rect 1460 -2470 1480 -2450
rect 1500 -2470 1520 -2450
rect 1540 -2470 1560 -2450
rect 1580 -2470 1600 -2450
rect 1620 -2470 1640 -2450
rect 1660 -2470 1680 -2450
rect 1700 -2470 1720 -2450
rect 1740 -2470 1760 -2450
rect 1780 -2470 1800 -2450
rect 1820 -2470 1840 -2450
rect 1860 -2470 1880 -2450
rect 1900 -2470 1920 -2450
rect 1940 -2470 1960 -2450
rect 1980 -2470 2000 -2450
rect 2020 -2470 2040 -2450
rect 2060 -2470 2080 -2450
rect 2100 -2470 2120 -2450
rect 2140 -2470 2160 -2450
rect 2180 -2470 2200 -2450
rect 2220 -2470 2240 -2450
rect 2260 -2470 2280 -2450
rect 2300 -2470 2320 -2450
rect 2340 -2470 2360 -2450
rect 2380 -2470 2400 -2450
rect 2420 -2470 2440 -2450
rect 2460 -2470 2480 -2450
rect 2500 -2470 2520 -2450
rect 2540 -2470 2560 -2450
rect 2590 -2470 2605 -2450
rect 105 -2480 2605 -2470
rect -70 -2495 85 -2485
rect -70 -2520 -60 -2495
rect -40 -2520 -20 -2495
rect 0 -2520 20 -2495
rect 40 -2520 60 -2495
rect -70 -2530 85 -2520
rect 105 -2545 2605 -2535
rect 105 -2565 120 -2545
rect 140 -2565 160 -2545
rect 180 -2565 200 -2545
rect 220 -2565 240 -2545
rect 260 -2565 280 -2545
rect 300 -2565 320 -2545
rect 340 -2565 360 -2545
rect 380 -2565 400 -2545
rect 420 -2565 440 -2545
rect 460 -2565 480 -2545
rect 500 -2565 520 -2545
rect 540 -2565 560 -2545
rect 580 -2565 600 -2545
rect 620 -2565 640 -2545
rect 660 -2565 680 -2545
rect 700 -2565 720 -2545
rect 740 -2565 760 -2545
rect 780 -2565 800 -2545
rect 820 -2565 840 -2545
rect 860 -2565 880 -2545
rect 900 -2565 920 -2545
rect 940 -2565 960 -2545
rect 980 -2565 1000 -2545
rect 1020 -2565 1040 -2545
rect 1060 -2565 1080 -2545
rect 1100 -2565 1120 -2545
rect 1140 -2565 1160 -2545
rect 1180 -2565 1200 -2545
rect 1220 -2565 1240 -2545
rect 1260 -2565 1280 -2545
rect 1300 -2565 1320 -2545
rect 1340 -2565 1360 -2545
rect 1380 -2565 1400 -2545
rect 1420 -2565 1440 -2545
rect 1460 -2565 1480 -2545
rect 1500 -2565 1520 -2545
rect 1540 -2565 1560 -2545
rect 1580 -2565 1600 -2545
rect 1620 -2565 1640 -2545
rect 1660 -2565 1680 -2545
rect 1700 -2565 1720 -2545
rect 1740 -2565 1760 -2545
rect 1780 -2565 1800 -2545
rect 1820 -2565 1840 -2545
rect 1860 -2565 1880 -2545
rect 1900 -2565 1920 -2545
rect 1940 -2565 1960 -2545
rect 1980 -2565 2000 -2545
rect 2020 -2565 2040 -2545
rect 2060 -2565 2080 -2545
rect 2100 -2565 2120 -2545
rect 2140 -2565 2160 -2545
rect 2180 -2565 2200 -2545
rect 2220 -2565 2240 -2545
rect 2260 -2565 2280 -2545
rect 2300 -2565 2320 -2545
rect 2340 -2565 2360 -2545
rect 2380 -2565 2400 -2545
rect 2420 -2565 2440 -2545
rect 2460 -2565 2480 -2545
rect 2500 -2565 2520 -2545
rect 2540 -2565 2560 -2545
rect 2590 -2565 2605 -2545
rect 105 -2575 2605 -2565
rect -70 -2590 85 -2580
rect -70 -2615 -60 -2590
rect -40 -2615 -20 -2590
rect 0 -2615 20 -2590
rect 40 -2615 60 -2590
rect -70 -2625 85 -2615
rect 105 -2640 2605 -2630
rect 105 -2660 120 -2640
rect 140 -2660 160 -2640
rect 180 -2660 200 -2640
rect 220 -2660 240 -2640
rect 260 -2660 280 -2640
rect 300 -2660 320 -2640
rect 340 -2660 360 -2640
rect 380 -2660 400 -2640
rect 420 -2660 440 -2640
rect 460 -2660 480 -2640
rect 500 -2660 520 -2640
rect 540 -2660 560 -2640
rect 580 -2660 600 -2640
rect 620 -2660 640 -2640
rect 660 -2660 680 -2640
rect 700 -2660 720 -2640
rect 740 -2660 760 -2640
rect 780 -2660 800 -2640
rect 820 -2660 840 -2640
rect 860 -2660 880 -2640
rect 900 -2660 920 -2640
rect 940 -2660 960 -2640
rect 980 -2660 1000 -2640
rect 1020 -2660 1040 -2640
rect 1060 -2660 1080 -2640
rect 1100 -2660 1120 -2640
rect 1140 -2660 1160 -2640
rect 1180 -2660 1200 -2640
rect 1220 -2660 1240 -2640
rect 1260 -2660 1280 -2640
rect 1300 -2660 1320 -2640
rect 1340 -2660 1360 -2640
rect 1380 -2660 1400 -2640
rect 1420 -2660 1440 -2640
rect 1460 -2660 1480 -2640
rect 1500 -2660 1520 -2640
rect 1540 -2660 1560 -2640
rect 1580 -2660 1600 -2640
rect 1620 -2660 1640 -2640
rect 1660 -2660 1680 -2640
rect 1700 -2660 1720 -2640
rect 1740 -2660 1760 -2640
rect 1780 -2660 1800 -2640
rect 1820 -2660 1840 -2640
rect 1860 -2660 1880 -2640
rect 1900 -2660 1920 -2640
rect 1940 -2660 1960 -2640
rect 1980 -2660 2000 -2640
rect 2020 -2660 2040 -2640
rect 2060 -2660 2080 -2640
rect 2100 -2660 2120 -2640
rect 2140 -2660 2160 -2640
rect 2180 -2660 2200 -2640
rect 2220 -2660 2240 -2640
rect 2260 -2660 2280 -2640
rect 2300 -2660 2320 -2640
rect 2340 -2660 2360 -2640
rect 2380 -2660 2400 -2640
rect 2420 -2660 2440 -2640
rect 2460 -2660 2480 -2640
rect 2500 -2660 2520 -2640
rect 2540 -2660 2560 -2640
rect 2590 -2660 2605 -2640
rect 105 -2670 2605 -2660
rect -70 -2685 85 -2675
rect -70 -2710 -60 -2685
rect -40 -2710 -20 -2685
rect 0 -2710 20 -2685
rect 40 -2710 60 -2685
rect -70 -2720 85 -2710
rect 105 -2735 2605 -2725
rect 105 -2755 120 -2735
rect 140 -2755 160 -2735
rect 180 -2755 200 -2735
rect 220 -2755 240 -2735
rect 260 -2755 280 -2735
rect 300 -2755 320 -2735
rect 340 -2755 360 -2735
rect 380 -2755 400 -2735
rect 420 -2755 440 -2735
rect 460 -2755 480 -2735
rect 500 -2755 520 -2735
rect 540 -2755 560 -2735
rect 580 -2755 600 -2735
rect 620 -2755 640 -2735
rect 660 -2755 680 -2735
rect 700 -2755 720 -2735
rect 740 -2755 760 -2735
rect 780 -2755 800 -2735
rect 820 -2755 840 -2735
rect 860 -2755 880 -2735
rect 900 -2755 920 -2735
rect 940 -2755 960 -2735
rect 980 -2755 1000 -2735
rect 1020 -2755 1040 -2735
rect 1060 -2755 1080 -2735
rect 1100 -2755 1120 -2735
rect 1140 -2755 1160 -2735
rect 1180 -2755 1200 -2735
rect 1220 -2755 1240 -2735
rect 1260 -2755 1280 -2735
rect 1300 -2755 1320 -2735
rect 1340 -2755 1360 -2735
rect 1380 -2755 1400 -2735
rect 1420 -2755 1440 -2735
rect 1460 -2755 1480 -2735
rect 1500 -2755 1520 -2735
rect 1540 -2755 1560 -2735
rect 1580 -2755 1600 -2735
rect 1620 -2755 1640 -2735
rect 1660 -2755 1680 -2735
rect 1700 -2755 1720 -2735
rect 1740 -2755 1760 -2735
rect 1780 -2755 1800 -2735
rect 1820 -2755 1840 -2735
rect 1860 -2755 1880 -2735
rect 1900 -2755 1920 -2735
rect 1940 -2755 1960 -2735
rect 1980 -2755 2000 -2735
rect 2020 -2755 2040 -2735
rect 2060 -2755 2080 -2735
rect 2100 -2755 2120 -2735
rect 2140 -2755 2160 -2735
rect 2180 -2755 2200 -2735
rect 2220 -2755 2240 -2735
rect 2260 -2755 2280 -2735
rect 2300 -2755 2320 -2735
rect 2340 -2755 2360 -2735
rect 2380 -2755 2400 -2735
rect 2420 -2755 2440 -2735
rect 2460 -2755 2480 -2735
rect 2500 -2755 2520 -2735
rect 2540 -2755 2560 -2735
rect 2590 -2755 2605 -2735
rect 105 -2775 2605 -2755
rect 105 -2795 120 -2775
rect 140 -2795 160 -2775
rect 180 -2795 200 -2775
rect 220 -2795 240 -2775
rect 260 -2795 280 -2775
rect 300 -2795 320 -2775
rect 340 -2795 360 -2775
rect 380 -2795 400 -2775
rect 420 -2795 440 -2775
rect 460 -2795 480 -2775
rect 500 -2795 520 -2775
rect 540 -2795 560 -2775
rect 580 -2795 600 -2775
rect 620 -2795 640 -2775
rect 660 -2795 680 -2775
rect 700 -2795 720 -2775
rect 740 -2795 760 -2775
rect 780 -2795 800 -2775
rect 820 -2795 840 -2775
rect 860 -2795 880 -2775
rect 900 -2795 920 -2775
rect 940 -2795 960 -2775
rect 980 -2795 1000 -2775
rect 1020 -2795 1040 -2775
rect 1060 -2795 1080 -2775
rect 1100 -2795 1120 -2775
rect 1140 -2795 1160 -2775
rect 1180 -2795 1200 -2775
rect 1220 -2795 1240 -2775
rect 1260 -2795 1280 -2775
rect 1300 -2795 1320 -2775
rect 1340 -2795 1360 -2775
rect 1380 -2795 1400 -2775
rect 1420 -2795 1440 -2775
rect 1460 -2795 1480 -2775
rect 1500 -2795 1520 -2775
rect 1540 -2795 1560 -2775
rect 1580 -2795 1600 -2775
rect 1620 -2795 1640 -2775
rect 1660 -2795 1680 -2775
rect 1700 -2795 1720 -2775
rect 1740 -2795 1760 -2775
rect 1780 -2795 1800 -2775
rect 1820 -2795 1840 -2775
rect 1860 -2795 1880 -2775
rect 1900 -2795 1920 -2775
rect 1940 -2795 1960 -2775
rect 1980 -2795 2000 -2775
rect 2020 -2795 2040 -2775
rect 2060 -2795 2080 -2775
rect 2100 -2795 2120 -2775
rect 2140 -2795 2160 -2775
rect 2180 -2795 2200 -2775
rect 2220 -2795 2240 -2775
rect 2260 -2795 2280 -2775
rect 2300 -2795 2320 -2775
rect 2340 -2795 2360 -2775
rect 2380 -2795 2400 -2775
rect 2420 -2795 2440 -2775
rect 2460 -2795 2480 -2775
rect 2500 -2795 2520 -2775
rect 2540 -2795 2560 -2775
rect 2590 -2795 2605 -2775
rect 105 -2805 2605 -2795
<< viali >>
rect 680 2240 700 2260
rect 720 2240 740 2260
rect 760 2240 780 2260
rect 800 2240 820 2260
rect 840 2240 860 2260
rect 880 2240 900 2260
rect 920 2240 940 2260
rect 960 2240 980 2260
rect 1000 2240 1020 2260
rect 1040 2240 1060 2260
rect 1080 2240 1100 2260
rect 1120 2240 1140 2260
rect 1160 2240 1180 2260
rect 1200 2240 1220 2260
rect 1240 2240 1260 2260
rect 1280 2240 1300 2260
rect 1320 2240 1340 2260
rect 1360 2240 1380 2260
rect 1400 2240 1420 2260
rect 1440 2240 1460 2260
rect 680 2197 700 2217
rect 720 2197 740 2217
rect 760 2197 780 2217
rect 800 2197 820 2217
rect 840 2197 860 2217
rect 880 2197 900 2217
rect 920 2197 940 2217
rect 960 2197 980 2217
rect 1000 2197 1020 2217
rect 1040 2197 1060 2217
rect 1080 2197 1100 2217
rect 1120 2197 1140 2217
rect 1160 2197 1180 2217
rect 1200 2197 1220 2217
rect 1240 2197 1260 2217
rect 1280 2197 1300 2217
rect 1320 2197 1340 2217
rect 1360 2197 1380 2217
rect 1400 2197 1420 2217
rect 1440 2197 1460 2217
rect 10 2155 30 2175
rect 50 2155 70 2175
rect 90 2155 110 2175
rect 130 2155 150 2175
rect 1760 2115 1780 2135
rect 1800 2115 1820 2135
rect 1840 2115 1860 2135
rect 1880 2115 1900 2135
rect 1920 2115 1940 2135
rect 1960 2115 1980 2135
rect 2000 2115 2020 2135
rect 2040 2115 2060 2135
rect 2080 2115 2100 2135
rect 2120 2115 2140 2135
rect 2160 2115 2180 2135
rect 2200 2115 2220 2135
rect 2240 2115 2260 2135
rect 2280 2115 2300 2135
rect 2320 2115 2340 2135
rect 2360 2115 2380 2135
rect 2400 2115 2420 2135
rect 2440 2115 2460 2135
rect 2480 2115 2500 2135
rect 2520 2115 2540 2135
rect 10 2075 30 2095
rect 50 2075 70 2095
rect 90 2075 110 2095
rect 130 2075 150 2095
rect 680 2033 700 2053
rect 720 2033 740 2053
rect 760 2033 780 2053
rect 800 2033 820 2053
rect 840 2033 860 2053
rect 880 2033 900 2053
rect 920 2033 940 2053
rect 960 2033 980 2053
rect 1000 2033 1020 2053
rect 1040 2033 1060 2053
rect 1080 2033 1100 2053
rect 1120 2033 1140 2053
rect 1160 2033 1180 2053
rect 1200 2033 1220 2053
rect 1240 2033 1260 2053
rect 1280 2033 1300 2053
rect 1320 2033 1340 2053
rect 1360 2033 1380 2053
rect 1400 2033 1420 2053
rect 1440 2033 1460 2053
rect 10 1990 30 2010
rect 50 1990 70 2010
rect 90 1990 110 2010
rect 130 1990 150 2010
rect 1760 1951 1780 1971
rect 1800 1951 1820 1971
rect 1840 1951 1860 1971
rect 1880 1951 1900 1971
rect 1920 1951 1940 1971
rect 1960 1951 1980 1971
rect 2000 1951 2020 1971
rect 2040 1951 2060 1971
rect 2080 1951 2100 1971
rect 2120 1951 2140 1971
rect 2160 1951 2180 1971
rect 2200 1951 2220 1971
rect 2240 1951 2260 1971
rect 2280 1951 2300 1971
rect 2320 1951 2340 1971
rect 2360 1951 2380 1971
rect 2400 1951 2420 1971
rect 2440 1951 2460 1971
rect 2480 1951 2500 1971
rect 2520 1951 2540 1971
rect 10 1910 30 1930
rect 50 1910 70 1930
rect 90 1910 110 1930
rect 130 1910 150 1930
rect 680 1869 700 1889
rect 720 1869 740 1889
rect 760 1869 780 1889
rect 800 1869 820 1889
rect 840 1869 860 1889
rect 880 1869 900 1889
rect 920 1869 940 1889
rect 960 1869 980 1889
rect 1000 1869 1020 1889
rect 1040 1869 1060 1889
rect 1080 1869 1100 1889
rect 1120 1869 1140 1889
rect 1160 1869 1180 1889
rect 1200 1869 1220 1889
rect 1240 1869 1260 1889
rect 1280 1869 1300 1889
rect 1320 1869 1340 1889
rect 1360 1869 1380 1889
rect 1400 1869 1420 1889
rect 1440 1869 1460 1889
rect 10 1830 30 1850
rect 50 1830 70 1850
rect 90 1830 110 1850
rect 130 1830 150 1850
rect 1760 1787 1780 1807
rect 1800 1787 1820 1807
rect 1840 1787 1860 1807
rect 1880 1787 1900 1807
rect 1920 1787 1940 1807
rect 1960 1787 1980 1807
rect 2000 1787 2020 1807
rect 2040 1787 2060 1807
rect 2080 1787 2100 1807
rect 2120 1787 2140 1807
rect 2160 1787 2180 1807
rect 2200 1787 2220 1807
rect 2240 1787 2260 1807
rect 2280 1787 2300 1807
rect 2320 1787 2340 1807
rect 2360 1787 2380 1807
rect 2400 1787 2420 1807
rect 2440 1787 2460 1807
rect 2480 1787 2500 1807
rect 2520 1787 2540 1807
rect 10 1745 30 1765
rect 50 1745 70 1765
rect 90 1745 110 1765
rect 130 1745 150 1765
rect 680 1705 700 1725
rect 720 1705 740 1725
rect 760 1705 780 1725
rect 800 1705 820 1725
rect 840 1705 860 1725
rect 880 1705 900 1725
rect 920 1705 940 1725
rect 960 1705 980 1725
rect 1000 1705 1020 1725
rect 1040 1705 1060 1725
rect 1080 1705 1100 1725
rect 1120 1705 1140 1725
rect 1160 1705 1180 1725
rect 1200 1705 1220 1725
rect 1240 1705 1260 1725
rect 1280 1705 1300 1725
rect 1320 1705 1340 1725
rect 1360 1705 1380 1725
rect 1400 1705 1420 1725
rect 1440 1705 1460 1725
rect 10 1665 30 1685
rect 50 1665 70 1685
rect 90 1665 110 1685
rect 130 1665 150 1685
rect 1760 1623 1780 1643
rect 1800 1623 1820 1643
rect 1840 1623 1860 1643
rect 1880 1623 1900 1643
rect 1920 1623 1940 1643
rect 1960 1623 1980 1643
rect 2000 1623 2020 1643
rect 2040 1623 2060 1643
rect 2080 1623 2100 1643
rect 2120 1623 2140 1643
rect 2160 1623 2180 1643
rect 2200 1623 2220 1643
rect 2240 1623 2260 1643
rect 2280 1623 2300 1643
rect 2320 1623 2340 1643
rect 2360 1623 2380 1643
rect 2400 1623 2420 1643
rect 2440 1623 2460 1643
rect 2480 1623 2500 1643
rect 2520 1623 2540 1643
rect 10 1580 30 1600
rect 50 1580 70 1600
rect 90 1580 110 1600
rect 130 1580 150 1600
rect 680 1541 700 1561
rect 720 1541 740 1561
rect 760 1541 780 1561
rect 800 1541 820 1561
rect 840 1541 860 1561
rect 880 1541 900 1561
rect 920 1541 940 1561
rect 960 1541 980 1561
rect 1000 1541 1020 1561
rect 1040 1541 1060 1561
rect 1080 1541 1100 1561
rect 1120 1541 1140 1561
rect 1160 1541 1180 1561
rect 1200 1541 1220 1561
rect 1240 1541 1260 1561
rect 1280 1541 1300 1561
rect 1320 1541 1340 1561
rect 1360 1541 1380 1561
rect 1400 1541 1420 1561
rect 1440 1541 1460 1561
rect 10 1500 30 1520
rect 50 1500 70 1520
rect 90 1500 110 1520
rect 130 1500 150 1520
rect 1760 1459 1780 1479
rect 1800 1459 1820 1479
rect 1840 1459 1860 1479
rect 1880 1459 1900 1479
rect 1920 1459 1940 1479
rect 1960 1459 1980 1479
rect 2000 1459 2020 1479
rect 2040 1459 2060 1479
rect 2080 1459 2100 1479
rect 2120 1459 2140 1479
rect 2160 1459 2180 1479
rect 2200 1459 2220 1479
rect 2240 1459 2260 1479
rect 2280 1459 2300 1479
rect 2320 1459 2340 1479
rect 2360 1459 2380 1479
rect 2400 1459 2420 1479
rect 2440 1459 2460 1479
rect 2480 1459 2500 1479
rect 2520 1459 2540 1479
rect 10 1420 30 1440
rect 50 1420 70 1440
rect 90 1420 110 1440
rect 130 1420 150 1440
rect 680 1377 700 1397
rect 720 1377 740 1397
rect 760 1377 780 1397
rect 800 1377 820 1397
rect 840 1377 860 1397
rect 880 1377 900 1397
rect 920 1377 940 1397
rect 960 1377 980 1397
rect 1000 1377 1020 1397
rect 1040 1377 1060 1397
rect 1080 1377 1100 1397
rect 1120 1377 1140 1397
rect 1160 1377 1180 1397
rect 1200 1377 1220 1397
rect 1240 1377 1260 1397
rect 1280 1377 1300 1397
rect 1320 1377 1340 1397
rect 1360 1377 1380 1397
rect 1400 1377 1420 1397
rect 1440 1377 1460 1397
rect 10 1335 30 1355
rect 50 1335 70 1355
rect 90 1335 110 1355
rect 130 1335 150 1355
rect 1760 1295 1780 1315
rect 1800 1295 1820 1315
rect 1840 1295 1860 1315
rect 1880 1295 1900 1315
rect 1920 1295 1940 1315
rect 1960 1295 1980 1315
rect 2000 1295 2020 1315
rect 2040 1295 2060 1315
rect 2080 1295 2100 1315
rect 2120 1295 2140 1315
rect 2160 1295 2180 1315
rect 2200 1295 2220 1315
rect 2240 1295 2260 1315
rect 2280 1295 2300 1315
rect 2320 1295 2340 1315
rect 2360 1295 2380 1315
rect 2400 1295 2420 1315
rect 2440 1295 2460 1315
rect 2480 1295 2500 1315
rect 2520 1295 2540 1315
rect 10 1255 30 1275
rect 50 1255 70 1275
rect 90 1255 110 1275
rect 130 1255 150 1275
rect 680 1213 700 1233
rect 720 1213 740 1233
rect 760 1213 780 1233
rect 800 1213 820 1233
rect 840 1213 860 1233
rect 880 1213 900 1233
rect 920 1213 940 1233
rect 960 1213 980 1233
rect 1000 1213 1020 1233
rect 1040 1213 1060 1233
rect 1080 1213 1100 1233
rect 1120 1213 1140 1233
rect 1160 1213 1180 1233
rect 1200 1213 1220 1233
rect 1240 1213 1260 1233
rect 1280 1213 1300 1233
rect 1320 1213 1340 1233
rect 1360 1213 1380 1233
rect 1400 1213 1420 1233
rect 1440 1213 1460 1233
rect 10 1170 30 1190
rect 50 1170 70 1190
rect 90 1170 110 1190
rect 130 1170 150 1190
rect 1760 1131 1780 1151
rect 1800 1131 1820 1151
rect 1840 1131 1860 1151
rect 1880 1131 1900 1151
rect 1920 1131 1940 1151
rect 1960 1131 1980 1151
rect 2000 1131 2020 1151
rect 2040 1131 2060 1151
rect 2080 1131 2100 1151
rect 2120 1131 2140 1151
rect 2160 1131 2180 1151
rect 2200 1131 2220 1151
rect 2240 1131 2260 1151
rect 2280 1131 2300 1151
rect 2320 1131 2340 1151
rect 2360 1131 2380 1151
rect 2400 1131 2420 1151
rect 2440 1131 2460 1151
rect 2480 1131 2500 1151
rect 2520 1131 2540 1151
rect 10 1090 30 1110
rect 50 1090 70 1110
rect 90 1090 110 1110
rect 130 1090 150 1110
rect 680 1049 700 1069
rect 720 1049 740 1069
rect 760 1049 780 1069
rect 800 1049 820 1069
rect 840 1049 860 1069
rect 880 1049 900 1069
rect 920 1049 940 1069
rect 960 1049 980 1069
rect 1000 1049 1020 1069
rect 1040 1049 1060 1069
rect 1080 1049 1100 1069
rect 1120 1049 1140 1069
rect 1160 1049 1180 1069
rect 1200 1049 1220 1069
rect 1240 1049 1260 1069
rect 1280 1049 1300 1069
rect 1320 1049 1340 1069
rect 1360 1049 1380 1069
rect 1400 1049 1420 1069
rect 1440 1049 1460 1069
rect 10 1010 30 1030
rect 50 1010 70 1030
rect 90 1010 110 1030
rect 130 1010 150 1030
rect 1760 967 1780 987
rect 1800 967 1820 987
rect 1840 967 1860 987
rect 1880 967 1900 987
rect 1920 967 1940 987
rect 1960 967 1980 987
rect 2000 967 2020 987
rect 2040 967 2060 987
rect 2080 967 2100 987
rect 2120 967 2140 987
rect 2160 967 2180 987
rect 2200 967 2220 987
rect 2240 967 2260 987
rect 2280 967 2300 987
rect 2320 967 2340 987
rect 2360 967 2380 987
rect 2400 967 2420 987
rect 2440 967 2460 987
rect 2480 967 2500 987
rect 2520 967 2540 987
rect 10 925 30 945
rect 50 925 70 945
rect 90 925 110 945
rect 130 925 150 945
rect 680 885 700 905
rect 720 885 740 905
rect 760 885 780 905
rect 800 885 820 905
rect 840 885 860 905
rect 880 885 900 905
rect 920 885 940 905
rect 960 885 980 905
rect 1000 885 1020 905
rect 1040 885 1060 905
rect 1080 885 1100 905
rect 1120 885 1140 905
rect 1160 885 1180 905
rect 1200 885 1220 905
rect 1240 885 1260 905
rect 1280 885 1300 905
rect 1320 885 1340 905
rect 1360 885 1380 905
rect 1400 885 1420 905
rect 1440 885 1460 905
rect 10 845 30 865
rect 50 845 70 865
rect 90 845 110 865
rect 130 845 150 865
rect 1760 803 1780 823
rect 1800 803 1820 823
rect 1840 803 1860 823
rect 1880 803 1900 823
rect 1920 803 1940 823
rect 1960 803 1980 823
rect 2000 803 2020 823
rect 2040 803 2060 823
rect 2080 803 2100 823
rect 2120 803 2140 823
rect 2160 803 2180 823
rect 2200 803 2220 823
rect 2240 803 2260 823
rect 2280 803 2300 823
rect 2320 803 2340 823
rect 2360 803 2380 823
rect 2400 803 2420 823
rect 2440 803 2460 823
rect 2480 803 2500 823
rect 2520 803 2540 823
rect 10 760 30 780
rect 50 760 70 780
rect 90 760 110 780
rect 130 760 150 780
rect 680 721 700 741
rect 720 721 740 741
rect 760 721 780 741
rect 800 721 820 741
rect 840 721 860 741
rect 880 721 900 741
rect 920 721 940 741
rect 960 721 980 741
rect 1000 721 1020 741
rect 1040 721 1060 741
rect 1080 721 1100 741
rect 1120 721 1140 741
rect 1160 721 1180 741
rect 1200 721 1220 741
rect 1240 721 1260 741
rect 1280 721 1300 741
rect 1320 721 1340 741
rect 1360 721 1380 741
rect 1400 721 1420 741
rect 1440 721 1460 741
rect 10 680 30 700
rect 50 680 70 700
rect 90 680 110 700
rect 130 680 150 700
rect 1760 639 1780 659
rect 1800 639 1820 659
rect 1840 639 1860 659
rect 1880 639 1900 659
rect 1920 639 1940 659
rect 1960 639 1980 659
rect 2000 639 2020 659
rect 2040 639 2060 659
rect 2080 639 2100 659
rect 2120 639 2140 659
rect 2160 639 2180 659
rect 2200 639 2220 659
rect 2240 639 2260 659
rect 2280 639 2300 659
rect 2320 639 2340 659
rect 2360 639 2380 659
rect 2400 639 2420 659
rect 2440 639 2460 659
rect 2480 639 2500 659
rect 2520 639 2540 659
rect 10 600 30 620
rect 50 600 70 620
rect 90 600 110 620
rect 130 600 150 620
rect 680 557 700 577
rect 720 557 740 577
rect 760 557 780 577
rect 800 557 820 577
rect 840 557 860 577
rect 880 557 900 577
rect 920 557 940 577
rect 960 557 980 577
rect 1000 557 1020 577
rect 1040 557 1060 577
rect 1080 557 1100 577
rect 1120 557 1140 577
rect 1160 557 1180 577
rect 1200 557 1220 577
rect 1240 557 1260 577
rect 1280 557 1300 577
rect 1320 557 1340 577
rect 1360 557 1380 577
rect 1400 557 1420 577
rect 1440 557 1460 577
rect 10 515 30 535
rect 50 515 70 535
rect 90 515 110 535
rect 130 515 150 535
rect 1760 475 1780 495
rect 1800 475 1820 495
rect 1840 475 1860 495
rect 1880 475 1900 495
rect 1920 475 1940 495
rect 1960 475 1980 495
rect 2000 475 2020 495
rect 2040 475 2060 495
rect 2080 475 2100 495
rect 2120 475 2140 495
rect 2160 475 2180 495
rect 2200 475 2220 495
rect 2240 475 2260 495
rect 2280 475 2300 495
rect 2320 475 2340 495
rect 2360 475 2380 495
rect 2400 475 2420 495
rect 2440 475 2460 495
rect 2480 475 2500 495
rect 2520 475 2540 495
rect 10 435 30 455
rect 50 435 70 455
rect 90 435 110 455
rect 130 435 150 455
rect 680 393 700 413
rect 720 393 740 413
rect 760 393 780 413
rect 800 393 820 413
rect 840 393 860 413
rect 880 393 900 413
rect 920 393 940 413
rect 960 393 980 413
rect 1000 393 1020 413
rect 1040 393 1060 413
rect 1080 393 1100 413
rect 1120 393 1140 413
rect 1160 393 1180 413
rect 1200 393 1220 413
rect 1240 393 1260 413
rect 1280 393 1300 413
rect 1320 393 1340 413
rect 1360 393 1380 413
rect 1400 393 1420 413
rect 1440 393 1460 413
rect 10 355 30 375
rect 50 355 70 375
rect 90 355 110 375
rect 130 355 150 375
rect 1760 311 1780 331
rect 1800 311 1820 331
rect 1840 311 1860 331
rect 1880 311 1900 331
rect 1920 311 1940 331
rect 1960 311 1980 331
rect 2000 311 2020 331
rect 2040 311 2060 331
rect 2080 311 2100 331
rect 2120 311 2140 331
rect 2160 311 2180 331
rect 2200 311 2220 331
rect 2240 311 2260 331
rect 2280 311 2300 331
rect 2320 311 2340 331
rect 2360 311 2380 331
rect 2400 311 2420 331
rect 2440 311 2460 331
rect 2480 311 2500 331
rect 2520 311 2540 331
rect 10 270 30 290
rect 50 270 70 290
rect 90 270 110 290
rect 130 270 150 290
rect 680 229 700 249
rect 720 229 740 249
rect 760 229 780 249
rect 800 229 820 249
rect 840 229 860 249
rect 880 229 900 249
rect 920 229 940 249
rect 960 229 980 249
rect 1000 229 1020 249
rect 1040 229 1060 249
rect 1080 229 1100 249
rect 1120 229 1140 249
rect 1160 229 1180 249
rect 1200 229 1220 249
rect 1240 229 1260 249
rect 1280 229 1300 249
rect 1320 229 1340 249
rect 1360 229 1380 249
rect 1400 229 1420 249
rect 1440 229 1460 249
rect 10 190 30 210
rect 50 190 70 210
rect 90 190 110 210
rect 130 190 150 210
rect 1760 147 1780 167
rect 1800 147 1820 167
rect 1840 147 1860 167
rect 1880 147 1900 167
rect 1920 147 1940 167
rect 1960 147 1980 167
rect 2000 147 2020 167
rect 2040 147 2060 167
rect 2080 147 2100 167
rect 2120 147 2140 167
rect 2160 147 2180 167
rect 2200 147 2220 167
rect 2240 147 2260 167
rect 2280 147 2300 167
rect 2320 147 2340 167
rect 2360 147 2380 167
rect 2400 147 2420 167
rect 2440 147 2460 167
rect 2480 147 2500 167
rect 2520 147 2540 167
rect 10 110 30 130
rect 50 110 70 130
rect 90 110 110 130
rect 130 110 150 130
rect 680 65 700 85
rect 720 65 740 85
rect 760 65 780 85
rect 800 65 820 85
rect 840 65 860 85
rect 880 65 900 85
rect 920 65 940 85
rect 960 65 980 85
rect 1000 65 1020 85
rect 1040 65 1060 85
rect 1080 65 1100 85
rect 1120 65 1140 85
rect 1160 65 1180 85
rect 1200 65 1220 85
rect 1240 65 1260 85
rect 1280 65 1300 85
rect 1320 65 1340 85
rect 1360 65 1380 85
rect 1400 65 1420 85
rect 1440 65 1460 85
rect 680 25 700 45
rect 720 25 740 45
rect 760 25 780 45
rect 800 25 820 45
rect 840 25 860 45
rect 880 25 900 45
rect 920 25 940 45
rect 960 25 980 45
rect 1000 25 1020 45
rect 1040 25 1060 45
rect 1080 25 1100 45
rect 1120 25 1140 45
rect 1160 25 1180 45
rect 1200 25 1220 45
rect 1240 25 1260 45
rect 1280 25 1300 45
rect 1320 25 1340 45
rect 1360 25 1380 45
rect 1400 25 1420 45
rect 1440 25 1460 45
rect 1760 -245 1780 -225
rect 1800 -245 1820 -225
rect 1840 -245 1860 -225
rect 1880 -245 1900 -225
rect 1920 -245 1940 -225
rect 1960 -245 1980 -225
rect 2000 -245 2020 -225
rect 2040 -245 2060 -225
rect 2080 -245 2100 -225
rect 2120 -245 2140 -225
rect 2160 -245 2180 -225
rect 2200 -245 2220 -225
rect 2240 -245 2260 -225
rect 2280 -245 2300 -225
rect 2320 -245 2340 -225
rect 2360 -245 2380 -225
rect 2400 -245 2420 -225
rect 2440 -245 2460 -225
rect 2480 -245 2500 -225
rect 2520 -245 2540 -225
rect 1760 -285 1780 -265
rect 1800 -285 1820 -265
rect 1840 -285 1860 -265
rect 1880 -285 1900 -265
rect 1920 -285 1940 -265
rect 1960 -285 1980 -265
rect 2000 -285 2020 -265
rect 2040 -285 2060 -265
rect 2080 -285 2100 -265
rect 2120 -285 2140 -265
rect 2160 -285 2180 -265
rect 2200 -285 2220 -265
rect 2240 -285 2260 -265
rect 2280 -285 2300 -265
rect 2320 -285 2340 -265
rect 2360 -285 2380 -265
rect 2400 -285 2420 -265
rect 2440 -285 2460 -265
rect 2480 -285 2500 -265
rect 2520 -285 2540 -265
rect -60 -335 -40 -310
rect -20 -335 0 -310
rect 20 -335 40 -310
rect 60 -335 80 -310
rect 680 -380 700 -360
rect 720 -380 740 -360
rect 760 -380 780 -360
rect 800 -380 820 -360
rect 840 -380 860 -360
rect 880 -380 900 -360
rect 920 -380 940 -360
rect 960 -380 980 -360
rect 1000 -380 1020 -360
rect 1040 -380 1060 -360
rect 1080 -380 1100 -360
rect 1120 -380 1140 -360
rect 1160 -380 1180 -360
rect 1200 -380 1220 -360
rect 1240 -380 1260 -360
rect 1280 -380 1300 -360
rect 1320 -380 1340 -360
rect 1360 -380 1380 -360
rect 1400 -380 1420 -360
rect 1440 -380 1460 -360
rect -60 -430 -40 -405
rect -20 -430 0 -405
rect 20 -430 40 -405
rect 60 -430 80 -405
rect 1760 -475 1780 -455
rect 1800 -475 1820 -455
rect 1840 -475 1860 -455
rect 1880 -475 1900 -455
rect 1920 -475 1940 -455
rect 1960 -475 1980 -455
rect 2000 -475 2020 -455
rect 2040 -475 2060 -455
rect 2080 -475 2100 -455
rect 2120 -475 2140 -455
rect 2160 -475 2180 -455
rect 2200 -475 2220 -455
rect 2240 -475 2260 -455
rect 2280 -475 2300 -455
rect 2320 -475 2340 -455
rect 2360 -475 2380 -455
rect 2400 -475 2420 -455
rect 2440 -475 2460 -455
rect 2480 -475 2500 -455
rect 2520 -475 2540 -455
rect -60 -525 -40 -500
rect -20 -525 0 -500
rect 20 -525 40 -500
rect 60 -525 80 -500
rect 680 -570 700 -550
rect 720 -570 740 -550
rect 760 -570 780 -550
rect 800 -570 820 -550
rect 840 -570 860 -550
rect 880 -570 900 -550
rect 920 -570 940 -550
rect 960 -570 980 -550
rect 1000 -570 1020 -550
rect 1040 -570 1060 -550
rect 1080 -570 1100 -550
rect 1120 -570 1140 -550
rect 1160 -570 1180 -550
rect 1200 -570 1220 -550
rect 1240 -570 1260 -550
rect 1280 -570 1300 -550
rect 1320 -570 1340 -550
rect 1360 -570 1380 -550
rect 1400 -570 1420 -550
rect 1440 -570 1460 -550
rect -60 -620 -40 -595
rect -20 -620 0 -595
rect 20 -620 40 -595
rect 60 -620 80 -595
rect 1760 -665 1780 -645
rect 1800 -665 1820 -645
rect 1840 -665 1860 -645
rect 1880 -665 1900 -645
rect 1920 -665 1940 -645
rect 1960 -665 1980 -645
rect 2000 -665 2020 -645
rect 2040 -665 2060 -645
rect 2080 -665 2100 -645
rect 2120 -665 2140 -645
rect 2160 -665 2180 -645
rect 2200 -665 2220 -645
rect 2240 -665 2260 -645
rect 2280 -665 2300 -645
rect 2320 -665 2340 -645
rect 2360 -665 2380 -645
rect 2400 -665 2420 -645
rect 2440 -665 2460 -645
rect 2480 -665 2500 -645
rect 2520 -665 2540 -645
rect -60 -715 -40 -690
rect -20 -715 0 -690
rect 20 -715 40 -690
rect 60 -715 80 -690
rect 680 -760 700 -740
rect 720 -760 740 -740
rect 760 -760 780 -740
rect 800 -760 820 -740
rect 840 -760 860 -740
rect 880 -760 900 -740
rect 920 -760 940 -740
rect 960 -760 980 -740
rect 1000 -760 1020 -740
rect 1040 -760 1060 -740
rect 1080 -760 1100 -740
rect 1120 -760 1140 -740
rect 1160 -760 1180 -740
rect 1200 -760 1220 -740
rect 1240 -760 1260 -740
rect 1280 -760 1300 -740
rect 1320 -760 1340 -740
rect 1360 -760 1380 -740
rect 1400 -760 1420 -740
rect 1440 -760 1460 -740
rect -60 -810 -40 -785
rect -20 -810 0 -785
rect 20 -810 40 -785
rect 60 -810 80 -785
rect 1760 -855 1780 -835
rect 1800 -855 1820 -835
rect 1840 -855 1860 -835
rect 1880 -855 1900 -835
rect 1920 -855 1940 -835
rect 1960 -855 1980 -835
rect 2000 -855 2020 -835
rect 2040 -855 2060 -835
rect 2080 -855 2100 -835
rect 2120 -855 2140 -835
rect 2160 -855 2180 -835
rect 2200 -855 2220 -835
rect 2240 -855 2260 -835
rect 2280 -855 2300 -835
rect 2320 -855 2340 -835
rect 2360 -855 2380 -835
rect 2400 -855 2420 -835
rect 2440 -855 2460 -835
rect 2480 -855 2500 -835
rect 2520 -855 2540 -835
rect -60 -905 -40 -880
rect -20 -905 0 -880
rect 20 -905 40 -880
rect 60 -905 80 -880
rect 680 -950 700 -930
rect 720 -950 740 -930
rect 760 -950 780 -930
rect 800 -950 820 -930
rect 840 -950 860 -930
rect 880 -950 900 -930
rect 920 -950 940 -930
rect 960 -950 980 -930
rect 1000 -950 1020 -930
rect 1040 -950 1060 -930
rect 1080 -950 1100 -930
rect 1120 -950 1140 -930
rect 1160 -950 1180 -930
rect 1200 -950 1220 -930
rect 1240 -950 1260 -930
rect 1280 -950 1300 -930
rect 1320 -950 1340 -930
rect 1360 -950 1380 -930
rect 1400 -950 1420 -930
rect 1440 -950 1460 -930
rect -60 -1000 -40 -975
rect -20 -1000 0 -975
rect 20 -1000 40 -975
rect 60 -1000 80 -975
rect 1760 -1045 1780 -1025
rect 1800 -1045 1820 -1025
rect 1840 -1045 1860 -1025
rect 1880 -1045 1900 -1025
rect 1920 -1045 1940 -1025
rect 1960 -1045 1980 -1025
rect 2000 -1045 2020 -1025
rect 2040 -1045 2060 -1025
rect 2080 -1045 2100 -1025
rect 2120 -1045 2140 -1025
rect 2160 -1045 2180 -1025
rect 2200 -1045 2220 -1025
rect 2240 -1045 2260 -1025
rect 2280 -1045 2300 -1025
rect 2320 -1045 2340 -1025
rect 2360 -1045 2380 -1025
rect 2400 -1045 2420 -1025
rect 2440 -1045 2460 -1025
rect 2480 -1045 2500 -1025
rect 2520 -1045 2540 -1025
rect -60 -1095 -40 -1070
rect -20 -1095 0 -1070
rect 20 -1095 40 -1070
rect 60 -1095 80 -1070
rect 680 -1140 700 -1120
rect 720 -1140 740 -1120
rect 760 -1140 780 -1120
rect 800 -1140 820 -1120
rect 840 -1140 860 -1120
rect 880 -1140 900 -1120
rect 920 -1140 940 -1120
rect 960 -1140 980 -1120
rect 1000 -1140 1020 -1120
rect 1040 -1140 1060 -1120
rect 1080 -1140 1100 -1120
rect 1120 -1140 1140 -1120
rect 1160 -1140 1180 -1120
rect 1200 -1140 1220 -1120
rect 1240 -1140 1260 -1120
rect 1280 -1140 1300 -1120
rect 1320 -1140 1340 -1120
rect 1360 -1140 1380 -1120
rect 1400 -1140 1420 -1120
rect 1440 -1140 1460 -1120
rect -60 -1190 -40 -1165
rect -20 -1190 0 -1165
rect 20 -1190 40 -1165
rect 60 -1190 80 -1165
rect 1760 -1235 1780 -1215
rect 1800 -1235 1820 -1215
rect 1840 -1235 1860 -1215
rect 1880 -1235 1900 -1215
rect 1920 -1235 1940 -1215
rect 1960 -1235 1980 -1215
rect 2000 -1235 2020 -1215
rect 2040 -1235 2060 -1215
rect 2080 -1235 2100 -1215
rect 2120 -1235 2140 -1215
rect 2160 -1235 2180 -1215
rect 2200 -1235 2220 -1215
rect 2240 -1235 2260 -1215
rect 2280 -1235 2300 -1215
rect 2320 -1235 2340 -1215
rect 2360 -1235 2380 -1215
rect 2400 -1235 2420 -1215
rect 2440 -1235 2460 -1215
rect 2480 -1235 2500 -1215
rect 2520 -1235 2540 -1215
rect -60 -1285 -40 -1260
rect -20 -1285 0 -1260
rect 20 -1285 40 -1260
rect 60 -1285 80 -1260
rect 680 -1330 700 -1310
rect 720 -1330 740 -1310
rect 760 -1330 780 -1310
rect 800 -1330 820 -1310
rect 840 -1330 860 -1310
rect 880 -1330 900 -1310
rect 920 -1330 940 -1310
rect 960 -1330 980 -1310
rect 1000 -1330 1020 -1310
rect 1040 -1330 1060 -1310
rect 1080 -1330 1100 -1310
rect 1120 -1330 1140 -1310
rect 1160 -1330 1180 -1310
rect 1200 -1330 1220 -1310
rect 1240 -1330 1260 -1310
rect 1280 -1330 1300 -1310
rect 1320 -1330 1340 -1310
rect 1360 -1330 1380 -1310
rect 1400 -1330 1420 -1310
rect 1440 -1330 1460 -1310
rect -60 -1380 -40 -1355
rect -20 -1380 0 -1355
rect 20 -1380 40 -1355
rect 60 -1380 80 -1355
rect 1760 -1425 1780 -1405
rect 1800 -1425 1820 -1405
rect 1840 -1425 1860 -1405
rect 1880 -1425 1900 -1405
rect 1920 -1425 1940 -1405
rect 1960 -1425 1980 -1405
rect 2000 -1425 2020 -1405
rect 2040 -1425 2060 -1405
rect 2080 -1425 2100 -1405
rect 2120 -1425 2140 -1405
rect 2160 -1425 2180 -1405
rect 2200 -1425 2220 -1405
rect 2240 -1425 2260 -1405
rect 2280 -1425 2300 -1405
rect 2320 -1425 2340 -1405
rect 2360 -1425 2380 -1405
rect 2400 -1425 2420 -1405
rect 2440 -1425 2460 -1405
rect 2480 -1425 2500 -1405
rect 2520 -1425 2540 -1405
rect -60 -1475 -40 -1450
rect -20 -1475 0 -1450
rect 20 -1475 40 -1450
rect 60 -1475 80 -1450
rect 680 -1520 700 -1500
rect 720 -1520 740 -1500
rect 760 -1520 780 -1500
rect 800 -1520 820 -1500
rect 840 -1520 860 -1500
rect 880 -1520 900 -1500
rect 920 -1520 940 -1500
rect 960 -1520 980 -1500
rect 1000 -1520 1020 -1500
rect 1040 -1520 1060 -1500
rect 1080 -1520 1100 -1500
rect 1120 -1520 1140 -1500
rect 1160 -1520 1180 -1500
rect 1200 -1520 1220 -1500
rect 1240 -1520 1260 -1500
rect 1280 -1520 1300 -1500
rect 1320 -1520 1340 -1500
rect 1360 -1520 1380 -1500
rect 1400 -1520 1420 -1500
rect 1440 -1520 1460 -1500
rect -60 -1570 -40 -1545
rect -20 -1570 0 -1545
rect 20 -1570 40 -1545
rect 60 -1570 80 -1545
rect 1760 -1615 1780 -1595
rect 1800 -1615 1820 -1595
rect 1840 -1615 1860 -1595
rect 1880 -1615 1900 -1595
rect 1920 -1615 1940 -1595
rect 1960 -1615 1980 -1595
rect 2000 -1615 2020 -1595
rect 2040 -1615 2060 -1595
rect 2080 -1615 2100 -1595
rect 2120 -1615 2140 -1595
rect 2160 -1615 2180 -1595
rect 2200 -1615 2220 -1595
rect 2240 -1615 2260 -1595
rect 2280 -1615 2300 -1595
rect 2320 -1615 2340 -1595
rect 2360 -1615 2380 -1595
rect 2400 -1615 2420 -1595
rect 2440 -1615 2460 -1595
rect 2480 -1615 2500 -1595
rect 2520 -1615 2540 -1595
rect -60 -1665 -40 -1640
rect -20 -1665 0 -1640
rect 20 -1665 40 -1640
rect 60 -1665 80 -1640
rect 680 -1710 700 -1690
rect 720 -1710 740 -1690
rect 760 -1710 780 -1690
rect 800 -1710 820 -1690
rect 840 -1710 860 -1690
rect 880 -1710 900 -1690
rect 920 -1710 940 -1690
rect 960 -1710 980 -1690
rect 1000 -1710 1020 -1690
rect 1040 -1710 1060 -1690
rect 1080 -1710 1100 -1690
rect 1120 -1710 1140 -1690
rect 1160 -1710 1180 -1690
rect 1200 -1710 1220 -1690
rect 1240 -1710 1260 -1690
rect 1280 -1710 1300 -1690
rect 1320 -1710 1340 -1690
rect 1360 -1710 1380 -1690
rect 1400 -1710 1420 -1690
rect 1440 -1710 1460 -1690
rect -60 -1760 -40 -1735
rect -20 -1760 0 -1735
rect 20 -1760 40 -1735
rect 60 -1760 80 -1735
rect 1760 -1805 1780 -1785
rect 1800 -1805 1820 -1785
rect 1840 -1805 1860 -1785
rect 1880 -1805 1900 -1785
rect 1920 -1805 1940 -1785
rect 1960 -1805 1980 -1785
rect 2000 -1805 2020 -1785
rect 2040 -1805 2060 -1785
rect 2080 -1805 2100 -1785
rect 2120 -1805 2140 -1785
rect 2160 -1805 2180 -1785
rect 2200 -1805 2220 -1785
rect 2240 -1805 2260 -1785
rect 2280 -1805 2300 -1785
rect 2320 -1805 2340 -1785
rect 2360 -1805 2380 -1785
rect 2400 -1805 2420 -1785
rect 2440 -1805 2460 -1785
rect 2480 -1805 2500 -1785
rect 2520 -1805 2540 -1785
rect -60 -1855 -40 -1830
rect -20 -1855 0 -1830
rect 20 -1855 40 -1830
rect 60 -1855 80 -1830
rect 680 -1900 700 -1880
rect 720 -1900 740 -1880
rect 760 -1900 780 -1880
rect 800 -1900 820 -1880
rect 840 -1900 860 -1880
rect 880 -1900 900 -1880
rect 920 -1900 940 -1880
rect 960 -1900 980 -1880
rect 1000 -1900 1020 -1880
rect 1040 -1900 1060 -1880
rect 1080 -1900 1100 -1880
rect 1120 -1900 1140 -1880
rect 1160 -1900 1180 -1880
rect 1200 -1900 1220 -1880
rect 1240 -1900 1260 -1880
rect 1280 -1900 1300 -1880
rect 1320 -1900 1340 -1880
rect 1360 -1900 1380 -1880
rect 1400 -1900 1420 -1880
rect 1440 -1900 1460 -1880
rect -60 -1950 -40 -1925
rect -20 -1950 0 -1925
rect 20 -1950 40 -1925
rect 60 -1950 80 -1925
rect 1760 -1995 1780 -1975
rect 1800 -1995 1820 -1975
rect 1840 -1995 1860 -1975
rect 1880 -1995 1900 -1975
rect 1920 -1995 1940 -1975
rect 1960 -1995 1980 -1975
rect 2000 -1995 2020 -1975
rect 2040 -1995 2060 -1975
rect 2080 -1995 2100 -1975
rect 2120 -1995 2140 -1975
rect 2160 -1995 2180 -1975
rect 2200 -1995 2220 -1975
rect 2240 -1995 2260 -1975
rect 2280 -1995 2300 -1975
rect 2320 -1995 2340 -1975
rect 2360 -1995 2380 -1975
rect 2400 -1995 2420 -1975
rect 2440 -1995 2460 -1975
rect 2480 -1995 2500 -1975
rect 2520 -1995 2540 -1975
rect -60 -2045 -40 -2020
rect -20 -2045 0 -2020
rect 20 -2045 40 -2020
rect 60 -2045 80 -2020
rect 680 -2090 700 -2070
rect 720 -2090 740 -2070
rect 760 -2090 780 -2070
rect 800 -2090 820 -2070
rect 840 -2090 860 -2070
rect 880 -2090 900 -2070
rect 920 -2090 940 -2070
rect 960 -2090 980 -2070
rect 1000 -2090 1020 -2070
rect 1040 -2090 1060 -2070
rect 1080 -2090 1100 -2070
rect 1120 -2090 1140 -2070
rect 1160 -2090 1180 -2070
rect 1200 -2090 1220 -2070
rect 1240 -2090 1260 -2070
rect 1280 -2090 1300 -2070
rect 1320 -2090 1340 -2070
rect 1360 -2090 1380 -2070
rect 1400 -2090 1420 -2070
rect 1440 -2090 1460 -2070
rect -60 -2140 -40 -2115
rect -20 -2140 0 -2115
rect 20 -2140 40 -2115
rect 60 -2140 80 -2115
rect 1760 -2185 1780 -2165
rect 1800 -2185 1820 -2165
rect 1840 -2185 1860 -2165
rect 1880 -2185 1900 -2165
rect 1920 -2185 1940 -2165
rect 1960 -2185 1980 -2165
rect 2000 -2185 2020 -2165
rect 2040 -2185 2060 -2165
rect 2080 -2185 2100 -2165
rect 2120 -2185 2140 -2165
rect 2160 -2185 2180 -2165
rect 2200 -2185 2220 -2165
rect 2240 -2185 2260 -2165
rect 2280 -2185 2300 -2165
rect 2320 -2185 2340 -2165
rect 2360 -2185 2380 -2165
rect 2400 -2185 2420 -2165
rect 2440 -2185 2460 -2165
rect 2480 -2185 2500 -2165
rect 2520 -2185 2540 -2165
rect -60 -2235 -40 -2210
rect -20 -2235 0 -2210
rect 20 -2235 40 -2210
rect 60 -2235 80 -2210
rect 680 -2280 700 -2260
rect 720 -2280 740 -2260
rect 760 -2280 780 -2260
rect 800 -2280 820 -2260
rect 840 -2280 860 -2260
rect 880 -2280 900 -2260
rect 920 -2280 940 -2260
rect 960 -2280 980 -2260
rect 1000 -2280 1020 -2260
rect 1040 -2280 1060 -2260
rect 1080 -2280 1100 -2260
rect 1120 -2280 1140 -2260
rect 1160 -2280 1180 -2260
rect 1200 -2280 1220 -2260
rect 1240 -2280 1260 -2260
rect 1280 -2280 1300 -2260
rect 1320 -2280 1340 -2260
rect 1360 -2280 1380 -2260
rect 1400 -2280 1420 -2260
rect 1440 -2280 1460 -2260
rect -60 -2330 -40 -2305
rect -20 -2330 0 -2305
rect 20 -2330 40 -2305
rect 60 -2330 80 -2305
rect 1760 -2375 1780 -2355
rect 1800 -2375 1820 -2355
rect 1840 -2375 1860 -2355
rect 1880 -2375 1900 -2355
rect 1920 -2375 1940 -2355
rect 1960 -2375 1980 -2355
rect 2000 -2375 2020 -2355
rect 2040 -2375 2060 -2355
rect 2080 -2375 2100 -2355
rect 2120 -2375 2140 -2355
rect 2160 -2375 2180 -2355
rect 2200 -2375 2220 -2355
rect 2240 -2375 2260 -2355
rect 2280 -2375 2300 -2355
rect 2320 -2375 2340 -2355
rect 2360 -2375 2380 -2355
rect 2400 -2375 2420 -2355
rect 2440 -2375 2460 -2355
rect 2480 -2375 2500 -2355
rect 2520 -2375 2540 -2355
rect -60 -2425 -40 -2400
rect -20 -2425 0 -2400
rect 20 -2425 40 -2400
rect 60 -2425 80 -2400
rect 680 -2470 700 -2450
rect 720 -2470 740 -2450
rect 760 -2470 780 -2450
rect 800 -2470 820 -2450
rect 840 -2470 860 -2450
rect 880 -2470 900 -2450
rect 920 -2470 940 -2450
rect 960 -2470 980 -2450
rect 1000 -2470 1020 -2450
rect 1040 -2470 1060 -2450
rect 1080 -2470 1100 -2450
rect 1120 -2470 1140 -2450
rect 1160 -2470 1180 -2450
rect 1200 -2470 1220 -2450
rect 1240 -2470 1260 -2450
rect 1280 -2470 1300 -2450
rect 1320 -2470 1340 -2450
rect 1360 -2470 1380 -2450
rect 1400 -2470 1420 -2450
rect 1440 -2470 1460 -2450
rect -60 -2520 -40 -2495
rect -20 -2520 0 -2495
rect 20 -2520 40 -2495
rect 60 -2520 80 -2495
rect 1760 -2565 1780 -2545
rect 1800 -2565 1820 -2545
rect 1840 -2565 1860 -2545
rect 1880 -2565 1900 -2545
rect 1920 -2565 1940 -2545
rect 1960 -2565 1980 -2545
rect 2000 -2565 2020 -2545
rect 2040 -2565 2060 -2545
rect 2080 -2565 2100 -2545
rect 2120 -2565 2140 -2545
rect 2160 -2565 2180 -2545
rect 2200 -2565 2220 -2545
rect 2240 -2565 2260 -2545
rect 2280 -2565 2300 -2545
rect 2320 -2565 2340 -2545
rect 2360 -2565 2380 -2545
rect 2400 -2565 2420 -2545
rect 2440 -2565 2460 -2545
rect 2480 -2565 2500 -2545
rect 2520 -2565 2540 -2545
rect -60 -2615 -40 -2590
rect -20 -2615 0 -2590
rect 20 -2615 40 -2590
rect 60 -2615 80 -2590
rect 680 -2660 700 -2640
rect 720 -2660 740 -2640
rect 760 -2660 780 -2640
rect 800 -2660 820 -2640
rect 840 -2660 860 -2640
rect 880 -2660 900 -2640
rect 920 -2660 940 -2640
rect 960 -2660 980 -2640
rect 1000 -2660 1020 -2640
rect 1040 -2660 1060 -2640
rect 1080 -2660 1100 -2640
rect 1120 -2660 1140 -2640
rect 1160 -2660 1180 -2640
rect 1200 -2660 1220 -2640
rect 1240 -2660 1260 -2640
rect 1280 -2660 1300 -2640
rect 1320 -2660 1340 -2640
rect 1360 -2660 1380 -2640
rect 1400 -2660 1420 -2640
rect 1440 -2660 1460 -2640
rect -60 -2710 -40 -2685
rect -20 -2710 0 -2685
rect 20 -2710 40 -2685
rect 60 -2710 80 -2685
rect 1760 -2755 1780 -2735
rect 1800 -2755 1820 -2735
rect 1840 -2755 1860 -2735
rect 1880 -2755 1900 -2735
rect 1920 -2755 1940 -2735
rect 1960 -2755 1980 -2735
rect 2000 -2755 2020 -2735
rect 2040 -2755 2060 -2735
rect 2080 -2755 2100 -2735
rect 2120 -2755 2140 -2735
rect 2160 -2755 2180 -2735
rect 2200 -2755 2220 -2735
rect 2240 -2755 2260 -2735
rect 2280 -2755 2300 -2735
rect 2320 -2755 2340 -2735
rect 2360 -2755 2380 -2735
rect 2400 -2755 2420 -2735
rect 2440 -2755 2460 -2735
rect 2480 -2755 2500 -2735
rect 2520 -2755 2540 -2735
rect 1760 -2795 1780 -2775
rect 1800 -2795 1820 -2775
rect 1840 -2795 1860 -2775
rect 1880 -2795 1900 -2775
rect 1920 -2795 1940 -2775
rect 1960 -2795 1980 -2775
rect 2000 -2795 2020 -2775
rect 2040 -2795 2060 -2775
rect 2080 -2795 2100 -2775
rect 2120 -2795 2140 -2775
rect 2160 -2795 2180 -2775
rect 2200 -2795 2220 -2775
rect 2240 -2795 2260 -2775
rect 2280 -2795 2300 -2775
rect 2320 -2795 2340 -2775
rect 2360 -2795 2380 -2775
rect 2400 -2795 2420 -2775
rect 2440 -2795 2460 -2775
rect 2480 -2795 2500 -2775
rect 2520 -2795 2540 -2775
<< metal1 >>
rect 670 2260 1470 2270
rect 670 2240 680 2260
rect 700 2240 720 2260
rect 740 2240 760 2260
rect 780 2240 800 2260
rect 820 2240 840 2260
rect 860 2240 880 2260
rect 900 2240 920 2260
rect 940 2240 960 2260
rect 980 2240 1000 2260
rect 1020 2240 1040 2260
rect 1060 2240 1080 2260
rect 1100 2240 1120 2260
rect 1140 2240 1160 2260
rect 1180 2240 1200 2260
rect 1220 2240 1240 2260
rect 1260 2240 1280 2260
rect 1300 2240 1320 2260
rect 1340 2240 1360 2260
rect 1380 2240 1400 2260
rect 1420 2240 1440 2260
rect 1460 2240 1470 2260
rect 670 2217 1470 2240
rect 670 2197 680 2217
rect 700 2197 720 2217
rect 740 2197 760 2217
rect 780 2197 800 2217
rect 820 2197 840 2217
rect 860 2197 880 2217
rect 900 2197 920 2217
rect 940 2197 960 2217
rect 980 2197 1000 2217
rect 1020 2197 1040 2217
rect 1060 2197 1080 2217
rect 1100 2197 1120 2217
rect 1140 2197 1160 2217
rect 1180 2197 1200 2217
rect 1220 2197 1240 2217
rect 1260 2197 1280 2217
rect 1300 2197 1320 2217
rect 1340 2197 1360 2217
rect 1380 2197 1400 2217
rect 1420 2197 1440 2217
rect 1460 2197 1470 2217
rect 0 2175 165 2185
rect 0 2155 10 2175
rect 30 2155 50 2175
rect 70 2155 90 2175
rect 110 2155 130 2175
rect 150 2155 165 2175
rect 0 2095 165 2155
rect 0 2075 10 2095
rect 30 2075 50 2095
rect 70 2075 90 2095
rect 110 2075 130 2095
rect 150 2075 165 2095
rect 0 2010 165 2075
rect 0 1990 10 2010
rect 30 1990 50 2010
rect 70 1990 90 2010
rect 110 1990 130 2010
rect 150 1990 165 2010
rect 0 1930 165 1990
rect 0 1910 10 1930
rect 30 1910 50 1930
rect 70 1910 90 1930
rect 110 1910 130 1930
rect 150 1910 165 1930
rect 0 1850 165 1910
rect 0 1830 10 1850
rect 30 1830 50 1850
rect 70 1830 90 1850
rect 110 1830 130 1850
rect 150 1830 165 1850
rect 0 1765 165 1830
rect 0 1745 10 1765
rect 30 1745 50 1765
rect 70 1745 90 1765
rect 110 1745 130 1765
rect 150 1745 165 1765
rect 0 1685 165 1745
rect 0 1665 10 1685
rect 30 1665 50 1685
rect 70 1665 90 1685
rect 110 1665 130 1685
rect 150 1665 165 1685
rect 0 1600 165 1665
rect 0 1580 10 1600
rect 30 1580 50 1600
rect 70 1580 90 1600
rect 110 1580 130 1600
rect 150 1580 165 1600
rect 0 1520 165 1580
rect 0 1500 10 1520
rect 30 1500 50 1520
rect 70 1500 90 1520
rect 110 1500 130 1520
rect 150 1500 165 1520
rect 0 1440 165 1500
rect 0 1420 10 1440
rect 30 1420 50 1440
rect 70 1420 90 1440
rect 110 1420 130 1440
rect 150 1420 165 1440
rect 0 1355 165 1420
rect 0 1335 10 1355
rect 30 1335 50 1355
rect 70 1335 90 1355
rect 110 1335 130 1355
rect 150 1335 165 1355
rect 0 1275 165 1335
rect 0 1255 10 1275
rect 30 1255 50 1275
rect 70 1255 90 1275
rect 110 1255 130 1275
rect 150 1255 165 1275
rect 0 1190 165 1255
rect 0 1170 10 1190
rect 30 1170 50 1190
rect 70 1170 90 1190
rect 110 1170 130 1190
rect 150 1170 165 1190
rect 0 1110 165 1170
rect 0 1090 10 1110
rect 30 1090 50 1110
rect 70 1090 90 1110
rect 110 1090 130 1110
rect 150 1090 165 1110
rect 0 1030 165 1090
rect 0 1010 10 1030
rect 30 1010 50 1030
rect 70 1010 90 1030
rect 110 1010 130 1030
rect 150 1010 165 1030
rect 0 945 165 1010
rect 0 925 10 945
rect 30 925 50 945
rect 70 925 90 945
rect 110 925 130 945
rect 150 925 165 945
rect 0 865 165 925
rect 0 845 10 865
rect 30 845 50 865
rect 70 845 90 865
rect 110 845 130 865
rect 150 845 165 865
rect 0 780 165 845
rect 0 760 10 780
rect 30 760 50 780
rect 70 760 90 780
rect 110 760 130 780
rect 150 760 165 780
rect 0 700 165 760
rect 0 680 10 700
rect 30 680 50 700
rect 70 680 90 700
rect 110 680 130 700
rect 150 680 165 700
rect 0 620 165 680
rect 0 600 10 620
rect 30 600 50 620
rect 70 600 90 620
rect 110 600 130 620
rect 150 600 165 620
rect 0 535 165 600
rect 0 515 10 535
rect 30 515 50 535
rect 70 515 90 535
rect 110 515 130 535
rect 150 515 165 535
rect 0 455 165 515
rect 0 435 10 455
rect 30 435 50 455
rect 70 435 90 455
rect 110 435 130 455
rect 150 435 165 455
rect 0 375 165 435
rect 0 355 10 375
rect 30 355 50 375
rect 70 355 90 375
rect 110 355 130 375
rect 150 355 165 375
rect 0 290 165 355
rect 0 270 10 290
rect 30 270 50 290
rect 70 270 90 290
rect 110 270 130 290
rect 150 270 165 290
rect 0 210 165 270
rect 0 190 10 210
rect 30 190 50 210
rect 70 190 90 210
rect 110 190 130 210
rect 150 190 165 210
rect 0 130 165 190
rect 0 110 10 130
rect 30 110 50 130
rect 70 110 90 130
rect 110 110 130 130
rect 150 110 165 130
rect 0 100 165 110
rect 670 2053 1470 2197
rect 670 2033 680 2053
rect 700 2033 720 2053
rect 740 2033 760 2053
rect 780 2033 800 2053
rect 820 2033 840 2053
rect 860 2033 880 2053
rect 900 2033 920 2053
rect 940 2033 960 2053
rect 980 2033 1000 2053
rect 1020 2033 1040 2053
rect 1060 2033 1080 2053
rect 1100 2033 1120 2053
rect 1140 2033 1160 2053
rect 1180 2033 1200 2053
rect 1220 2033 1240 2053
rect 1260 2033 1280 2053
rect 1300 2033 1320 2053
rect 1340 2033 1360 2053
rect 1380 2033 1400 2053
rect 1420 2033 1440 2053
rect 1460 2033 1470 2053
rect 670 1889 1470 2033
rect 670 1869 680 1889
rect 700 1869 720 1889
rect 740 1869 760 1889
rect 780 1869 800 1889
rect 820 1869 840 1889
rect 860 1869 880 1889
rect 900 1869 920 1889
rect 940 1869 960 1889
rect 980 1869 1000 1889
rect 1020 1869 1040 1889
rect 1060 1869 1080 1889
rect 1100 1869 1120 1889
rect 1140 1869 1160 1889
rect 1180 1869 1200 1889
rect 1220 1869 1240 1889
rect 1260 1869 1280 1889
rect 1300 1869 1320 1889
rect 1340 1869 1360 1889
rect 1380 1869 1400 1889
rect 1420 1869 1440 1889
rect 1460 1869 1470 1889
rect 670 1725 1470 1869
rect 670 1705 680 1725
rect 700 1705 720 1725
rect 740 1705 760 1725
rect 780 1705 800 1725
rect 820 1705 840 1725
rect 860 1705 880 1725
rect 900 1705 920 1725
rect 940 1705 960 1725
rect 980 1705 1000 1725
rect 1020 1705 1040 1725
rect 1060 1705 1080 1725
rect 1100 1705 1120 1725
rect 1140 1705 1160 1725
rect 1180 1705 1200 1725
rect 1220 1705 1240 1725
rect 1260 1705 1280 1725
rect 1300 1705 1320 1725
rect 1340 1705 1360 1725
rect 1380 1705 1400 1725
rect 1420 1705 1440 1725
rect 1460 1705 1470 1725
rect 670 1561 1470 1705
rect 670 1541 680 1561
rect 700 1541 720 1561
rect 740 1541 760 1561
rect 780 1541 800 1561
rect 820 1541 840 1561
rect 860 1541 880 1561
rect 900 1541 920 1561
rect 940 1541 960 1561
rect 980 1541 1000 1561
rect 1020 1541 1040 1561
rect 1060 1541 1080 1561
rect 1100 1541 1120 1561
rect 1140 1541 1160 1561
rect 1180 1541 1200 1561
rect 1220 1541 1240 1561
rect 1260 1541 1280 1561
rect 1300 1541 1320 1561
rect 1340 1541 1360 1561
rect 1380 1541 1400 1561
rect 1420 1541 1440 1561
rect 1460 1541 1470 1561
rect 670 1397 1470 1541
rect 670 1377 680 1397
rect 700 1377 720 1397
rect 740 1377 760 1397
rect 780 1377 800 1397
rect 820 1377 840 1397
rect 860 1377 880 1397
rect 900 1377 920 1397
rect 940 1377 960 1397
rect 980 1377 1000 1397
rect 1020 1377 1040 1397
rect 1060 1377 1080 1397
rect 1100 1377 1120 1397
rect 1140 1377 1160 1397
rect 1180 1377 1200 1397
rect 1220 1377 1240 1397
rect 1260 1377 1280 1397
rect 1300 1377 1320 1397
rect 1340 1377 1360 1397
rect 1380 1377 1400 1397
rect 1420 1377 1440 1397
rect 1460 1377 1470 1397
rect 670 1233 1470 1377
rect 670 1213 680 1233
rect 700 1213 720 1233
rect 740 1213 760 1233
rect 780 1213 800 1233
rect 820 1213 840 1233
rect 860 1213 880 1233
rect 900 1213 920 1233
rect 940 1213 960 1233
rect 980 1213 1000 1233
rect 1020 1213 1040 1233
rect 1060 1213 1080 1233
rect 1100 1213 1120 1233
rect 1140 1213 1160 1233
rect 1180 1213 1200 1233
rect 1220 1213 1240 1233
rect 1260 1213 1280 1233
rect 1300 1213 1320 1233
rect 1340 1213 1360 1233
rect 1380 1213 1400 1233
rect 1420 1213 1440 1233
rect 1460 1213 1470 1233
rect 670 1069 1470 1213
rect 670 1049 680 1069
rect 700 1049 720 1069
rect 740 1049 760 1069
rect 780 1049 800 1069
rect 820 1049 840 1069
rect 860 1049 880 1069
rect 900 1049 920 1069
rect 940 1049 960 1069
rect 980 1049 1000 1069
rect 1020 1049 1040 1069
rect 1060 1049 1080 1069
rect 1100 1049 1120 1069
rect 1140 1049 1160 1069
rect 1180 1049 1200 1069
rect 1220 1049 1240 1069
rect 1260 1049 1280 1069
rect 1300 1049 1320 1069
rect 1340 1049 1360 1069
rect 1380 1049 1400 1069
rect 1420 1049 1440 1069
rect 1460 1049 1470 1069
rect 670 905 1470 1049
rect 670 885 680 905
rect 700 885 720 905
rect 740 885 760 905
rect 780 885 800 905
rect 820 885 840 905
rect 860 885 880 905
rect 900 885 920 905
rect 940 885 960 905
rect 980 885 1000 905
rect 1020 885 1040 905
rect 1060 885 1080 905
rect 1100 885 1120 905
rect 1140 885 1160 905
rect 1180 885 1200 905
rect 1220 885 1240 905
rect 1260 885 1280 905
rect 1300 885 1320 905
rect 1340 885 1360 905
rect 1380 885 1400 905
rect 1420 885 1440 905
rect 1460 885 1470 905
rect 670 741 1470 885
rect 670 721 680 741
rect 700 721 720 741
rect 740 721 760 741
rect 780 721 800 741
rect 820 721 840 741
rect 860 721 880 741
rect 900 721 920 741
rect 940 721 960 741
rect 980 721 1000 741
rect 1020 721 1040 741
rect 1060 721 1080 741
rect 1100 721 1120 741
rect 1140 721 1160 741
rect 1180 721 1200 741
rect 1220 721 1240 741
rect 1260 721 1280 741
rect 1300 721 1320 741
rect 1340 721 1360 741
rect 1380 721 1400 741
rect 1420 721 1440 741
rect 1460 721 1470 741
rect 670 577 1470 721
rect 670 557 680 577
rect 700 557 720 577
rect 740 557 760 577
rect 780 557 800 577
rect 820 557 840 577
rect 860 557 880 577
rect 900 557 920 577
rect 940 557 960 577
rect 980 557 1000 577
rect 1020 557 1040 577
rect 1060 557 1080 577
rect 1100 557 1120 577
rect 1140 557 1160 577
rect 1180 557 1200 577
rect 1220 557 1240 577
rect 1260 557 1280 577
rect 1300 557 1320 577
rect 1340 557 1360 577
rect 1380 557 1400 577
rect 1420 557 1440 577
rect 1460 557 1470 577
rect 670 413 1470 557
rect 670 393 680 413
rect 700 393 720 413
rect 740 393 760 413
rect 780 393 800 413
rect 820 393 840 413
rect 860 393 880 413
rect 900 393 920 413
rect 940 393 960 413
rect 980 393 1000 413
rect 1020 393 1040 413
rect 1060 393 1080 413
rect 1100 393 1120 413
rect 1140 393 1160 413
rect 1180 393 1200 413
rect 1220 393 1240 413
rect 1260 393 1280 413
rect 1300 393 1320 413
rect 1340 393 1360 413
rect 1380 393 1400 413
rect 1420 393 1440 413
rect 1460 393 1470 413
rect 670 249 1470 393
rect 670 229 680 249
rect 700 229 720 249
rect 740 229 760 249
rect 780 229 800 249
rect 820 229 840 249
rect 860 229 880 249
rect 900 229 920 249
rect 940 229 960 249
rect 980 229 1000 249
rect 1020 229 1040 249
rect 1060 229 1080 249
rect 1100 229 1120 249
rect 1140 229 1160 249
rect 1180 229 1200 249
rect 1220 229 1240 249
rect 1260 229 1280 249
rect 1300 229 1320 249
rect 1340 229 1360 249
rect 1380 229 1400 249
rect 1420 229 1440 249
rect 1460 229 1470 249
rect 670 85 1470 229
rect 670 65 680 85
rect 700 65 720 85
rect 740 65 760 85
rect 780 65 800 85
rect 820 65 840 85
rect 860 65 880 85
rect 900 65 920 85
rect 940 65 960 85
rect 980 65 1000 85
rect 1020 65 1040 85
rect 1060 65 1080 85
rect 1100 65 1120 85
rect 1140 65 1160 85
rect 1180 65 1200 85
rect 1220 65 1240 85
rect 1260 65 1280 85
rect 1300 65 1320 85
rect 1340 65 1360 85
rect 1380 65 1400 85
rect 1420 65 1440 85
rect 1460 65 1470 85
rect 670 45 1470 65
rect 670 25 680 45
rect 700 25 720 45
rect 740 25 760 45
rect 780 25 800 45
rect 820 25 840 45
rect 860 25 880 45
rect 900 25 920 45
rect 940 25 960 45
rect 980 25 1000 45
rect 1020 25 1040 45
rect 1060 25 1080 45
rect 1100 25 1120 45
rect 1140 25 1160 45
rect 1180 25 1200 45
rect 1220 25 1240 45
rect 1260 25 1280 45
rect 1300 25 1320 45
rect 1340 25 1360 45
rect 1380 25 1400 45
rect 1420 25 1440 45
rect 1460 25 1470 45
rect -70 -310 85 -300
rect -70 -335 -60 -310
rect -40 -335 -20 -310
rect 0 -335 20 -310
rect 40 -335 60 -310
rect 80 -335 85 -310
rect -70 -405 85 -335
rect -70 -430 -60 -405
rect -40 -430 -20 -405
rect 0 -430 20 -405
rect 40 -430 60 -405
rect 80 -430 85 -405
rect -70 -500 85 -430
rect -70 -525 -60 -500
rect -40 -525 -20 -500
rect 0 -525 20 -500
rect 40 -525 60 -500
rect 80 -525 85 -500
rect -70 -595 85 -525
rect -70 -620 -60 -595
rect -40 -620 -20 -595
rect 0 -620 20 -595
rect 40 -620 60 -595
rect 80 -620 85 -595
rect -70 -690 85 -620
rect -70 -715 -60 -690
rect -40 -715 -20 -690
rect 0 -715 20 -690
rect 40 -715 60 -690
rect 80 -715 85 -690
rect -70 -785 85 -715
rect -70 -810 -60 -785
rect -40 -810 -20 -785
rect 0 -810 20 -785
rect 40 -810 60 -785
rect 80 -810 85 -785
rect -70 -880 85 -810
rect -70 -905 -60 -880
rect -40 -905 -20 -880
rect 0 -905 20 -880
rect 40 -905 60 -880
rect 80 -905 85 -880
rect -70 -975 85 -905
rect -70 -1000 -60 -975
rect -40 -1000 -20 -975
rect 0 -1000 20 -975
rect 40 -1000 60 -975
rect 80 -1000 85 -975
rect -70 -1070 85 -1000
rect -70 -1095 -60 -1070
rect -40 -1095 -20 -1070
rect 0 -1095 20 -1070
rect 40 -1095 60 -1070
rect 80 -1095 85 -1070
rect -70 -1165 85 -1095
rect -70 -1190 -60 -1165
rect -40 -1190 -20 -1165
rect 0 -1190 20 -1165
rect 40 -1190 60 -1165
rect 80 -1190 85 -1165
rect -70 -1260 85 -1190
rect -70 -1285 -60 -1260
rect -40 -1285 -20 -1260
rect 0 -1285 20 -1260
rect 40 -1285 60 -1260
rect 80 -1285 85 -1260
rect -70 -1355 85 -1285
rect -70 -1380 -60 -1355
rect -40 -1380 -20 -1355
rect 0 -1380 20 -1355
rect 40 -1380 60 -1355
rect 80 -1380 85 -1355
rect -70 -1450 85 -1380
rect -70 -1475 -60 -1450
rect -40 -1475 -20 -1450
rect 0 -1475 20 -1450
rect 40 -1475 60 -1450
rect 80 -1475 85 -1450
rect -70 -1545 85 -1475
rect -70 -1570 -60 -1545
rect -40 -1570 -20 -1545
rect 0 -1570 20 -1545
rect 40 -1570 60 -1545
rect 80 -1570 85 -1545
rect -70 -1640 85 -1570
rect -70 -1665 -60 -1640
rect -40 -1665 -20 -1640
rect 0 -1665 20 -1640
rect 40 -1665 60 -1640
rect 80 -1665 85 -1640
rect -70 -1735 85 -1665
rect -70 -1760 -60 -1735
rect -40 -1760 -20 -1735
rect 0 -1760 20 -1735
rect 40 -1760 60 -1735
rect 80 -1760 85 -1735
rect -70 -1830 85 -1760
rect -70 -1855 -60 -1830
rect -40 -1855 -20 -1830
rect 0 -1855 20 -1830
rect 40 -1855 60 -1830
rect 80 -1855 85 -1830
rect -70 -1925 85 -1855
rect -70 -1950 -60 -1925
rect -40 -1950 -20 -1925
rect 0 -1950 20 -1925
rect 40 -1950 60 -1925
rect 80 -1950 85 -1925
rect -70 -2020 85 -1950
rect -70 -2045 -60 -2020
rect -40 -2045 -20 -2020
rect 0 -2045 20 -2020
rect 40 -2045 60 -2020
rect 80 -2045 85 -2020
rect -70 -2115 85 -2045
rect -70 -2140 -60 -2115
rect -40 -2140 -20 -2115
rect 0 -2140 20 -2115
rect 40 -2140 60 -2115
rect 80 -2140 85 -2115
rect -70 -2210 85 -2140
rect -70 -2235 -60 -2210
rect -40 -2235 -20 -2210
rect 0 -2235 20 -2210
rect 40 -2235 60 -2210
rect 80 -2235 85 -2210
rect -70 -2305 85 -2235
rect -70 -2330 -60 -2305
rect -40 -2330 -20 -2305
rect 0 -2330 20 -2305
rect 40 -2330 60 -2305
rect 80 -2330 85 -2305
rect -70 -2400 85 -2330
rect -70 -2425 -60 -2400
rect -40 -2425 -20 -2400
rect 0 -2425 20 -2400
rect 40 -2425 60 -2400
rect 80 -2425 85 -2400
rect -70 -2495 85 -2425
rect -70 -2520 -60 -2495
rect -40 -2520 -20 -2495
rect 0 -2520 20 -2495
rect 40 -2520 60 -2495
rect 80 -2520 85 -2495
rect -70 -2590 85 -2520
rect -70 -2615 -60 -2590
rect -40 -2615 -20 -2590
rect 0 -2615 20 -2590
rect 40 -2615 60 -2590
rect 80 -2615 85 -2590
rect -70 -2685 85 -2615
rect 670 -360 1470 25
rect 1750 2135 2550 2385
rect 1750 2115 1760 2135
rect 1780 2115 1800 2135
rect 1820 2115 1840 2135
rect 1860 2115 1880 2135
rect 1900 2115 1920 2135
rect 1940 2115 1960 2135
rect 1980 2115 2000 2135
rect 2020 2115 2040 2135
rect 2060 2115 2080 2135
rect 2100 2115 2120 2135
rect 2140 2115 2160 2135
rect 2180 2115 2200 2135
rect 2220 2115 2240 2135
rect 2260 2115 2280 2135
rect 2300 2115 2320 2135
rect 2340 2115 2360 2135
rect 2380 2115 2400 2135
rect 2420 2115 2440 2135
rect 2460 2115 2480 2135
rect 2500 2115 2520 2135
rect 2540 2115 2550 2135
rect 1750 1971 2550 2115
rect 1750 1951 1760 1971
rect 1780 1951 1800 1971
rect 1820 1951 1840 1971
rect 1860 1951 1880 1971
rect 1900 1951 1920 1971
rect 1940 1951 1960 1971
rect 1980 1951 2000 1971
rect 2020 1951 2040 1971
rect 2060 1951 2080 1971
rect 2100 1951 2120 1971
rect 2140 1951 2160 1971
rect 2180 1951 2200 1971
rect 2220 1951 2240 1971
rect 2260 1951 2280 1971
rect 2300 1951 2320 1971
rect 2340 1951 2360 1971
rect 2380 1951 2400 1971
rect 2420 1951 2440 1971
rect 2460 1951 2480 1971
rect 2500 1951 2520 1971
rect 2540 1951 2550 1971
rect 1750 1807 2550 1951
rect 1750 1787 1760 1807
rect 1780 1787 1800 1807
rect 1820 1787 1840 1807
rect 1860 1787 1880 1807
rect 1900 1787 1920 1807
rect 1940 1787 1960 1807
rect 1980 1787 2000 1807
rect 2020 1787 2040 1807
rect 2060 1787 2080 1807
rect 2100 1787 2120 1807
rect 2140 1787 2160 1807
rect 2180 1787 2200 1807
rect 2220 1787 2240 1807
rect 2260 1787 2280 1807
rect 2300 1787 2320 1807
rect 2340 1787 2360 1807
rect 2380 1787 2400 1807
rect 2420 1787 2440 1807
rect 2460 1787 2480 1807
rect 2500 1787 2520 1807
rect 2540 1787 2550 1807
rect 1750 1643 2550 1787
rect 1750 1623 1760 1643
rect 1780 1623 1800 1643
rect 1820 1623 1840 1643
rect 1860 1623 1880 1643
rect 1900 1623 1920 1643
rect 1940 1623 1960 1643
rect 1980 1623 2000 1643
rect 2020 1623 2040 1643
rect 2060 1623 2080 1643
rect 2100 1623 2120 1643
rect 2140 1623 2160 1643
rect 2180 1623 2200 1643
rect 2220 1623 2240 1643
rect 2260 1623 2280 1643
rect 2300 1623 2320 1643
rect 2340 1623 2360 1643
rect 2380 1623 2400 1643
rect 2420 1623 2440 1643
rect 2460 1623 2480 1643
rect 2500 1623 2520 1643
rect 2540 1623 2550 1643
rect 1750 1479 2550 1623
rect 1750 1459 1760 1479
rect 1780 1459 1800 1479
rect 1820 1459 1840 1479
rect 1860 1459 1880 1479
rect 1900 1459 1920 1479
rect 1940 1459 1960 1479
rect 1980 1459 2000 1479
rect 2020 1459 2040 1479
rect 2060 1459 2080 1479
rect 2100 1459 2120 1479
rect 2140 1459 2160 1479
rect 2180 1459 2200 1479
rect 2220 1459 2240 1479
rect 2260 1459 2280 1479
rect 2300 1459 2320 1479
rect 2340 1459 2360 1479
rect 2380 1459 2400 1479
rect 2420 1459 2440 1479
rect 2460 1459 2480 1479
rect 2500 1459 2520 1479
rect 2540 1459 2550 1479
rect 1750 1315 2550 1459
rect 1750 1295 1760 1315
rect 1780 1295 1800 1315
rect 1820 1295 1840 1315
rect 1860 1295 1880 1315
rect 1900 1295 1920 1315
rect 1940 1295 1960 1315
rect 1980 1295 2000 1315
rect 2020 1295 2040 1315
rect 2060 1295 2080 1315
rect 2100 1295 2120 1315
rect 2140 1295 2160 1315
rect 2180 1295 2200 1315
rect 2220 1295 2240 1315
rect 2260 1295 2280 1315
rect 2300 1295 2320 1315
rect 2340 1295 2360 1315
rect 2380 1295 2400 1315
rect 2420 1295 2440 1315
rect 2460 1295 2480 1315
rect 2500 1295 2520 1315
rect 2540 1295 2550 1315
rect 1750 1151 2550 1295
rect 1750 1131 1760 1151
rect 1780 1131 1800 1151
rect 1820 1131 1840 1151
rect 1860 1131 1880 1151
rect 1900 1131 1920 1151
rect 1940 1131 1960 1151
rect 1980 1131 2000 1151
rect 2020 1131 2040 1151
rect 2060 1131 2080 1151
rect 2100 1131 2120 1151
rect 2140 1131 2160 1151
rect 2180 1131 2200 1151
rect 2220 1131 2240 1151
rect 2260 1131 2280 1151
rect 2300 1131 2320 1151
rect 2340 1131 2360 1151
rect 2380 1131 2400 1151
rect 2420 1131 2440 1151
rect 2460 1131 2480 1151
rect 2500 1131 2520 1151
rect 2540 1131 2550 1151
rect 1750 987 2550 1131
rect 1750 967 1760 987
rect 1780 967 1800 987
rect 1820 967 1840 987
rect 1860 967 1880 987
rect 1900 967 1920 987
rect 1940 967 1960 987
rect 1980 967 2000 987
rect 2020 967 2040 987
rect 2060 967 2080 987
rect 2100 967 2120 987
rect 2140 967 2160 987
rect 2180 967 2200 987
rect 2220 967 2240 987
rect 2260 967 2280 987
rect 2300 967 2320 987
rect 2340 967 2360 987
rect 2380 967 2400 987
rect 2420 967 2440 987
rect 2460 967 2480 987
rect 2500 967 2520 987
rect 2540 967 2550 987
rect 1750 823 2550 967
rect 1750 803 1760 823
rect 1780 803 1800 823
rect 1820 803 1840 823
rect 1860 803 1880 823
rect 1900 803 1920 823
rect 1940 803 1960 823
rect 1980 803 2000 823
rect 2020 803 2040 823
rect 2060 803 2080 823
rect 2100 803 2120 823
rect 2140 803 2160 823
rect 2180 803 2200 823
rect 2220 803 2240 823
rect 2260 803 2280 823
rect 2300 803 2320 823
rect 2340 803 2360 823
rect 2380 803 2400 823
rect 2420 803 2440 823
rect 2460 803 2480 823
rect 2500 803 2520 823
rect 2540 803 2550 823
rect 1750 659 2550 803
rect 1750 639 1760 659
rect 1780 639 1800 659
rect 1820 639 1840 659
rect 1860 639 1880 659
rect 1900 639 1920 659
rect 1940 639 1960 659
rect 1980 639 2000 659
rect 2020 639 2040 659
rect 2060 639 2080 659
rect 2100 639 2120 659
rect 2140 639 2160 659
rect 2180 639 2200 659
rect 2220 639 2240 659
rect 2260 639 2280 659
rect 2300 639 2320 659
rect 2340 639 2360 659
rect 2380 639 2400 659
rect 2420 639 2440 659
rect 2460 639 2480 659
rect 2500 639 2520 659
rect 2540 639 2550 659
rect 1750 495 2550 639
rect 1750 475 1760 495
rect 1780 475 1800 495
rect 1820 475 1840 495
rect 1860 475 1880 495
rect 1900 475 1920 495
rect 1940 475 1960 495
rect 1980 475 2000 495
rect 2020 475 2040 495
rect 2060 475 2080 495
rect 2100 475 2120 495
rect 2140 475 2160 495
rect 2180 475 2200 495
rect 2220 475 2240 495
rect 2260 475 2280 495
rect 2300 475 2320 495
rect 2340 475 2360 495
rect 2380 475 2400 495
rect 2420 475 2440 495
rect 2460 475 2480 495
rect 2500 475 2520 495
rect 2540 475 2550 495
rect 1750 331 2550 475
rect 1750 311 1760 331
rect 1780 311 1800 331
rect 1820 311 1840 331
rect 1860 311 1880 331
rect 1900 311 1920 331
rect 1940 311 1960 331
rect 1980 311 2000 331
rect 2020 311 2040 331
rect 2060 311 2080 331
rect 2100 311 2120 331
rect 2140 311 2160 331
rect 2180 311 2200 331
rect 2220 311 2240 331
rect 2260 311 2280 331
rect 2300 311 2320 331
rect 2340 311 2360 331
rect 2380 311 2400 331
rect 2420 311 2440 331
rect 2460 311 2480 331
rect 2500 311 2520 331
rect 2540 311 2550 331
rect 1750 167 2550 311
rect 1750 147 1760 167
rect 1780 147 1800 167
rect 1820 147 1840 167
rect 1860 147 1880 167
rect 1900 147 1920 167
rect 1940 147 1960 167
rect 1980 147 2000 167
rect 2020 147 2040 167
rect 2060 147 2080 167
rect 2100 147 2120 167
rect 2140 147 2160 167
rect 2180 147 2200 167
rect 2220 147 2240 167
rect 2260 147 2280 167
rect 2300 147 2320 167
rect 2340 147 2360 167
rect 2380 147 2400 167
rect 2420 147 2440 167
rect 2460 147 2480 167
rect 2500 147 2520 167
rect 2540 147 2550 167
rect 1750 15 2550 147
rect 670 -380 680 -360
rect 700 -380 720 -360
rect 740 -380 760 -360
rect 780 -380 800 -360
rect 820 -380 840 -360
rect 860 -380 880 -360
rect 900 -380 920 -360
rect 940 -380 960 -360
rect 980 -380 1000 -360
rect 1020 -380 1040 -360
rect 1060 -380 1080 -360
rect 1100 -380 1120 -360
rect 1140 -380 1160 -360
rect 1180 -380 1200 -360
rect 1220 -380 1240 -360
rect 1260 -380 1280 -360
rect 1300 -380 1320 -360
rect 1340 -380 1360 -360
rect 1380 -380 1400 -360
rect 1420 -380 1440 -360
rect 1460 -380 1470 -360
rect 670 -550 1470 -380
rect 670 -570 680 -550
rect 700 -570 720 -550
rect 740 -570 760 -550
rect 780 -570 800 -550
rect 820 -570 840 -550
rect 860 -570 880 -550
rect 900 -570 920 -550
rect 940 -570 960 -550
rect 980 -570 1000 -550
rect 1020 -570 1040 -550
rect 1060 -570 1080 -550
rect 1100 -570 1120 -550
rect 1140 -570 1160 -550
rect 1180 -570 1200 -550
rect 1220 -570 1240 -550
rect 1260 -570 1280 -550
rect 1300 -570 1320 -550
rect 1340 -570 1360 -550
rect 1380 -570 1400 -550
rect 1420 -570 1440 -550
rect 1460 -570 1470 -550
rect 670 -740 1470 -570
rect 670 -760 680 -740
rect 700 -760 720 -740
rect 740 -760 760 -740
rect 780 -760 800 -740
rect 820 -760 840 -740
rect 860 -760 880 -740
rect 900 -760 920 -740
rect 940 -760 960 -740
rect 980 -760 1000 -740
rect 1020 -760 1040 -740
rect 1060 -760 1080 -740
rect 1100 -760 1120 -740
rect 1140 -760 1160 -740
rect 1180 -760 1200 -740
rect 1220 -760 1240 -740
rect 1260 -760 1280 -740
rect 1300 -760 1320 -740
rect 1340 -760 1360 -740
rect 1380 -760 1400 -740
rect 1420 -760 1440 -740
rect 1460 -760 1470 -740
rect 670 -930 1470 -760
rect 670 -950 680 -930
rect 700 -950 720 -930
rect 740 -950 760 -930
rect 780 -950 800 -930
rect 820 -950 840 -930
rect 860 -950 880 -930
rect 900 -950 920 -930
rect 940 -950 960 -930
rect 980 -950 1000 -930
rect 1020 -950 1040 -930
rect 1060 -950 1080 -930
rect 1100 -950 1120 -930
rect 1140 -950 1160 -930
rect 1180 -950 1200 -930
rect 1220 -950 1240 -930
rect 1260 -950 1280 -930
rect 1300 -950 1320 -930
rect 1340 -950 1360 -930
rect 1380 -950 1400 -930
rect 1420 -950 1440 -930
rect 1460 -950 1470 -930
rect 670 -1120 1470 -950
rect 670 -1140 680 -1120
rect 700 -1140 720 -1120
rect 740 -1140 760 -1120
rect 780 -1140 800 -1120
rect 820 -1140 840 -1120
rect 860 -1140 880 -1120
rect 900 -1140 920 -1120
rect 940 -1140 960 -1120
rect 980 -1140 1000 -1120
rect 1020 -1140 1040 -1120
rect 1060 -1140 1080 -1120
rect 1100 -1140 1120 -1120
rect 1140 -1140 1160 -1120
rect 1180 -1140 1200 -1120
rect 1220 -1140 1240 -1120
rect 1260 -1140 1280 -1120
rect 1300 -1140 1320 -1120
rect 1340 -1140 1360 -1120
rect 1380 -1140 1400 -1120
rect 1420 -1140 1440 -1120
rect 1460 -1140 1470 -1120
rect 670 -1310 1470 -1140
rect 670 -1330 680 -1310
rect 700 -1330 720 -1310
rect 740 -1330 760 -1310
rect 780 -1330 800 -1310
rect 820 -1330 840 -1310
rect 860 -1330 880 -1310
rect 900 -1330 920 -1310
rect 940 -1330 960 -1310
rect 980 -1330 1000 -1310
rect 1020 -1330 1040 -1310
rect 1060 -1330 1080 -1310
rect 1100 -1330 1120 -1310
rect 1140 -1330 1160 -1310
rect 1180 -1330 1200 -1310
rect 1220 -1330 1240 -1310
rect 1260 -1330 1280 -1310
rect 1300 -1330 1320 -1310
rect 1340 -1330 1360 -1310
rect 1380 -1330 1400 -1310
rect 1420 -1330 1440 -1310
rect 1460 -1330 1470 -1310
rect 670 -1500 1470 -1330
rect 670 -1520 680 -1500
rect 700 -1520 720 -1500
rect 740 -1520 760 -1500
rect 780 -1520 800 -1500
rect 820 -1520 840 -1500
rect 860 -1520 880 -1500
rect 900 -1520 920 -1500
rect 940 -1520 960 -1500
rect 980 -1520 1000 -1500
rect 1020 -1520 1040 -1500
rect 1060 -1520 1080 -1500
rect 1100 -1520 1120 -1500
rect 1140 -1520 1160 -1500
rect 1180 -1520 1200 -1500
rect 1220 -1520 1240 -1500
rect 1260 -1520 1280 -1500
rect 1300 -1520 1320 -1500
rect 1340 -1520 1360 -1500
rect 1380 -1520 1400 -1500
rect 1420 -1520 1440 -1500
rect 1460 -1520 1470 -1500
rect 670 -1690 1470 -1520
rect 670 -1710 680 -1690
rect 700 -1710 720 -1690
rect 740 -1710 760 -1690
rect 780 -1710 800 -1690
rect 820 -1710 840 -1690
rect 860 -1710 880 -1690
rect 900 -1710 920 -1690
rect 940 -1710 960 -1690
rect 980 -1710 1000 -1690
rect 1020 -1710 1040 -1690
rect 1060 -1710 1080 -1690
rect 1100 -1710 1120 -1690
rect 1140 -1710 1160 -1690
rect 1180 -1710 1200 -1690
rect 1220 -1710 1240 -1690
rect 1260 -1710 1280 -1690
rect 1300 -1710 1320 -1690
rect 1340 -1710 1360 -1690
rect 1380 -1710 1400 -1690
rect 1420 -1710 1440 -1690
rect 1460 -1710 1470 -1690
rect 670 -1880 1470 -1710
rect 670 -1900 680 -1880
rect 700 -1900 720 -1880
rect 740 -1900 760 -1880
rect 780 -1900 800 -1880
rect 820 -1900 840 -1880
rect 860 -1900 880 -1880
rect 900 -1900 920 -1880
rect 940 -1900 960 -1880
rect 980 -1900 1000 -1880
rect 1020 -1900 1040 -1880
rect 1060 -1900 1080 -1880
rect 1100 -1900 1120 -1880
rect 1140 -1900 1160 -1880
rect 1180 -1900 1200 -1880
rect 1220 -1900 1240 -1880
rect 1260 -1900 1280 -1880
rect 1300 -1900 1320 -1880
rect 1340 -1900 1360 -1880
rect 1380 -1900 1400 -1880
rect 1420 -1900 1440 -1880
rect 1460 -1900 1470 -1880
rect 670 -2070 1470 -1900
rect 670 -2090 680 -2070
rect 700 -2090 720 -2070
rect 740 -2090 760 -2070
rect 780 -2090 800 -2070
rect 820 -2090 840 -2070
rect 860 -2090 880 -2070
rect 900 -2090 920 -2070
rect 940 -2090 960 -2070
rect 980 -2090 1000 -2070
rect 1020 -2090 1040 -2070
rect 1060 -2090 1080 -2070
rect 1100 -2090 1120 -2070
rect 1140 -2090 1160 -2070
rect 1180 -2090 1200 -2070
rect 1220 -2090 1240 -2070
rect 1260 -2090 1280 -2070
rect 1300 -2090 1320 -2070
rect 1340 -2090 1360 -2070
rect 1380 -2090 1400 -2070
rect 1420 -2090 1440 -2070
rect 1460 -2090 1470 -2070
rect 670 -2260 1470 -2090
rect 670 -2280 680 -2260
rect 700 -2280 720 -2260
rect 740 -2280 760 -2260
rect 780 -2280 800 -2260
rect 820 -2280 840 -2260
rect 860 -2280 880 -2260
rect 900 -2280 920 -2260
rect 940 -2280 960 -2260
rect 980 -2280 1000 -2260
rect 1020 -2280 1040 -2260
rect 1060 -2280 1080 -2260
rect 1100 -2280 1120 -2260
rect 1140 -2280 1160 -2260
rect 1180 -2280 1200 -2260
rect 1220 -2280 1240 -2260
rect 1260 -2280 1280 -2260
rect 1300 -2280 1320 -2260
rect 1340 -2280 1360 -2260
rect 1380 -2280 1400 -2260
rect 1420 -2280 1440 -2260
rect 1460 -2280 1470 -2260
rect 670 -2450 1470 -2280
rect 670 -2470 680 -2450
rect 700 -2470 720 -2450
rect 740 -2470 760 -2450
rect 780 -2470 800 -2450
rect 820 -2470 840 -2450
rect 860 -2470 880 -2450
rect 900 -2470 920 -2450
rect 940 -2470 960 -2450
rect 980 -2470 1000 -2450
rect 1020 -2470 1040 -2450
rect 1060 -2470 1080 -2450
rect 1100 -2470 1120 -2450
rect 1140 -2470 1160 -2450
rect 1180 -2470 1200 -2450
rect 1220 -2470 1240 -2450
rect 1260 -2470 1280 -2450
rect 1300 -2470 1320 -2450
rect 1340 -2470 1360 -2450
rect 1380 -2470 1400 -2450
rect 1420 -2470 1440 -2450
rect 1460 -2470 1470 -2450
rect 670 -2640 1470 -2470
rect 670 -2660 680 -2640
rect 700 -2660 720 -2640
rect 740 -2660 760 -2640
rect 780 -2660 800 -2640
rect 820 -2660 840 -2640
rect 860 -2660 880 -2640
rect 900 -2660 920 -2640
rect 940 -2660 960 -2640
rect 980 -2660 1000 -2640
rect 1020 -2660 1040 -2640
rect 1060 -2660 1080 -2640
rect 1100 -2660 1120 -2640
rect 1140 -2660 1160 -2640
rect 1180 -2660 1200 -2640
rect 1220 -2660 1240 -2640
rect 1260 -2660 1280 -2640
rect 1300 -2660 1320 -2640
rect 1340 -2660 1360 -2640
rect 1380 -2660 1400 -2640
rect 1420 -2660 1440 -2640
rect 1460 -2660 1470 -2640
rect 670 -2670 1470 -2660
rect 1750 -225 2550 -215
rect 1750 -245 1760 -225
rect 1780 -245 1800 -225
rect 1820 -245 1840 -225
rect 1860 -245 1880 -225
rect 1900 -245 1920 -225
rect 1940 -245 1960 -225
rect 1980 -245 2000 -225
rect 2020 -245 2040 -225
rect 2060 -245 2080 -225
rect 2100 -245 2120 -225
rect 2140 -245 2160 -225
rect 2180 -245 2200 -225
rect 2220 -245 2240 -225
rect 2260 -245 2280 -225
rect 2300 -245 2320 -225
rect 2340 -245 2360 -225
rect 2380 -245 2400 -225
rect 2420 -245 2440 -225
rect 2460 -245 2480 -225
rect 2500 -245 2520 -225
rect 2540 -245 2550 -225
rect 1750 -265 2550 -245
rect 1750 -285 1760 -265
rect 1780 -285 1800 -265
rect 1820 -285 1840 -265
rect 1860 -285 1880 -265
rect 1900 -285 1920 -265
rect 1940 -285 1960 -265
rect 1980 -285 2000 -265
rect 2020 -285 2040 -265
rect 2060 -285 2080 -265
rect 2100 -285 2120 -265
rect 2140 -285 2160 -265
rect 2180 -285 2200 -265
rect 2220 -285 2240 -265
rect 2260 -285 2280 -265
rect 2300 -285 2320 -265
rect 2340 -285 2360 -265
rect 2380 -285 2400 -265
rect 2420 -285 2440 -265
rect 2460 -285 2480 -265
rect 2500 -285 2520 -265
rect 2540 -285 2550 -265
rect 1750 -455 2550 -285
rect 1750 -475 1760 -455
rect 1780 -475 1800 -455
rect 1820 -475 1840 -455
rect 1860 -475 1880 -455
rect 1900 -475 1920 -455
rect 1940 -475 1960 -455
rect 1980 -475 2000 -455
rect 2020 -475 2040 -455
rect 2060 -475 2080 -455
rect 2100 -475 2120 -455
rect 2140 -475 2160 -455
rect 2180 -475 2200 -455
rect 2220 -475 2240 -455
rect 2260 -475 2280 -455
rect 2300 -475 2320 -455
rect 2340 -475 2360 -455
rect 2380 -475 2400 -455
rect 2420 -475 2440 -455
rect 2460 -475 2480 -455
rect 2500 -475 2520 -455
rect 2540 -475 2550 -455
rect 1750 -645 2550 -475
rect 1750 -665 1760 -645
rect 1780 -665 1800 -645
rect 1820 -665 1840 -645
rect 1860 -665 1880 -645
rect 1900 -665 1920 -645
rect 1940 -665 1960 -645
rect 1980 -665 2000 -645
rect 2020 -665 2040 -645
rect 2060 -665 2080 -645
rect 2100 -665 2120 -645
rect 2140 -665 2160 -645
rect 2180 -665 2200 -645
rect 2220 -665 2240 -645
rect 2260 -665 2280 -645
rect 2300 -665 2320 -645
rect 2340 -665 2360 -645
rect 2380 -665 2400 -645
rect 2420 -665 2440 -645
rect 2460 -665 2480 -645
rect 2500 -665 2520 -645
rect 2540 -665 2550 -645
rect 1750 -835 2550 -665
rect 1750 -855 1760 -835
rect 1780 -855 1800 -835
rect 1820 -855 1840 -835
rect 1860 -855 1880 -835
rect 1900 -855 1920 -835
rect 1940 -855 1960 -835
rect 1980 -855 2000 -835
rect 2020 -855 2040 -835
rect 2060 -855 2080 -835
rect 2100 -855 2120 -835
rect 2140 -855 2160 -835
rect 2180 -855 2200 -835
rect 2220 -855 2240 -835
rect 2260 -855 2280 -835
rect 2300 -855 2320 -835
rect 2340 -855 2360 -835
rect 2380 -855 2400 -835
rect 2420 -855 2440 -835
rect 2460 -855 2480 -835
rect 2500 -855 2520 -835
rect 2540 -855 2550 -835
rect 1750 -1025 2550 -855
rect 1750 -1045 1760 -1025
rect 1780 -1045 1800 -1025
rect 1820 -1045 1840 -1025
rect 1860 -1045 1880 -1025
rect 1900 -1045 1920 -1025
rect 1940 -1045 1960 -1025
rect 1980 -1045 2000 -1025
rect 2020 -1045 2040 -1025
rect 2060 -1045 2080 -1025
rect 2100 -1045 2120 -1025
rect 2140 -1045 2160 -1025
rect 2180 -1045 2200 -1025
rect 2220 -1045 2240 -1025
rect 2260 -1045 2280 -1025
rect 2300 -1045 2320 -1025
rect 2340 -1045 2360 -1025
rect 2380 -1045 2400 -1025
rect 2420 -1045 2440 -1025
rect 2460 -1045 2480 -1025
rect 2500 -1045 2520 -1025
rect 2540 -1045 2550 -1025
rect 1750 -1215 2550 -1045
rect 1750 -1235 1760 -1215
rect 1780 -1235 1800 -1215
rect 1820 -1235 1840 -1215
rect 1860 -1235 1880 -1215
rect 1900 -1235 1920 -1215
rect 1940 -1235 1960 -1215
rect 1980 -1235 2000 -1215
rect 2020 -1235 2040 -1215
rect 2060 -1235 2080 -1215
rect 2100 -1235 2120 -1215
rect 2140 -1235 2160 -1215
rect 2180 -1235 2200 -1215
rect 2220 -1235 2240 -1215
rect 2260 -1235 2280 -1215
rect 2300 -1235 2320 -1215
rect 2340 -1235 2360 -1215
rect 2380 -1235 2400 -1215
rect 2420 -1235 2440 -1215
rect 2460 -1235 2480 -1215
rect 2500 -1235 2520 -1215
rect 2540 -1235 2550 -1215
rect 1750 -1405 2550 -1235
rect 1750 -1425 1760 -1405
rect 1780 -1425 1800 -1405
rect 1820 -1425 1840 -1405
rect 1860 -1425 1880 -1405
rect 1900 -1425 1920 -1405
rect 1940 -1425 1960 -1405
rect 1980 -1425 2000 -1405
rect 2020 -1425 2040 -1405
rect 2060 -1425 2080 -1405
rect 2100 -1425 2120 -1405
rect 2140 -1425 2160 -1405
rect 2180 -1425 2200 -1405
rect 2220 -1425 2240 -1405
rect 2260 -1425 2280 -1405
rect 2300 -1425 2320 -1405
rect 2340 -1425 2360 -1405
rect 2380 -1425 2400 -1405
rect 2420 -1425 2440 -1405
rect 2460 -1425 2480 -1405
rect 2500 -1425 2520 -1405
rect 2540 -1425 2550 -1405
rect 1750 -1595 2550 -1425
rect 1750 -1615 1760 -1595
rect 1780 -1615 1800 -1595
rect 1820 -1615 1840 -1595
rect 1860 -1615 1880 -1595
rect 1900 -1615 1920 -1595
rect 1940 -1615 1960 -1595
rect 1980 -1615 2000 -1595
rect 2020 -1615 2040 -1595
rect 2060 -1615 2080 -1595
rect 2100 -1615 2120 -1595
rect 2140 -1615 2160 -1595
rect 2180 -1615 2200 -1595
rect 2220 -1615 2240 -1595
rect 2260 -1615 2280 -1595
rect 2300 -1615 2320 -1595
rect 2340 -1615 2360 -1595
rect 2380 -1615 2400 -1595
rect 2420 -1615 2440 -1595
rect 2460 -1615 2480 -1595
rect 2500 -1615 2520 -1595
rect 2540 -1615 2550 -1595
rect 1750 -1785 2550 -1615
rect 1750 -1805 1760 -1785
rect 1780 -1805 1800 -1785
rect 1820 -1805 1840 -1785
rect 1860 -1805 1880 -1785
rect 1900 -1805 1920 -1785
rect 1940 -1805 1960 -1785
rect 1980 -1805 2000 -1785
rect 2020 -1805 2040 -1785
rect 2060 -1805 2080 -1785
rect 2100 -1805 2120 -1785
rect 2140 -1805 2160 -1785
rect 2180 -1805 2200 -1785
rect 2220 -1805 2240 -1785
rect 2260 -1805 2280 -1785
rect 2300 -1805 2320 -1785
rect 2340 -1805 2360 -1785
rect 2380 -1805 2400 -1785
rect 2420 -1805 2440 -1785
rect 2460 -1805 2480 -1785
rect 2500 -1805 2520 -1785
rect 2540 -1805 2550 -1785
rect 1750 -1975 2550 -1805
rect 1750 -1995 1760 -1975
rect 1780 -1995 1800 -1975
rect 1820 -1995 1840 -1975
rect 1860 -1995 1880 -1975
rect 1900 -1995 1920 -1975
rect 1940 -1995 1960 -1975
rect 1980 -1995 2000 -1975
rect 2020 -1995 2040 -1975
rect 2060 -1995 2080 -1975
rect 2100 -1995 2120 -1975
rect 2140 -1995 2160 -1975
rect 2180 -1995 2200 -1975
rect 2220 -1995 2240 -1975
rect 2260 -1995 2280 -1975
rect 2300 -1995 2320 -1975
rect 2340 -1995 2360 -1975
rect 2380 -1995 2400 -1975
rect 2420 -1995 2440 -1975
rect 2460 -1995 2480 -1975
rect 2500 -1995 2520 -1975
rect 2540 -1995 2550 -1975
rect 1750 -2165 2550 -1995
rect 1750 -2185 1760 -2165
rect 1780 -2185 1800 -2165
rect 1820 -2185 1840 -2165
rect 1860 -2185 1880 -2165
rect 1900 -2185 1920 -2165
rect 1940 -2185 1960 -2165
rect 1980 -2185 2000 -2165
rect 2020 -2185 2040 -2165
rect 2060 -2185 2080 -2165
rect 2100 -2185 2120 -2165
rect 2140 -2185 2160 -2165
rect 2180 -2185 2200 -2165
rect 2220 -2185 2240 -2165
rect 2260 -2185 2280 -2165
rect 2300 -2185 2320 -2165
rect 2340 -2185 2360 -2165
rect 2380 -2185 2400 -2165
rect 2420 -2185 2440 -2165
rect 2460 -2185 2480 -2165
rect 2500 -2185 2520 -2165
rect 2540 -2185 2550 -2165
rect 1750 -2355 2550 -2185
rect 1750 -2375 1760 -2355
rect 1780 -2375 1800 -2355
rect 1820 -2375 1840 -2355
rect 1860 -2375 1880 -2355
rect 1900 -2375 1920 -2355
rect 1940 -2375 1960 -2355
rect 1980 -2375 2000 -2355
rect 2020 -2375 2040 -2355
rect 2060 -2375 2080 -2355
rect 2100 -2375 2120 -2355
rect 2140 -2375 2160 -2355
rect 2180 -2375 2200 -2355
rect 2220 -2375 2240 -2355
rect 2260 -2375 2280 -2355
rect 2300 -2375 2320 -2355
rect 2340 -2375 2360 -2355
rect 2380 -2375 2400 -2355
rect 2420 -2375 2440 -2355
rect 2460 -2375 2480 -2355
rect 2500 -2375 2520 -2355
rect 2540 -2375 2550 -2355
rect 1750 -2545 2550 -2375
rect 1750 -2565 1760 -2545
rect 1780 -2565 1800 -2545
rect 1820 -2565 1840 -2545
rect 1860 -2565 1880 -2545
rect 1900 -2565 1920 -2545
rect 1940 -2565 1960 -2545
rect 1980 -2565 2000 -2545
rect 2020 -2565 2040 -2545
rect 2060 -2565 2080 -2545
rect 2100 -2565 2120 -2545
rect 2140 -2565 2160 -2545
rect 2180 -2565 2200 -2545
rect 2220 -2565 2240 -2545
rect 2260 -2565 2280 -2545
rect 2300 -2565 2320 -2545
rect 2340 -2565 2360 -2545
rect 2380 -2565 2400 -2545
rect 2420 -2565 2440 -2545
rect 2460 -2565 2480 -2545
rect 2500 -2565 2520 -2545
rect 2540 -2565 2550 -2545
rect -70 -2710 -60 -2685
rect -40 -2710 -20 -2685
rect 0 -2710 20 -2685
rect 40 -2710 60 -2685
rect 80 -2710 85 -2685
rect -70 -2720 85 -2710
rect 1750 -2735 2550 -2565
rect 1750 -2755 1760 -2735
rect 1780 -2755 1800 -2735
rect 1820 -2755 1840 -2735
rect 1860 -2755 1880 -2735
rect 1900 -2755 1920 -2735
rect 1940 -2755 1960 -2735
rect 1980 -2755 2000 -2735
rect 2020 -2755 2040 -2735
rect 2060 -2755 2080 -2735
rect 2100 -2755 2120 -2735
rect 2140 -2755 2160 -2735
rect 2180 -2755 2200 -2735
rect 2220 -2755 2240 -2735
rect 2260 -2755 2280 -2735
rect 2300 -2755 2320 -2735
rect 2340 -2755 2360 -2735
rect 2380 -2755 2400 -2735
rect 2420 -2755 2440 -2735
rect 2460 -2755 2480 -2735
rect 2500 -2755 2520 -2735
rect 2540 -2755 2550 -2735
rect 1750 -2775 2550 -2755
rect 1750 -2795 1760 -2775
rect 1780 -2795 1800 -2775
rect 1820 -2795 1840 -2775
rect 1860 -2795 1880 -2775
rect 1900 -2795 1920 -2775
rect 1940 -2795 1960 -2775
rect 1980 -2795 2000 -2775
rect 2020 -2795 2040 -2775
rect 2060 -2795 2080 -2775
rect 2100 -2795 2120 -2775
rect 2140 -2795 2160 -2775
rect 2180 -2795 2200 -2775
rect 2220 -2795 2240 -2775
rect 2260 -2795 2280 -2775
rect 2300 -2795 2320 -2775
rect 2340 -2795 2360 -2775
rect 2380 -2795 2400 -2775
rect 2420 -2795 2440 -2775
rect 2460 -2795 2480 -2775
rect 2500 -2795 2520 -2775
rect 2540 -2795 2550 -2775
rect 1750 -2810 2550 -2795
<< comment >>
rect -75 -85 -70 -80
<< labels >>
rlabel metal1 9 1084 9 1084 1 g_u
port 3 n
rlabel metal1 1070 -95 1070 -95 1 Vout
port 1 n
rlabel metal1 2150 -1110 2150 -1110 1 GND
port 8 n
rlabel metal1 -59 -1509 -59 -1509 1 g_d
port 4 n
rlabel metal1 2235 2380 2235 2380 1 VDD
port 9 n
<< end >>
