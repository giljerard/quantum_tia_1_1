magic
tech sky130A
timestamp 1640986943
<< dnwell >>
rect -5805 6155 -2885 8650
rect -2255 6155 665 8650
<< nwell >>
rect -5845 8545 -2845 8690
rect -5845 6260 -5700 8545
rect -2990 6260 -2845 8545
rect -5845 6115 -2845 6260
rect -2295 8545 705 8690
rect -2295 6260 -2150 8545
rect 560 6260 705 8545
rect -2295 6115 705 6260
<< pwell >>
rect -5700 6260 -2990 8545
rect -2150 6260 560 8545
<< nmos >>
rect -5595 5965 -3095 6010
rect -2045 5965 455 6010
rect -5595 5870 -3095 5915
rect -2045 5870 455 5915
rect -5595 5775 -3095 5820
rect -2045 5775 455 5820
rect -5595 5680 -3095 5725
rect -2045 5680 455 5725
rect -5595 5585 -3095 5630
rect -2045 5585 455 5630
rect -5595 5490 -3095 5535
rect -2045 5490 455 5535
rect -5595 5395 -3095 5440
rect -2045 5395 455 5440
rect -5595 5300 -3095 5345
rect -2045 5300 455 5345
rect -5595 5205 -3095 5250
rect -2045 5205 455 5250
rect -5595 5110 -3095 5155
rect -2045 5110 455 5155
rect -5595 5015 -3095 5060
rect -2045 5015 455 5060
rect -5595 4920 -3095 4965
rect -2045 4920 455 4965
rect -5595 4825 -3095 4870
rect -2045 4825 455 4870
rect -5595 4730 -3095 4775
rect -2045 4730 455 4775
rect -5595 4635 -3095 4680
rect -2045 4635 455 4680
rect -5595 4540 -3095 4585
rect -2045 4540 455 4585
rect -5595 4445 -3095 4490
rect -2045 4445 455 4490
rect -5595 4350 -3095 4395
rect -2045 4350 455 4395
rect -5595 4255 -3095 4300
rect -2045 4255 455 4300
rect -5595 4160 -3095 4205
rect -2045 4160 455 4205
rect -5595 4065 -3095 4110
rect -2045 4065 455 4110
rect -5595 3970 -3095 4015
rect -2045 3970 455 4015
rect -5595 3875 -3095 3920
rect -2045 3875 455 3920
rect -5595 3780 -3095 3825
rect -2045 3780 455 3825
rect -5595 3685 -3095 3730
rect -2045 3685 455 3730
rect -5595 3590 -3095 3635
rect -2045 3590 455 3635
<< nmoslvt >>
rect -5665 8410 -3165 8442
rect -5665 8328 -3165 8360
rect -5665 8246 -3165 8278
rect -5665 8164 -3165 8196
rect -5665 8082 -3165 8114
rect -5665 8000 -3165 8032
rect -5665 7918 -3165 7950
rect -5665 7836 -3165 7868
rect -5665 7754 -3165 7786
rect -5665 7672 -3165 7704
rect -5665 7590 -3165 7622
rect -5665 7508 -3165 7540
rect -5665 7426 -3165 7458
rect -5665 7344 -3165 7376
rect -5665 7262 -3165 7294
rect -5665 7180 -3165 7212
rect -5665 7098 -3165 7130
rect -5665 7016 -3165 7048
rect -5665 6934 -3165 6966
rect -5665 6852 -3165 6884
rect -5665 6770 -3165 6802
rect -5665 6688 -3165 6720
rect -5665 6606 -3165 6638
rect -5665 6524 -3165 6556
rect -5665 6442 -3165 6474
rect -5665 6360 -3165 6392
rect -1975 8410 525 8442
rect -1975 8328 525 8360
rect -1975 8246 525 8278
rect -1975 8164 525 8196
rect -1975 8082 525 8114
rect -1975 8000 525 8032
rect -1975 7918 525 7950
rect -1975 7836 525 7868
rect -1975 7754 525 7786
rect -1975 7672 525 7704
rect -1975 7590 525 7622
rect -1975 7508 525 7540
rect -1975 7426 525 7458
rect -1975 7344 525 7376
rect -1975 7262 525 7294
rect -1975 7180 525 7212
rect -1975 7098 525 7130
rect -1975 7016 525 7048
rect -1975 6934 525 6966
rect -1975 6852 525 6884
rect -1975 6770 525 6802
rect -1975 6688 525 6720
rect -1975 6606 525 6638
rect -1975 6524 525 6556
rect -1975 6442 525 6474
rect -1975 6360 525 6392
<< ndiff >>
rect -5665 8477 -3165 8490
rect -5665 8457 -5650 8477
rect -5630 8457 -5610 8477
rect -5590 8457 -5570 8477
rect -5550 8457 -5530 8477
rect -5510 8457 -5490 8477
rect -5470 8457 -5450 8477
rect -5430 8457 -5410 8477
rect -5390 8457 -5370 8477
rect -5350 8457 -5330 8477
rect -5310 8457 -5290 8477
rect -5270 8457 -5250 8477
rect -5230 8457 -5210 8477
rect -5190 8457 -5170 8477
rect -5150 8457 -5130 8477
rect -5110 8457 -5090 8477
rect -5070 8457 -5050 8477
rect -5030 8457 -5010 8477
rect -4990 8457 -4970 8477
rect -4950 8457 -4930 8477
rect -4910 8457 -4890 8477
rect -4870 8457 -4850 8477
rect -4830 8457 -4810 8477
rect -4790 8457 -4770 8477
rect -4750 8457 -4730 8477
rect -4710 8457 -4690 8477
rect -4670 8457 -4650 8477
rect -4630 8457 -4610 8477
rect -4590 8457 -4570 8477
rect -4550 8457 -4530 8477
rect -4510 8457 -4490 8477
rect -4470 8457 -4450 8477
rect -4430 8457 -4410 8477
rect -4390 8457 -4370 8477
rect -4350 8457 -4330 8477
rect -4310 8457 -4290 8477
rect -4270 8457 -4250 8477
rect -4230 8457 -4210 8477
rect -4190 8457 -4170 8477
rect -4150 8457 -4130 8477
rect -4110 8457 -4090 8477
rect -4070 8457 -4050 8477
rect -4030 8457 -4010 8477
rect -3990 8457 -3970 8477
rect -3950 8457 -3930 8477
rect -3910 8457 -3890 8477
rect -3870 8457 -3850 8477
rect -3830 8457 -3810 8477
rect -3790 8457 -3770 8477
rect -3750 8457 -3730 8477
rect -3710 8457 -3690 8477
rect -3670 8457 -3650 8477
rect -3630 8457 -3610 8477
rect -3590 8457 -3570 8477
rect -3550 8457 -3530 8477
rect -3510 8457 -3490 8477
rect -3470 8457 -3450 8477
rect -3430 8457 -3410 8477
rect -3390 8457 -3370 8477
rect -3350 8457 -3330 8477
rect -3310 8457 -3290 8477
rect -3270 8457 -3250 8477
rect -3230 8457 -3210 8477
rect -3190 8457 -3165 8477
rect -5665 8442 -3165 8457
rect -5665 8395 -3165 8410
rect -5665 8375 -5650 8395
rect -5630 8375 -5610 8395
rect -5590 8375 -5570 8395
rect -5550 8375 -5530 8395
rect -5510 8375 -5490 8395
rect -5470 8375 -5450 8395
rect -5430 8375 -5410 8395
rect -5390 8375 -5370 8395
rect -5350 8375 -5330 8395
rect -5310 8375 -5290 8395
rect -5270 8375 -5250 8395
rect -5230 8375 -5210 8395
rect -5190 8375 -5170 8395
rect -5150 8375 -5130 8395
rect -5110 8375 -5090 8395
rect -5070 8375 -5050 8395
rect -5030 8375 -5010 8395
rect -4990 8375 -4970 8395
rect -4950 8375 -4930 8395
rect -4910 8375 -4890 8395
rect -4870 8375 -4850 8395
rect -4830 8375 -4810 8395
rect -4790 8375 -4770 8395
rect -4750 8375 -4730 8395
rect -4710 8375 -4690 8395
rect -4670 8375 -4650 8395
rect -4630 8375 -4610 8395
rect -4590 8375 -4570 8395
rect -4550 8375 -4530 8395
rect -4510 8375 -4490 8395
rect -4470 8375 -4450 8395
rect -4430 8375 -4410 8395
rect -4390 8375 -4370 8395
rect -4350 8375 -4330 8395
rect -4310 8375 -4290 8395
rect -4270 8375 -4250 8395
rect -4230 8375 -4210 8395
rect -4190 8375 -4170 8395
rect -4150 8375 -4130 8395
rect -4110 8375 -4090 8395
rect -4070 8375 -4050 8395
rect -4030 8375 -4010 8395
rect -3990 8375 -3970 8395
rect -3950 8375 -3930 8395
rect -3910 8375 -3890 8395
rect -3870 8375 -3850 8395
rect -3830 8375 -3810 8395
rect -3790 8375 -3770 8395
rect -3750 8375 -3730 8395
rect -3710 8375 -3690 8395
rect -3670 8375 -3650 8395
rect -3630 8375 -3610 8395
rect -3590 8375 -3570 8395
rect -3550 8375 -3530 8395
rect -3510 8375 -3490 8395
rect -3470 8375 -3450 8395
rect -3430 8375 -3410 8395
rect -3390 8375 -3370 8395
rect -3350 8375 -3330 8395
rect -3310 8375 -3290 8395
rect -3270 8375 -3250 8395
rect -3230 8375 -3210 8395
rect -3190 8375 -3165 8395
rect -5665 8360 -3165 8375
rect -5665 8313 -3165 8328
rect -5665 8293 -5650 8313
rect -5630 8293 -5610 8313
rect -5590 8293 -5570 8313
rect -5550 8293 -5530 8313
rect -5510 8293 -5490 8313
rect -5470 8293 -5450 8313
rect -5430 8293 -5410 8313
rect -5390 8293 -5370 8313
rect -5350 8293 -5330 8313
rect -5310 8293 -5290 8313
rect -5270 8293 -5250 8313
rect -5230 8293 -5210 8313
rect -5190 8293 -5170 8313
rect -5150 8293 -5130 8313
rect -5110 8293 -5090 8313
rect -5070 8293 -5050 8313
rect -5030 8293 -5010 8313
rect -4990 8293 -4970 8313
rect -4950 8293 -4930 8313
rect -4910 8293 -4890 8313
rect -4870 8293 -4850 8313
rect -4830 8293 -4810 8313
rect -4790 8293 -4770 8313
rect -4750 8293 -4730 8313
rect -4710 8293 -4690 8313
rect -4670 8293 -4650 8313
rect -4630 8293 -4610 8313
rect -4590 8293 -4570 8313
rect -4550 8293 -4530 8313
rect -4510 8293 -4490 8313
rect -4470 8293 -4450 8313
rect -4430 8293 -4410 8313
rect -4390 8293 -4370 8313
rect -4350 8293 -4330 8313
rect -4310 8293 -4290 8313
rect -4270 8293 -4250 8313
rect -4230 8293 -4210 8313
rect -4190 8293 -4170 8313
rect -4150 8293 -4130 8313
rect -4110 8293 -4090 8313
rect -4070 8293 -4050 8313
rect -4030 8293 -4010 8313
rect -3990 8293 -3970 8313
rect -3950 8293 -3930 8313
rect -3910 8293 -3890 8313
rect -3870 8293 -3850 8313
rect -3830 8293 -3810 8313
rect -3790 8293 -3770 8313
rect -3750 8293 -3730 8313
rect -3710 8293 -3690 8313
rect -3670 8293 -3650 8313
rect -3630 8293 -3610 8313
rect -3590 8293 -3570 8313
rect -3550 8293 -3530 8313
rect -3510 8293 -3490 8313
rect -3470 8293 -3450 8313
rect -3430 8293 -3410 8313
rect -3390 8293 -3370 8313
rect -3350 8293 -3330 8313
rect -3310 8293 -3290 8313
rect -3270 8293 -3250 8313
rect -3230 8293 -3210 8313
rect -3190 8293 -3165 8313
rect -5665 8278 -3165 8293
rect -5665 8231 -3165 8246
rect -5665 8211 -5650 8231
rect -5630 8211 -5610 8231
rect -5590 8211 -5570 8231
rect -5550 8211 -5530 8231
rect -5510 8211 -5490 8231
rect -5470 8211 -5450 8231
rect -5430 8211 -5410 8231
rect -5390 8211 -5370 8231
rect -5350 8211 -5330 8231
rect -5310 8211 -5290 8231
rect -5270 8211 -5250 8231
rect -5230 8211 -5210 8231
rect -5190 8211 -5170 8231
rect -5150 8211 -5130 8231
rect -5110 8211 -5090 8231
rect -5070 8211 -5050 8231
rect -5030 8211 -5010 8231
rect -4990 8211 -4970 8231
rect -4950 8211 -4930 8231
rect -4910 8211 -4890 8231
rect -4870 8211 -4850 8231
rect -4830 8211 -4810 8231
rect -4790 8211 -4770 8231
rect -4750 8211 -4730 8231
rect -4710 8211 -4690 8231
rect -4670 8211 -4650 8231
rect -4630 8211 -4610 8231
rect -4590 8211 -4570 8231
rect -4550 8211 -4530 8231
rect -4510 8211 -4490 8231
rect -4470 8211 -4450 8231
rect -4430 8211 -4410 8231
rect -4390 8211 -4370 8231
rect -4350 8211 -4330 8231
rect -4310 8211 -4290 8231
rect -4270 8211 -4250 8231
rect -4230 8211 -4210 8231
rect -4190 8211 -4170 8231
rect -4150 8211 -4130 8231
rect -4110 8211 -4090 8231
rect -4070 8211 -4050 8231
rect -4030 8211 -4010 8231
rect -3990 8211 -3970 8231
rect -3950 8211 -3930 8231
rect -3910 8211 -3890 8231
rect -3870 8211 -3850 8231
rect -3830 8211 -3810 8231
rect -3790 8211 -3770 8231
rect -3750 8211 -3730 8231
rect -3710 8211 -3690 8231
rect -3670 8211 -3650 8231
rect -3630 8211 -3610 8231
rect -3590 8211 -3570 8231
rect -3550 8211 -3530 8231
rect -3510 8211 -3490 8231
rect -3470 8211 -3450 8231
rect -3430 8211 -3410 8231
rect -3390 8211 -3370 8231
rect -3350 8211 -3330 8231
rect -3310 8211 -3290 8231
rect -3270 8211 -3250 8231
rect -3230 8211 -3210 8231
rect -3190 8211 -3165 8231
rect -5665 8196 -3165 8211
rect -5665 8149 -3165 8164
rect -5665 8129 -5650 8149
rect -5630 8129 -5610 8149
rect -5590 8129 -5570 8149
rect -5550 8129 -5530 8149
rect -5510 8129 -5490 8149
rect -5470 8129 -5450 8149
rect -5430 8129 -5410 8149
rect -5390 8129 -5370 8149
rect -5350 8129 -5330 8149
rect -5310 8129 -5290 8149
rect -5270 8129 -5250 8149
rect -5230 8129 -5210 8149
rect -5190 8129 -5170 8149
rect -5150 8129 -5130 8149
rect -5110 8129 -5090 8149
rect -5070 8129 -5050 8149
rect -5030 8129 -5010 8149
rect -4990 8129 -4970 8149
rect -4950 8129 -4930 8149
rect -4910 8129 -4890 8149
rect -4870 8129 -4850 8149
rect -4830 8129 -4810 8149
rect -4790 8129 -4770 8149
rect -4750 8129 -4730 8149
rect -4710 8129 -4690 8149
rect -4670 8129 -4650 8149
rect -4630 8129 -4610 8149
rect -4590 8129 -4570 8149
rect -4550 8129 -4530 8149
rect -4510 8129 -4490 8149
rect -4470 8129 -4450 8149
rect -4430 8129 -4410 8149
rect -4390 8129 -4370 8149
rect -4350 8129 -4330 8149
rect -4310 8129 -4290 8149
rect -4270 8129 -4250 8149
rect -4230 8129 -4210 8149
rect -4190 8129 -4170 8149
rect -4150 8129 -4130 8149
rect -4110 8129 -4090 8149
rect -4070 8129 -4050 8149
rect -4030 8129 -4010 8149
rect -3990 8129 -3970 8149
rect -3950 8129 -3930 8149
rect -3910 8129 -3890 8149
rect -3870 8129 -3850 8149
rect -3830 8129 -3810 8149
rect -3790 8129 -3770 8149
rect -3750 8129 -3730 8149
rect -3710 8129 -3690 8149
rect -3670 8129 -3650 8149
rect -3630 8129 -3610 8149
rect -3590 8129 -3570 8149
rect -3550 8129 -3530 8149
rect -3510 8129 -3490 8149
rect -3470 8129 -3450 8149
rect -3430 8129 -3410 8149
rect -3390 8129 -3370 8149
rect -3350 8129 -3330 8149
rect -3310 8129 -3290 8149
rect -3270 8129 -3250 8149
rect -3230 8129 -3210 8149
rect -3190 8129 -3165 8149
rect -5665 8114 -3165 8129
rect -5665 8067 -3165 8082
rect -5665 8047 -5650 8067
rect -5630 8047 -5610 8067
rect -5590 8047 -5570 8067
rect -5550 8047 -5530 8067
rect -5510 8047 -5490 8067
rect -5470 8047 -5450 8067
rect -5430 8047 -5410 8067
rect -5390 8047 -5370 8067
rect -5350 8047 -5330 8067
rect -5310 8047 -5290 8067
rect -5270 8047 -5250 8067
rect -5230 8047 -5210 8067
rect -5190 8047 -5170 8067
rect -5150 8047 -5130 8067
rect -5110 8047 -5090 8067
rect -5070 8047 -5050 8067
rect -5030 8047 -5010 8067
rect -4990 8047 -4970 8067
rect -4950 8047 -4930 8067
rect -4910 8047 -4890 8067
rect -4870 8047 -4850 8067
rect -4830 8047 -4810 8067
rect -4790 8047 -4770 8067
rect -4750 8047 -4730 8067
rect -4710 8047 -4690 8067
rect -4670 8047 -4650 8067
rect -4630 8047 -4610 8067
rect -4590 8047 -4570 8067
rect -4550 8047 -4530 8067
rect -4510 8047 -4490 8067
rect -4470 8047 -4450 8067
rect -4430 8047 -4410 8067
rect -4390 8047 -4370 8067
rect -4350 8047 -4330 8067
rect -4310 8047 -4290 8067
rect -4270 8047 -4250 8067
rect -4230 8047 -4210 8067
rect -4190 8047 -4170 8067
rect -4150 8047 -4130 8067
rect -4110 8047 -4090 8067
rect -4070 8047 -4050 8067
rect -4030 8047 -4010 8067
rect -3990 8047 -3970 8067
rect -3950 8047 -3930 8067
rect -3910 8047 -3890 8067
rect -3870 8047 -3850 8067
rect -3830 8047 -3810 8067
rect -3790 8047 -3770 8067
rect -3750 8047 -3730 8067
rect -3710 8047 -3690 8067
rect -3670 8047 -3650 8067
rect -3630 8047 -3610 8067
rect -3590 8047 -3570 8067
rect -3550 8047 -3530 8067
rect -3510 8047 -3490 8067
rect -3470 8047 -3450 8067
rect -3430 8047 -3410 8067
rect -3390 8047 -3370 8067
rect -3350 8047 -3330 8067
rect -3310 8047 -3290 8067
rect -3270 8047 -3250 8067
rect -3230 8047 -3210 8067
rect -3190 8047 -3165 8067
rect -5665 8032 -3165 8047
rect -5665 7985 -3165 8000
rect -5665 7965 -5650 7985
rect -5630 7965 -5610 7985
rect -5590 7965 -5570 7985
rect -5550 7965 -5530 7985
rect -5510 7965 -5490 7985
rect -5470 7965 -5450 7985
rect -5430 7965 -5410 7985
rect -5390 7965 -5370 7985
rect -5350 7965 -5330 7985
rect -5310 7965 -5290 7985
rect -5270 7965 -5250 7985
rect -5230 7965 -5210 7985
rect -5190 7965 -5170 7985
rect -5150 7965 -5130 7985
rect -5110 7965 -5090 7985
rect -5070 7965 -5050 7985
rect -5030 7965 -5010 7985
rect -4990 7965 -4970 7985
rect -4950 7965 -4930 7985
rect -4910 7965 -4890 7985
rect -4870 7965 -4850 7985
rect -4830 7965 -4810 7985
rect -4790 7965 -4770 7985
rect -4750 7965 -4730 7985
rect -4710 7965 -4690 7985
rect -4670 7965 -4650 7985
rect -4630 7965 -4610 7985
rect -4590 7965 -4570 7985
rect -4550 7965 -4530 7985
rect -4510 7965 -4490 7985
rect -4470 7965 -4450 7985
rect -4430 7965 -4410 7985
rect -4390 7965 -4370 7985
rect -4350 7965 -4330 7985
rect -4310 7965 -4290 7985
rect -4270 7965 -4250 7985
rect -4230 7965 -4210 7985
rect -4190 7965 -4170 7985
rect -4150 7965 -4130 7985
rect -4110 7965 -4090 7985
rect -4070 7965 -4050 7985
rect -4030 7965 -4010 7985
rect -3990 7965 -3970 7985
rect -3950 7965 -3930 7985
rect -3910 7965 -3890 7985
rect -3870 7965 -3850 7985
rect -3830 7965 -3810 7985
rect -3790 7965 -3770 7985
rect -3750 7965 -3730 7985
rect -3710 7965 -3690 7985
rect -3670 7965 -3650 7985
rect -3630 7965 -3610 7985
rect -3590 7965 -3570 7985
rect -3550 7965 -3530 7985
rect -3510 7965 -3490 7985
rect -3470 7965 -3450 7985
rect -3430 7965 -3410 7985
rect -3390 7965 -3370 7985
rect -3350 7965 -3330 7985
rect -3310 7965 -3290 7985
rect -3270 7965 -3250 7985
rect -3230 7965 -3210 7985
rect -3190 7965 -3165 7985
rect -5665 7950 -3165 7965
rect -5665 7903 -3165 7918
rect -5665 7883 -5650 7903
rect -5630 7883 -5610 7903
rect -5590 7883 -5570 7903
rect -5550 7883 -5530 7903
rect -5510 7883 -5490 7903
rect -5470 7883 -5450 7903
rect -5430 7883 -5410 7903
rect -5390 7883 -5370 7903
rect -5350 7883 -5330 7903
rect -5310 7883 -5290 7903
rect -5270 7883 -5250 7903
rect -5230 7883 -5210 7903
rect -5190 7883 -5170 7903
rect -5150 7883 -5130 7903
rect -5110 7883 -5090 7903
rect -5070 7883 -5050 7903
rect -5030 7883 -5010 7903
rect -4990 7883 -4970 7903
rect -4950 7883 -4930 7903
rect -4910 7883 -4890 7903
rect -4870 7883 -4850 7903
rect -4830 7883 -4810 7903
rect -4790 7883 -4770 7903
rect -4750 7883 -4730 7903
rect -4710 7883 -4690 7903
rect -4670 7883 -4650 7903
rect -4630 7883 -4610 7903
rect -4590 7883 -4570 7903
rect -4550 7883 -4530 7903
rect -4510 7883 -4490 7903
rect -4470 7883 -4450 7903
rect -4430 7883 -4410 7903
rect -4390 7883 -4370 7903
rect -4350 7883 -4330 7903
rect -4310 7883 -4290 7903
rect -4270 7883 -4250 7903
rect -4230 7883 -4210 7903
rect -4190 7883 -4170 7903
rect -4150 7883 -4130 7903
rect -4110 7883 -4090 7903
rect -4070 7883 -4050 7903
rect -4030 7883 -4010 7903
rect -3990 7883 -3970 7903
rect -3950 7883 -3930 7903
rect -3910 7883 -3890 7903
rect -3870 7883 -3850 7903
rect -3830 7883 -3810 7903
rect -3790 7883 -3770 7903
rect -3750 7883 -3730 7903
rect -3710 7883 -3690 7903
rect -3670 7883 -3650 7903
rect -3630 7883 -3610 7903
rect -3590 7883 -3570 7903
rect -3550 7883 -3530 7903
rect -3510 7883 -3490 7903
rect -3470 7883 -3450 7903
rect -3430 7883 -3410 7903
rect -3390 7883 -3370 7903
rect -3350 7883 -3330 7903
rect -3310 7883 -3290 7903
rect -3270 7883 -3250 7903
rect -3230 7883 -3210 7903
rect -3190 7883 -3165 7903
rect -5665 7868 -3165 7883
rect -5665 7821 -3165 7836
rect -5665 7801 -5650 7821
rect -5630 7801 -5610 7821
rect -5590 7801 -5570 7821
rect -5550 7801 -5530 7821
rect -5510 7801 -5490 7821
rect -5470 7801 -5450 7821
rect -5430 7801 -5410 7821
rect -5390 7801 -5370 7821
rect -5350 7801 -5330 7821
rect -5310 7801 -5290 7821
rect -5270 7801 -5250 7821
rect -5230 7801 -5210 7821
rect -5190 7801 -5170 7821
rect -5150 7801 -5130 7821
rect -5110 7801 -5090 7821
rect -5070 7801 -5050 7821
rect -5030 7801 -5010 7821
rect -4990 7801 -4970 7821
rect -4950 7801 -4930 7821
rect -4910 7801 -4890 7821
rect -4870 7801 -4850 7821
rect -4830 7801 -4810 7821
rect -4790 7801 -4770 7821
rect -4750 7801 -4730 7821
rect -4710 7801 -4690 7821
rect -4670 7801 -4650 7821
rect -4630 7801 -4610 7821
rect -4590 7801 -4570 7821
rect -4550 7801 -4530 7821
rect -4510 7801 -4490 7821
rect -4470 7801 -4450 7821
rect -4430 7801 -4410 7821
rect -4390 7801 -4370 7821
rect -4350 7801 -4330 7821
rect -4310 7801 -4290 7821
rect -4270 7801 -4250 7821
rect -4230 7801 -4210 7821
rect -4190 7801 -4170 7821
rect -4150 7801 -4130 7821
rect -4110 7801 -4090 7821
rect -4070 7801 -4050 7821
rect -4030 7801 -4010 7821
rect -3990 7801 -3970 7821
rect -3950 7801 -3930 7821
rect -3910 7801 -3890 7821
rect -3870 7801 -3850 7821
rect -3830 7801 -3810 7821
rect -3790 7801 -3770 7821
rect -3750 7801 -3730 7821
rect -3710 7801 -3690 7821
rect -3670 7801 -3650 7821
rect -3630 7801 -3610 7821
rect -3590 7801 -3570 7821
rect -3550 7801 -3530 7821
rect -3510 7801 -3490 7821
rect -3470 7801 -3450 7821
rect -3430 7801 -3410 7821
rect -3390 7801 -3370 7821
rect -3350 7801 -3330 7821
rect -3310 7801 -3290 7821
rect -3270 7801 -3250 7821
rect -3230 7801 -3210 7821
rect -3190 7801 -3165 7821
rect -5665 7786 -3165 7801
rect -5665 7739 -3165 7754
rect -5665 7719 -5650 7739
rect -5630 7719 -5610 7739
rect -5590 7719 -5570 7739
rect -5550 7719 -5530 7739
rect -5510 7719 -5490 7739
rect -5470 7719 -5450 7739
rect -5430 7719 -5410 7739
rect -5390 7719 -5370 7739
rect -5350 7719 -5330 7739
rect -5310 7719 -5290 7739
rect -5270 7719 -5250 7739
rect -5230 7719 -5210 7739
rect -5190 7719 -5170 7739
rect -5150 7719 -5130 7739
rect -5110 7719 -5090 7739
rect -5070 7719 -5050 7739
rect -5030 7719 -5010 7739
rect -4990 7719 -4970 7739
rect -4950 7719 -4930 7739
rect -4910 7719 -4890 7739
rect -4870 7719 -4850 7739
rect -4830 7719 -4810 7739
rect -4790 7719 -4770 7739
rect -4750 7719 -4730 7739
rect -4710 7719 -4690 7739
rect -4670 7719 -4650 7739
rect -4630 7719 -4610 7739
rect -4590 7719 -4570 7739
rect -4550 7719 -4530 7739
rect -4510 7719 -4490 7739
rect -4470 7719 -4450 7739
rect -4430 7719 -4410 7739
rect -4390 7719 -4370 7739
rect -4350 7719 -4330 7739
rect -4310 7719 -4290 7739
rect -4270 7719 -4250 7739
rect -4230 7719 -4210 7739
rect -4190 7719 -4170 7739
rect -4150 7719 -4130 7739
rect -4110 7719 -4090 7739
rect -4070 7719 -4050 7739
rect -4030 7719 -4010 7739
rect -3990 7719 -3970 7739
rect -3950 7719 -3930 7739
rect -3910 7719 -3890 7739
rect -3870 7719 -3850 7739
rect -3830 7719 -3810 7739
rect -3790 7719 -3770 7739
rect -3750 7719 -3730 7739
rect -3710 7719 -3690 7739
rect -3670 7719 -3650 7739
rect -3630 7719 -3610 7739
rect -3590 7719 -3570 7739
rect -3550 7719 -3530 7739
rect -3510 7719 -3490 7739
rect -3470 7719 -3450 7739
rect -3430 7719 -3410 7739
rect -3390 7719 -3370 7739
rect -3350 7719 -3330 7739
rect -3310 7719 -3290 7739
rect -3270 7719 -3250 7739
rect -3230 7719 -3210 7739
rect -3190 7719 -3165 7739
rect -5665 7704 -3165 7719
rect -5665 7657 -3165 7672
rect -5665 7637 -5650 7657
rect -5630 7637 -5610 7657
rect -5590 7637 -5570 7657
rect -5550 7637 -5530 7657
rect -5510 7637 -5490 7657
rect -5470 7637 -5450 7657
rect -5430 7637 -5410 7657
rect -5390 7637 -5370 7657
rect -5350 7637 -5330 7657
rect -5310 7637 -5290 7657
rect -5270 7637 -5250 7657
rect -5230 7637 -5210 7657
rect -5190 7637 -5170 7657
rect -5150 7637 -5130 7657
rect -5110 7637 -5090 7657
rect -5070 7637 -5050 7657
rect -5030 7637 -5010 7657
rect -4990 7637 -4970 7657
rect -4950 7637 -4930 7657
rect -4910 7637 -4890 7657
rect -4870 7637 -4850 7657
rect -4830 7637 -4810 7657
rect -4790 7637 -4770 7657
rect -4750 7637 -4730 7657
rect -4710 7637 -4690 7657
rect -4670 7637 -4650 7657
rect -4630 7637 -4610 7657
rect -4590 7637 -4570 7657
rect -4550 7637 -4530 7657
rect -4510 7637 -4490 7657
rect -4470 7637 -4450 7657
rect -4430 7637 -4410 7657
rect -4390 7637 -4370 7657
rect -4350 7637 -4330 7657
rect -4310 7637 -4290 7657
rect -4270 7637 -4250 7657
rect -4230 7637 -4210 7657
rect -4190 7637 -4170 7657
rect -4150 7637 -4130 7657
rect -4110 7637 -4090 7657
rect -4070 7637 -4050 7657
rect -4030 7637 -4010 7657
rect -3990 7637 -3970 7657
rect -3950 7637 -3930 7657
rect -3910 7637 -3890 7657
rect -3870 7637 -3850 7657
rect -3830 7637 -3810 7657
rect -3790 7637 -3770 7657
rect -3750 7637 -3730 7657
rect -3710 7637 -3690 7657
rect -3670 7637 -3650 7657
rect -3630 7637 -3610 7657
rect -3590 7637 -3570 7657
rect -3550 7637 -3530 7657
rect -3510 7637 -3490 7657
rect -3470 7637 -3450 7657
rect -3430 7637 -3410 7657
rect -3390 7637 -3370 7657
rect -3350 7637 -3330 7657
rect -3310 7637 -3290 7657
rect -3270 7637 -3250 7657
rect -3230 7637 -3210 7657
rect -3190 7637 -3165 7657
rect -5665 7622 -3165 7637
rect -5665 7575 -3165 7590
rect -5665 7555 -5650 7575
rect -5630 7555 -5610 7575
rect -5590 7555 -5570 7575
rect -5550 7555 -5530 7575
rect -5510 7555 -5490 7575
rect -5470 7555 -5450 7575
rect -5430 7555 -5410 7575
rect -5390 7555 -5370 7575
rect -5350 7555 -5330 7575
rect -5310 7555 -5290 7575
rect -5270 7555 -5250 7575
rect -5230 7555 -5210 7575
rect -5190 7555 -5170 7575
rect -5150 7555 -5130 7575
rect -5110 7555 -5090 7575
rect -5070 7555 -5050 7575
rect -5030 7555 -5010 7575
rect -4990 7555 -4970 7575
rect -4950 7555 -4930 7575
rect -4910 7555 -4890 7575
rect -4870 7555 -4850 7575
rect -4830 7555 -4810 7575
rect -4790 7555 -4770 7575
rect -4750 7555 -4730 7575
rect -4710 7555 -4690 7575
rect -4670 7555 -4650 7575
rect -4630 7555 -4610 7575
rect -4590 7555 -4570 7575
rect -4550 7555 -4530 7575
rect -4510 7555 -4490 7575
rect -4470 7555 -4450 7575
rect -4430 7555 -4410 7575
rect -4390 7555 -4370 7575
rect -4350 7555 -4330 7575
rect -4310 7555 -4290 7575
rect -4270 7555 -4250 7575
rect -4230 7555 -4210 7575
rect -4190 7555 -4170 7575
rect -4150 7555 -4130 7575
rect -4110 7555 -4090 7575
rect -4070 7555 -4050 7575
rect -4030 7555 -4010 7575
rect -3990 7555 -3970 7575
rect -3950 7555 -3930 7575
rect -3910 7555 -3890 7575
rect -3870 7555 -3850 7575
rect -3830 7555 -3810 7575
rect -3790 7555 -3770 7575
rect -3750 7555 -3730 7575
rect -3710 7555 -3690 7575
rect -3670 7555 -3650 7575
rect -3630 7555 -3610 7575
rect -3590 7555 -3570 7575
rect -3550 7555 -3530 7575
rect -3510 7555 -3490 7575
rect -3470 7555 -3450 7575
rect -3430 7555 -3410 7575
rect -3390 7555 -3370 7575
rect -3350 7555 -3330 7575
rect -3310 7555 -3290 7575
rect -3270 7555 -3250 7575
rect -3230 7555 -3210 7575
rect -3190 7555 -3165 7575
rect -5665 7540 -3165 7555
rect -5665 7493 -3165 7508
rect -5665 7473 -5650 7493
rect -5630 7473 -5610 7493
rect -5590 7473 -5570 7493
rect -5550 7473 -5530 7493
rect -5510 7473 -5490 7493
rect -5470 7473 -5450 7493
rect -5430 7473 -5410 7493
rect -5390 7473 -5370 7493
rect -5350 7473 -5330 7493
rect -5310 7473 -5290 7493
rect -5270 7473 -5250 7493
rect -5230 7473 -5210 7493
rect -5190 7473 -5170 7493
rect -5150 7473 -5130 7493
rect -5110 7473 -5090 7493
rect -5070 7473 -5050 7493
rect -5030 7473 -5010 7493
rect -4990 7473 -4970 7493
rect -4950 7473 -4930 7493
rect -4910 7473 -4890 7493
rect -4870 7473 -4850 7493
rect -4830 7473 -4810 7493
rect -4790 7473 -4770 7493
rect -4750 7473 -4730 7493
rect -4710 7473 -4690 7493
rect -4670 7473 -4650 7493
rect -4630 7473 -4610 7493
rect -4590 7473 -4570 7493
rect -4550 7473 -4530 7493
rect -4510 7473 -4490 7493
rect -4470 7473 -4450 7493
rect -4430 7473 -4410 7493
rect -4390 7473 -4370 7493
rect -4350 7473 -4330 7493
rect -4310 7473 -4290 7493
rect -4270 7473 -4250 7493
rect -4230 7473 -4210 7493
rect -4190 7473 -4170 7493
rect -4150 7473 -4130 7493
rect -4110 7473 -4090 7493
rect -4070 7473 -4050 7493
rect -4030 7473 -4010 7493
rect -3990 7473 -3970 7493
rect -3950 7473 -3930 7493
rect -3910 7473 -3890 7493
rect -3870 7473 -3850 7493
rect -3830 7473 -3810 7493
rect -3790 7473 -3770 7493
rect -3750 7473 -3730 7493
rect -3710 7473 -3690 7493
rect -3670 7473 -3650 7493
rect -3630 7473 -3610 7493
rect -3590 7473 -3570 7493
rect -3550 7473 -3530 7493
rect -3510 7473 -3490 7493
rect -3470 7473 -3450 7493
rect -3430 7473 -3410 7493
rect -3390 7473 -3370 7493
rect -3350 7473 -3330 7493
rect -3310 7473 -3290 7493
rect -3270 7473 -3250 7493
rect -3230 7473 -3210 7493
rect -3190 7473 -3165 7493
rect -5665 7458 -3165 7473
rect -5665 7411 -3165 7426
rect -5665 7391 -5650 7411
rect -5630 7391 -5610 7411
rect -5590 7391 -5570 7411
rect -5550 7391 -5530 7411
rect -5510 7391 -5490 7411
rect -5470 7391 -5450 7411
rect -5430 7391 -5410 7411
rect -5390 7391 -5370 7411
rect -5350 7391 -5330 7411
rect -5310 7391 -5290 7411
rect -5270 7391 -5250 7411
rect -5230 7391 -5210 7411
rect -5190 7391 -5170 7411
rect -5150 7391 -5130 7411
rect -5110 7391 -5090 7411
rect -5070 7391 -5050 7411
rect -5030 7391 -5010 7411
rect -4990 7391 -4970 7411
rect -4950 7391 -4930 7411
rect -4910 7391 -4890 7411
rect -4870 7391 -4850 7411
rect -4830 7391 -4810 7411
rect -4790 7391 -4770 7411
rect -4750 7391 -4730 7411
rect -4710 7391 -4690 7411
rect -4670 7391 -4650 7411
rect -4630 7391 -4610 7411
rect -4590 7391 -4570 7411
rect -4550 7391 -4530 7411
rect -4510 7391 -4490 7411
rect -4470 7391 -4450 7411
rect -4430 7391 -4410 7411
rect -4390 7391 -4370 7411
rect -4350 7391 -4330 7411
rect -4310 7391 -4290 7411
rect -4270 7391 -4250 7411
rect -4230 7391 -4210 7411
rect -4190 7391 -4170 7411
rect -4150 7391 -4130 7411
rect -4110 7391 -4090 7411
rect -4070 7391 -4050 7411
rect -4030 7391 -4010 7411
rect -3990 7391 -3970 7411
rect -3950 7391 -3930 7411
rect -3910 7391 -3890 7411
rect -3870 7391 -3850 7411
rect -3830 7391 -3810 7411
rect -3790 7391 -3770 7411
rect -3750 7391 -3730 7411
rect -3710 7391 -3690 7411
rect -3670 7391 -3650 7411
rect -3630 7391 -3610 7411
rect -3590 7391 -3570 7411
rect -3550 7391 -3530 7411
rect -3510 7391 -3490 7411
rect -3470 7391 -3450 7411
rect -3430 7391 -3410 7411
rect -3390 7391 -3370 7411
rect -3350 7391 -3330 7411
rect -3310 7391 -3290 7411
rect -3270 7391 -3250 7411
rect -3230 7391 -3210 7411
rect -3190 7391 -3165 7411
rect -5665 7376 -3165 7391
rect -5665 7329 -3165 7344
rect -5665 7309 -5650 7329
rect -5630 7309 -5610 7329
rect -5590 7309 -5570 7329
rect -5550 7309 -5530 7329
rect -5510 7309 -5490 7329
rect -5470 7309 -5450 7329
rect -5430 7309 -5410 7329
rect -5390 7309 -5370 7329
rect -5350 7309 -5330 7329
rect -5310 7309 -5290 7329
rect -5270 7309 -5250 7329
rect -5230 7309 -5210 7329
rect -5190 7309 -5170 7329
rect -5150 7309 -5130 7329
rect -5110 7309 -5090 7329
rect -5070 7309 -5050 7329
rect -5030 7309 -5010 7329
rect -4990 7309 -4970 7329
rect -4950 7309 -4930 7329
rect -4910 7309 -4890 7329
rect -4870 7309 -4850 7329
rect -4830 7309 -4810 7329
rect -4790 7309 -4770 7329
rect -4750 7309 -4730 7329
rect -4710 7309 -4690 7329
rect -4670 7309 -4650 7329
rect -4630 7309 -4610 7329
rect -4590 7309 -4570 7329
rect -4550 7309 -4530 7329
rect -4510 7309 -4490 7329
rect -4470 7309 -4450 7329
rect -4430 7309 -4410 7329
rect -4390 7309 -4370 7329
rect -4350 7309 -4330 7329
rect -4310 7309 -4290 7329
rect -4270 7309 -4250 7329
rect -4230 7309 -4210 7329
rect -4190 7309 -4170 7329
rect -4150 7309 -4130 7329
rect -4110 7309 -4090 7329
rect -4070 7309 -4050 7329
rect -4030 7309 -4010 7329
rect -3990 7309 -3970 7329
rect -3950 7309 -3930 7329
rect -3910 7309 -3890 7329
rect -3870 7309 -3850 7329
rect -3830 7309 -3810 7329
rect -3790 7309 -3770 7329
rect -3750 7309 -3730 7329
rect -3710 7309 -3690 7329
rect -3670 7309 -3650 7329
rect -3630 7309 -3610 7329
rect -3590 7309 -3570 7329
rect -3550 7309 -3530 7329
rect -3510 7309 -3490 7329
rect -3470 7309 -3450 7329
rect -3430 7309 -3410 7329
rect -3390 7309 -3370 7329
rect -3350 7309 -3330 7329
rect -3310 7309 -3290 7329
rect -3270 7309 -3250 7329
rect -3230 7309 -3210 7329
rect -3190 7309 -3165 7329
rect -5665 7294 -3165 7309
rect -5665 7247 -3165 7262
rect -5665 7227 -5650 7247
rect -5630 7227 -5610 7247
rect -5590 7227 -5570 7247
rect -5550 7227 -5530 7247
rect -5510 7227 -5490 7247
rect -5470 7227 -5450 7247
rect -5430 7227 -5410 7247
rect -5390 7227 -5370 7247
rect -5350 7227 -5330 7247
rect -5310 7227 -5290 7247
rect -5270 7227 -5250 7247
rect -5230 7227 -5210 7247
rect -5190 7227 -5170 7247
rect -5150 7227 -5130 7247
rect -5110 7227 -5090 7247
rect -5070 7227 -5050 7247
rect -5030 7227 -5010 7247
rect -4990 7227 -4970 7247
rect -4950 7227 -4930 7247
rect -4910 7227 -4890 7247
rect -4870 7227 -4850 7247
rect -4830 7227 -4810 7247
rect -4790 7227 -4770 7247
rect -4750 7227 -4730 7247
rect -4710 7227 -4690 7247
rect -4670 7227 -4650 7247
rect -4630 7227 -4610 7247
rect -4590 7227 -4570 7247
rect -4550 7227 -4530 7247
rect -4510 7227 -4490 7247
rect -4470 7227 -4450 7247
rect -4430 7227 -4410 7247
rect -4390 7227 -4370 7247
rect -4350 7227 -4330 7247
rect -4310 7227 -4290 7247
rect -4270 7227 -4250 7247
rect -4230 7227 -4210 7247
rect -4190 7227 -4170 7247
rect -4150 7227 -4130 7247
rect -4110 7227 -4090 7247
rect -4070 7227 -4050 7247
rect -4030 7227 -4010 7247
rect -3990 7227 -3970 7247
rect -3950 7227 -3930 7247
rect -3910 7227 -3890 7247
rect -3870 7227 -3850 7247
rect -3830 7227 -3810 7247
rect -3790 7227 -3770 7247
rect -3750 7227 -3730 7247
rect -3710 7227 -3690 7247
rect -3670 7227 -3650 7247
rect -3630 7227 -3610 7247
rect -3590 7227 -3570 7247
rect -3550 7227 -3530 7247
rect -3510 7227 -3490 7247
rect -3470 7227 -3450 7247
rect -3430 7227 -3410 7247
rect -3390 7227 -3370 7247
rect -3350 7227 -3330 7247
rect -3310 7227 -3290 7247
rect -3270 7227 -3250 7247
rect -3230 7227 -3210 7247
rect -3190 7227 -3165 7247
rect -5665 7212 -3165 7227
rect -5665 7165 -3165 7180
rect -5665 7145 -5650 7165
rect -5630 7145 -5610 7165
rect -5590 7145 -5570 7165
rect -5550 7145 -5530 7165
rect -5510 7145 -5490 7165
rect -5470 7145 -5450 7165
rect -5430 7145 -5410 7165
rect -5390 7145 -5370 7165
rect -5350 7145 -5330 7165
rect -5310 7145 -5290 7165
rect -5270 7145 -5250 7165
rect -5230 7145 -5210 7165
rect -5190 7145 -5170 7165
rect -5150 7145 -5130 7165
rect -5110 7145 -5090 7165
rect -5070 7145 -5050 7165
rect -5030 7145 -5010 7165
rect -4990 7145 -4970 7165
rect -4950 7145 -4930 7165
rect -4910 7145 -4890 7165
rect -4870 7145 -4850 7165
rect -4830 7145 -4810 7165
rect -4790 7145 -4770 7165
rect -4750 7145 -4730 7165
rect -4710 7145 -4690 7165
rect -4670 7145 -4650 7165
rect -4630 7145 -4610 7165
rect -4590 7145 -4570 7165
rect -4550 7145 -4530 7165
rect -4510 7145 -4490 7165
rect -4470 7145 -4450 7165
rect -4430 7145 -4410 7165
rect -4390 7145 -4370 7165
rect -4350 7145 -4330 7165
rect -4310 7145 -4290 7165
rect -4270 7145 -4250 7165
rect -4230 7145 -4210 7165
rect -4190 7145 -4170 7165
rect -4150 7145 -4130 7165
rect -4110 7145 -4090 7165
rect -4070 7145 -4050 7165
rect -4030 7145 -4010 7165
rect -3990 7145 -3970 7165
rect -3950 7145 -3930 7165
rect -3910 7145 -3890 7165
rect -3870 7145 -3850 7165
rect -3830 7145 -3810 7165
rect -3790 7145 -3770 7165
rect -3750 7145 -3730 7165
rect -3710 7145 -3690 7165
rect -3670 7145 -3650 7165
rect -3630 7145 -3610 7165
rect -3590 7145 -3570 7165
rect -3550 7145 -3530 7165
rect -3510 7145 -3490 7165
rect -3470 7145 -3450 7165
rect -3430 7145 -3410 7165
rect -3390 7145 -3370 7165
rect -3350 7145 -3330 7165
rect -3310 7145 -3290 7165
rect -3270 7145 -3250 7165
rect -3230 7145 -3210 7165
rect -3190 7145 -3165 7165
rect -5665 7130 -3165 7145
rect -5665 7083 -3165 7098
rect -5665 7063 -5650 7083
rect -5630 7063 -5610 7083
rect -5590 7063 -5570 7083
rect -5550 7063 -5530 7083
rect -5510 7063 -5490 7083
rect -5470 7063 -5450 7083
rect -5430 7063 -5410 7083
rect -5390 7063 -5370 7083
rect -5350 7063 -5330 7083
rect -5310 7063 -5290 7083
rect -5270 7063 -5250 7083
rect -5230 7063 -5210 7083
rect -5190 7063 -5170 7083
rect -5150 7063 -5130 7083
rect -5110 7063 -5090 7083
rect -5070 7063 -5050 7083
rect -5030 7063 -5010 7083
rect -4990 7063 -4970 7083
rect -4950 7063 -4930 7083
rect -4910 7063 -4890 7083
rect -4870 7063 -4850 7083
rect -4830 7063 -4810 7083
rect -4790 7063 -4770 7083
rect -4750 7063 -4730 7083
rect -4710 7063 -4690 7083
rect -4670 7063 -4650 7083
rect -4630 7063 -4610 7083
rect -4590 7063 -4570 7083
rect -4550 7063 -4530 7083
rect -4510 7063 -4490 7083
rect -4470 7063 -4450 7083
rect -4430 7063 -4410 7083
rect -4390 7063 -4370 7083
rect -4350 7063 -4330 7083
rect -4310 7063 -4290 7083
rect -4270 7063 -4250 7083
rect -4230 7063 -4210 7083
rect -4190 7063 -4170 7083
rect -4150 7063 -4130 7083
rect -4110 7063 -4090 7083
rect -4070 7063 -4050 7083
rect -4030 7063 -4010 7083
rect -3990 7063 -3970 7083
rect -3950 7063 -3930 7083
rect -3910 7063 -3890 7083
rect -3870 7063 -3850 7083
rect -3830 7063 -3810 7083
rect -3790 7063 -3770 7083
rect -3750 7063 -3730 7083
rect -3710 7063 -3690 7083
rect -3670 7063 -3650 7083
rect -3630 7063 -3610 7083
rect -3590 7063 -3570 7083
rect -3550 7063 -3530 7083
rect -3510 7063 -3490 7083
rect -3470 7063 -3450 7083
rect -3430 7063 -3410 7083
rect -3390 7063 -3370 7083
rect -3350 7063 -3330 7083
rect -3310 7063 -3290 7083
rect -3270 7063 -3250 7083
rect -3230 7063 -3210 7083
rect -3190 7063 -3165 7083
rect -5665 7048 -3165 7063
rect -5665 7001 -3165 7016
rect -5665 6981 -5650 7001
rect -5630 6981 -5610 7001
rect -5590 6981 -5570 7001
rect -5550 6981 -5530 7001
rect -5510 6981 -5490 7001
rect -5470 6981 -5450 7001
rect -5430 6981 -5410 7001
rect -5390 6981 -5370 7001
rect -5350 6981 -5330 7001
rect -5310 6981 -5290 7001
rect -5270 6981 -5250 7001
rect -5230 6981 -5210 7001
rect -5190 6981 -5170 7001
rect -5150 6981 -5130 7001
rect -5110 6981 -5090 7001
rect -5070 6981 -5050 7001
rect -5030 6981 -5010 7001
rect -4990 6981 -4970 7001
rect -4950 6981 -4930 7001
rect -4910 6981 -4890 7001
rect -4870 6981 -4850 7001
rect -4830 6981 -4810 7001
rect -4790 6981 -4770 7001
rect -4750 6981 -4730 7001
rect -4710 6981 -4690 7001
rect -4670 6981 -4650 7001
rect -4630 6981 -4610 7001
rect -4590 6981 -4570 7001
rect -4550 6981 -4530 7001
rect -4510 6981 -4490 7001
rect -4470 6981 -4450 7001
rect -4430 6981 -4410 7001
rect -4390 6981 -4370 7001
rect -4350 6981 -4330 7001
rect -4310 6981 -4290 7001
rect -4270 6981 -4250 7001
rect -4230 6981 -4210 7001
rect -4190 6981 -4170 7001
rect -4150 6981 -4130 7001
rect -4110 6981 -4090 7001
rect -4070 6981 -4050 7001
rect -4030 6981 -4010 7001
rect -3990 6981 -3970 7001
rect -3950 6981 -3930 7001
rect -3910 6981 -3890 7001
rect -3870 6981 -3850 7001
rect -3830 6981 -3810 7001
rect -3790 6981 -3770 7001
rect -3750 6981 -3730 7001
rect -3710 6981 -3690 7001
rect -3670 6981 -3650 7001
rect -3630 6981 -3610 7001
rect -3590 6981 -3570 7001
rect -3550 6981 -3530 7001
rect -3510 6981 -3490 7001
rect -3470 6981 -3450 7001
rect -3430 6981 -3410 7001
rect -3390 6981 -3370 7001
rect -3350 6981 -3330 7001
rect -3310 6981 -3290 7001
rect -3270 6981 -3250 7001
rect -3230 6981 -3210 7001
rect -3190 6981 -3165 7001
rect -5665 6966 -3165 6981
rect -5665 6919 -3165 6934
rect -5665 6899 -5650 6919
rect -5630 6899 -5610 6919
rect -5590 6899 -5570 6919
rect -5550 6899 -5530 6919
rect -5510 6899 -5490 6919
rect -5470 6899 -5450 6919
rect -5430 6899 -5410 6919
rect -5390 6899 -5370 6919
rect -5350 6899 -5330 6919
rect -5310 6899 -5290 6919
rect -5270 6899 -5250 6919
rect -5230 6899 -5210 6919
rect -5190 6899 -5170 6919
rect -5150 6899 -5130 6919
rect -5110 6899 -5090 6919
rect -5070 6899 -5050 6919
rect -5030 6899 -5010 6919
rect -4990 6899 -4970 6919
rect -4950 6899 -4930 6919
rect -4910 6899 -4890 6919
rect -4870 6899 -4850 6919
rect -4830 6899 -4810 6919
rect -4790 6899 -4770 6919
rect -4750 6899 -4730 6919
rect -4710 6899 -4690 6919
rect -4670 6899 -4650 6919
rect -4630 6899 -4610 6919
rect -4590 6899 -4570 6919
rect -4550 6899 -4530 6919
rect -4510 6899 -4490 6919
rect -4470 6899 -4450 6919
rect -4430 6899 -4410 6919
rect -4390 6899 -4370 6919
rect -4350 6899 -4330 6919
rect -4310 6899 -4290 6919
rect -4270 6899 -4250 6919
rect -4230 6899 -4210 6919
rect -4190 6899 -4170 6919
rect -4150 6899 -4130 6919
rect -4110 6899 -4090 6919
rect -4070 6899 -4050 6919
rect -4030 6899 -4010 6919
rect -3990 6899 -3970 6919
rect -3950 6899 -3930 6919
rect -3910 6899 -3890 6919
rect -3870 6899 -3850 6919
rect -3830 6899 -3810 6919
rect -3790 6899 -3770 6919
rect -3750 6899 -3730 6919
rect -3710 6899 -3690 6919
rect -3670 6899 -3650 6919
rect -3630 6899 -3610 6919
rect -3590 6899 -3570 6919
rect -3550 6899 -3530 6919
rect -3510 6899 -3490 6919
rect -3470 6899 -3450 6919
rect -3430 6899 -3410 6919
rect -3390 6899 -3370 6919
rect -3350 6899 -3330 6919
rect -3310 6899 -3290 6919
rect -3270 6899 -3250 6919
rect -3230 6899 -3210 6919
rect -3190 6899 -3165 6919
rect -5665 6884 -3165 6899
rect -5665 6837 -3165 6852
rect -5665 6817 -5650 6837
rect -5630 6817 -5610 6837
rect -5590 6817 -5570 6837
rect -5550 6817 -5530 6837
rect -5510 6817 -5490 6837
rect -5470 6817 -5450 6837
rect -5430 6817 -5410 6837
rect -5390 6817 -5370 6837
rect -5350 6817 -5330 6837
rect -5310 6817 -5290 6837
rect -5270 6817 -5250 6837
rect -5230 6817 -5210 6837
rect -5190 6817 -5170 6837
rect -5150 6817 -5130 6837
rect -5110 6817 -5090 6837
rect -5070 6817 -5050 6837
rect -5030 6817 -5010 6837
rect -4990 6817 -4970 6837
rect -4950 6817 -4930 6837
rect -4910 6817 -4890 6837
rect -4870 6817 -4850 6837
rect -4830 6817 -4810 6837
rect -4790 6817 -4770 6837
rect -4750 6817 -4730 6837
rect -4710 6817 -4690 6837
rect -4670 6817 -4650 6837
rect -4630 6817 -4610 6837
rect -4590 6817 -4570 6837
rect -4550 6817 -4530 6837
rect -4510 6817 -4490 6837
rect -4470 6817 -4450 6837
rect -4430 6817 -4410 6837
rect -4390 6817 -4370 6837
rect -4350 6817 -4330 6837
rect -4310 6817 -4290 6837
rect -4270 6817 -4250 6837
rect -4230 6817 -4210 6837
rect -4190 6817 -4170 6837
rect -4150 6817 -4130 6837
rect -4110 6817 -4090 6837
rect -4070 6817 -4050 6837
rect -4030 6817 -4010 6837
rect -3990 6817 -3970 6837
rect -3950 6817 -3930 6837
rect -3910 6817 -3890 6837
rect -3870 6817 -3850 6837
rect -3830 6817 -3810 6837
rect -3790 6817 -3770 6837
rect -3750 6817 -3730 6837
rect -3710 6817 -3690 6837
rect -3670 6817 -3650 6837
rect -3630 6817 -3610 6837
rect -3590 6817 -3570 6837
rect -3550 6817 -3530 6837
rect -3510 6817 -3490 6837
rect -3470 6817 -3450 6837
rect -3430 6817 -3410 6837
rect -3390 6817 -3370 6837
rect -3350 6817 -3330 6837
rect -3310 6817 -3290 6837
rect -3270 6817 -3250 6837
rect -3230 6817 -3210 6837
rect -3190 6817 -3165 6837
rect -5665 6802 -3165 6817
rect -5665 6755 -3165 6770
rect -5665 6735 -5650 6755
rect -5630 6735 -5610 6755
rect -5590 6735 -5570 6755
rect -5550 6735 -5530 6755
rect -5510 6735 -5490 6755
rect -5470 6735 -5450 6755
rect -5430 6735 -5410 6755
rect -5390 6735 -5370 6755
rect -5350 6735 -5330 6755
rect -5310 6735 -5290 6755
rect -5270 6735 -5250 6755
rect -5230 6735 -5210 6755
rect -5190 6735 -5170 6755
rect -5150 6735 -5130 6755
rect -5110 6735 -5090 6755
rect -5070 6735 -5050 6755
rect -5030 6735 -5010 6755
rect -4990 6735 -4970 6755
rect -4950 6735 -4930 6755
rect -4910 6735 -4890 6755
rect -4870 6735 -4850 6755
rect -4830 6735 -4810 6755
rect -4790 6735 -4770 6755
rect -4750 6735 -4730 6755
rect -4710 6735 -4690 6755
rect -4670 6735 -4650 6755
rect -4630 6735 -4610 6755
rect -4590 6735 -4570 6755
rect -4550 6735 -4530 6755
rect -4510 6735 -4490 6755
rect -4470 6735 -4450 6755
rect -4430 6735 -4410 6755
rect -4390 6735 -4370 6755
rect -4350 6735 -4330 6755
rect -4310 6735 -4290 6755
rect -4270 6735 -4250 6755
rect -4230 6735 -4210 6755
rect -4190 6735 -4170 6755
rect -4150 6735 -4130 6755
rect -4110 6735 -4090 6755
rect -4070 6735 -4050 6755
rect -4030 6735 -4010 6755
rect -3990 6735 -3970 6755
rect -3950 6735 -3930 6755
rect -3910 6735 -3890 6755
rect -3870 6735 -3850 6755
rect -3830 6735 -3810 6755
rect -3790 6735 -3770 6755
rect -3750 6735 -3730 6755
rect -3710 6735 -3690 6755
rect -3670 6735 -3650 6755
rect -3630 6735 -3610 6755
rect -3590 6735 -3570 6755
rect -3550 6735 -3530 6755
rect -3510 6735 -3490 6755
rect -3470 6735 -3450 6755
rect -3430 6735 -3410 6755
rect -3390 6735 -3370 6755
rect -3350 6735 -3330 6755
rect -3310 6735 -3290 6755
rect -3270 6735 -3250 6755
rect -3230 6735 -3210 6755
rect -3190 6735 -3165 6755
rect -5665 6720 -3165 6735
rect -5665 6673 -3165 6688
rect -5665 6653 -5650 6673
rect -5630 6653 -5610 6673
rect -5590 6653 -5570 6673
rect -5550 6653 -5530 6673
rect -5510 6653 -5490 6673
rect -5470 6653 -5450 6673
rect -5430 6653 -5410 6673
rect -5390 6653 -5370 6673
rect -5350 6653 -5330 6673
rect -5310 6653 -5290 6673
rect -5270 6653 -5250 6673
rect -5230 6653 -5210 6673
rect -5190 6653 -5170 6673
rect -5150 6653 -5130 6673
rect -5110 6653 -5090 6673
rect -5070 6653 -5050 6673
rect -5030 6653 -5010 6673
rect -4990 6653 -4970 6673
rect -4950 6653 -4930 6673
rect -4910 6653 -4890 6673
rect -4870 6653 -4850 6673
rect -4830 6653 -4810 6673
rect -4790 6653 -4770 6673
rect -4750 6653 -4730 6673
rect -4710 6653 -4690 6673
rect -4670 6653 -4650 6673
rect -4630 6653 -4610 6673
rect -4590 6653 -4570 6673
rect -4550 6653 -4530 6673
rect -4510 6653 -4490 6673
rect -4470 6653 -4450 6673
rect -4430 6653 -4410 6673
rect -4390 6653 -4370 6673
rect -4350 6653 -4330 6673
rect -4310 6653 -4290 6673
rect -4270 6653 -4250 6673
rect -4230 6653 -4210 6673
rect -4190 6653 -4170 6673
rect -4150 6653 -4130 6673
rect -4110 6653 -4090 6673
rect -4070 6653 -4050 6673
rect -4030 6653 -4010 6673
rect -3990 6653 -3970 6673
rect -3950 6653 -3930 6673
rect -3910 6653 -3890 6673
rect -3870 6653 -3850 6673
rect -3830 6653 -3810 6673
rect -3790 6653 -3770 6673
rect -3750 6653 -3730 6673
rect -3710 6653 -3690 6673
rect -3670 6653 -3650 6673
rect -3630 6653 -3610 6673
rect -3590 6653 -3570 6673
rect -3550 6653 -3530 6673
rect -3510 6653 -3490 6673
rect -3470 6653 -3450 6673
rect -3430 6653 -3410 6673
rect -3390 6653 -3370 6673
rect -3350 6653 -3330 6673
rect -3310 6653 -3290 6673
rect -3270 6653 -3250 6673
rect -3230 6653 -3210 6673
rect -3190 6653 -3165 6673
rect -5665 6638 -3165 6653
rect -5665 6591 -3165 6606
rect -5665 6571 -5650 6591
rect -5630 6571 -5610 6591
rect -5590 6571 -5570 6591
rect -5550 6571 -5530 6591
rect -5510 6571 -5490 6591
rect -5470 6571 -5450 6591
rect -5430 6571 -5410 6591
rect -5390 6571 -5370 6591
rect -5350 6571 -5330 6591
rect -5310 6571 -5290 6591
rect -5270 6571 -5250 6591
rect -5230 6571 -5210 6591
rect -5190 6571 -5170 6591
rect -5150 6571 -5130 6591
rect -5110 6571 -5090 6591
rect -5070 6571 -5050 6591
rect -5030 6571 -5010 6591
rect -4990 6571 -4970 6591
rect -4950 6571 -4930 6591
rect -4910 6571 -4890 6591
rect -4870 6571 -4850 6591
rect -4830 6571 -4810 6591
rect -4790 6571 -4770 6591
rect -4750 6571 -4730 6591
rect -4710 6571 -4690 6591
rect -4670 6571 -4650 6591
rect -4630 6571 -4610 6591
rect -4590 6571 -4570 6591
rect -4550 6571 -4530 6591
rect -4510 6571 -4490 6591
rect -4470 6571 -4450 6591
rect -4430 6571 -4410 6591
rect -4390 6571 -4370 6591
rect -4350 6571 -4330 6591
rect -4310 6571 -4290 6591
rect -4270 6571 -4250 6591
rect -4230 6571 -4210 6591
rect -4190 6571 -4170 6591
rect -4150 6571 -4130 6591
rect -4110 6571 -4090 6591
rect -4070 6571 -4050 6591
rect -4030 6571 -4010 6591
rect -3990 6571 -3970 6591
rect -3950 6571 -3930 6591
rect -3910 6571 -3890 6591
rect -3870 6571 -3850 6591
rect -3830 6571 -3810 6591
rect -3790 6571 -3770 6591
rect -3750 6571 -3730 6591
rect -3710 6571 -3690 6591
rect -3670 6571 -3650 6591
rect -3630 6571 -3610 6591
rect -3590 6571 -3570 6591
rect -3550 6571 -3530 6591
rect -3510 6571 -3490 6591
rect -3470 6571 -3450 6591
rect -3430 6571 -3410 6591
rect -3390 6571 -3370 6591
rect -3350 6571 -3330 6591
rect -3310 6571 -3290 6591
rect -3270 6571 -3250 6591
rect -3230 6571 -3210 6591
rect -3190 6571 -3165 6591
rect -5665 6556 -3165 6571
rect -5665 6509 -3165 6524
rect -5665 6489 -5650 6509
rect -5630 6489 -5610 6509
rect -5590 6489 -5570 6509
rect -5550 6489 -5530 6509
rect -5510 6489 -5490 6509
rect -5470 6489 -5450 6509
rect -5430 6489 -5410 6509
rect -5390 6489 -5370 6509
rect -5350 6489 -5330 6509
rect -5310 6489 -5290 6509
rect -5270 6489 -5250 6509
rect -5230 6489 -5210 6509
rect -5190 6489 -5170 6509
rect -5150 6489 -5130 6509
rect -5110 6489 -5090 6509
rect -5070 6489 -5050 6509
rect -5030 6489 -5010 6509
rect -4990 6489 -4970 6509
rect -4950 6489 -4930 6509
rect -4910 6489 -4890 6509
rect -4870 6489 -4850 6509
rect -4830 6489 -4810 6509
rect -4790 6489 -4770 6509
rect -4750 6489 -4730 6509
rect -4710 6489 -4690 6509
rect -4670 6489 -4650 6509
rect -4630 6489 -4610 6509
rect -4590 6489 -4570 6509
rect -4550 6489 -4530 6509
rect -4510 6489 -4490 6509
rect -4470 6489 -4450 6509
rect -4430 6489 -4410 6509
rect -4390 6489 -4370 6509
rect -4350 6489 -4330 6509
rect -4310 6489 -4290 6509
rect -4270 6489 -4250 6509
rect -4230 6489 -4210 6509
rect -4190 6489 -4170 6509
rect -4150 6489 -4130 6509
rect -4110 6489 -4090 6509
rect -4070 6489 -4050 6509
rect -4030 6489 -4010 6509
rect -3990 6489 -3970 6509
rect -3950 6489 -3930 6509
rect -3910 6489 -3890 6509
rect -3870 6489 -3850 6509
rect -3830 6489 -3810 6509
rect -3790 6489 -3770 6509
rect -3750 6489 -3730 6509
rect -3710 6489 -3690 6509
rect -3670 6489 -3650 6509
rect -3630 6489 -3610 6509
rect -3590 6489 -3570 6509
rect -3550 6489 -3530 6509
rect -3510 6489 -3490 6509
rect -3470 6489 -3450 6509
rect -3430 6489 -3410 6509
rect -3390 6489 -3370 6509
rect -3350 6489 -3330 6509
rect -3310 6489 -3290 6509
rect -3270 6489 -3250 6509
rect -3230 6489 -3210 6509
rect -3190 6489 -3165 6509
rect -5665 6474 -3165 6489
rect -5665 6427 -3165 6442
rect -5665 6407 -5650 6427
rect -5630 6407 -5610 6427
rect -5590 6407 -5570 6427
rect -5550 6407 -5530 6427
rect -5510 6407 -5490 6427
rect -5470 6407 -5450 6427
rect -5430 6407 -5410 6427
rect -5390 6407 -5370 6427
rect -5350 6407 -5330 6427
rect -5310 6407 -5290 6427
rect -5270 6407 -5250 6427
rect -5230 6407 -5210 6427
rect -5190 6407 -5170 6427
rect -5150 6407 -5130 6427
rect -5110 6407 -5090 6427
rect -5070 6407 -5050 6427
rect -5030 6407 -5010 6427
rect -4990 6407 -4970 6427
rect -4950 6407 -4930 6427
rect -4910 6407 -4890 6427
rect -4870 6407 -4850 6427
rect -4830 6407 -4810 6427
rect -4790 6407 -4770 6427
rect -4750 6407 -4730 6427
rect -4710 6407 -4690 6427
rect -4670 6407 -4650 6427
rect -4630 6407 -4610 6427
rect -4590 6407 -4570 6427
rect -4550 6407 -4530 6427
rect -4510 6407 -4490 6427
rect -4470 6407 -4450 6427
rect -4430 6407 -4410 6427
rect -4390 6407 -4370 6427
rect -4350 6407 -4330 6427
rect -4310 6407 -4290 6427
rect -4270 6407 -4250 6427
rect -4230 6407 -4210 6427
rect -4190 6407 -4170 6427
rect -4150 6407 -4130 6427
rect -4110 6407 -4090 6427
rect -4070 6407 -4050 6427
rect -4030 6407 -4010 6427
rect -3990 6407 -3970 6427
rect -3950 6407 -3930 6427
rect -3910 6407 -3890 6427
rect -3870 6407 -3850 6427
rect -3830 6407 -3810 6427
rect -3790 6407 -3770 6427
rect -3750 6407 -3730 6427
rect -3710 6407 -3690 6427
rect -3670 6407 -3650 6427
rect -3630 6407 -3610 6427
rect -3590 6407 -3570 6427
rect -3550 6407 -3530 6427
rect -3510 6407 -3490 6427
rect -3470 6407 -3450 6427
rect -3430 6407 -3410 6427
rect -3390 6407 -3370 6427
rect -3350 6407 -3330 6427
rect -3310 6407 -3290 6427
rect -3270 6407 -3250 6427
rect -3230 6407 -3210 6427
rect -3190 6407 -3165 6427
rect -5665 6392 -3165 6407
rect -5665 6345 -3165 6360
rect -5665 6325 -5650 6345
rect -5630 6325 -5610 6345
rect -5590 6325 -5570 6345
rect -5550 6325 -5530 6345
rect -5510 6325 -5490 6345
rect -5470 6325 -5450 6345
rect -5430 6325 -5410 6345
rect -5390 6325 -5370 6345
rect -5350 6325 -5330 6345
rect -5310 6325 -5290 6345
rect -5270 6325 -5250 6345
rect -5230 6325 -5210 6345
rect -5190 6325 -5170 6345
rect -5150 6325 -5130 6345
rect -5110 6325 -5090 6345
rect -5070 6325 -5050 6345
rect -5030 6325 -5010 6345
rect -4990 6325 -4970 6345
rect -4950 6325 -4930 6345
rect -4910 6325 -4890 6345
rect -4870 6325 -4850 6345
rect -4830 6325 -4810 6345
rect -4790 6325 -4770 6345
rect -4750 6325 -4730 6345
rect -4710 6325 -4690 6345
rect -4670 6325 -4650 6345
rect -4630 6325 -4610 6345
rect -4590 6325 -4570 6345
rect -4550 6325 -4530 6345
rect -4510 6325 -4490 6345
rect -4470 6325 -4450 6345
rect -4430 6325 -4410 6345
rect -4390 6325 -4370 6345
rect -4350 6325 -4330 6345
rect -4310 6325 -4290 6345
rect -4270 6325 -4250 6345
rect -4230 6325 -4210 6345
rect -4190 6325 -4170 6345
rect -4150 6325 -4130 6345
rect -4110 6325 -4090 6345
rect -4070 6325 -4050 6345
rect -4030 6325 -4010 6345
rect -3990 6325 -3970 6345
rect -3950 6325 -3930 6345
rect -3910 6325 -3890 6345
rect -3870 6325 -3850 6345
rect -3830 6325 -3810 6345
rect -3790 6325 -3770 6345
rect -3750 6325 -3730 6345
rect -3710 6325 -3690 6345
rect -3670 6325 -3650 6345
rect -3630 6325 -3610 6345
rect -3590 6325 -3570 6345
rect -3550 6325 -3530 6345
rect -3510 6325 -3490 6345
rect -3470 6325 -3450 6345
rect -3430 6325 -3410 6345
rect -3390 6325 -3370 6345
rect -3350 6325 -3330 6345
rect -3310 6325 -3290 6345
rect -3270 6325 -3250 6345
rect -3230 6325 -3210 6345
rect -3190 6325 -3165 6345
rect -5665 6315 -3165 6325
rect -1975 8477 525 8490
rect -1975 8457 -1950 8477
rect -1930 8457 -1910 8477
rect -1890 8457 -1870 8477
rect -1850 8457 -1830 8477
rect -1810 8457 -1790 8477
rect -1770 8457 -1750 8477
rect -1730 8457 -1710 8477
rect -1690 8457 -1670 8477
rect -1650 8457 -1630 8477
rect -1610 8457 -1590 8477
rect -1570 8457 -1550 8477
rect -1530 8457 -1510 8477
rect -1490 8457 -1470 8477
rect -1450 8457 -1430 8477
rect -1410 8457 -1390 8477
rect -1370 8457 -1350 8477
rect -1330 8457 -1310 8477
rect -1290 8457 -1270 8477
rect -1250 8457 -1230 8477
rect -1210 8457 -1190 8477
rect -1170 8457 -1150 8477
rect -1130 8457 -1110 8477
rect -1090 8457 -1070 8477
rect -1050 8457 -1030 8477
rect -1010 8457 -990 8477
rect -970 8457 -950 8477
rect -930 8457 -910 8477
rect -890 8457 -870 8477
rect -850 8457 -830 8477
rect -810 8457 -790 8477
rect -770 8457 -750 8477
rect -730 8457 -710 8477
rect -690 8457 -670 8477
rect -650 8457 -630 8477
rect -610 8457 -590 8477
rect -570 8457 -550 8477
rect -530 8457 -510 8477
rect -490 8457 -470 8477
rect -450 8457 -430 8477
rect -410 8457 -390 8477
rect -370 8457 -350 8477
rect -330 8457 -310 8477
rect -290 8457 -270 8477
rect -250 8457 -230 8477
rect -210 8457 -190 8477
rect -170 8457 -150 8477
rect -130 8457 -110 8477
rect -90 8457 -70 8477
rect -50 8457 -30 8477
rect -10 8457 10 8477
rect 30 8457 50 8477
rect 70 8457 90 8477
rect 110 8457 130 8477
rect 150 8457 170 8477
rect 190 8457 210 8477
rect 230 8457 250 8477
rect 270 8457 290 8477
rect 310 8457 330 8477
rect 350 8457 370 8477
rect 390 8457 410 8477
rect 430 8457 450 8477
rect 470 8457 490 8477
rect 510 8457 525 8477
rect -1975 8442 525 8457
rect -1975 8395 525 8410
rect -1975 8375 -1950 8395
rect -1930 8375 -1910 8395
rect -1890 8375 -1870 8395
rect -1850 8375 -1830 8395
rect -1810 8375 -1790 8395
rect -1770 8375 -1750 8395
rect -1730 8375 -1710 8395
rect -1690 8375 -1670 8395
rect -1650 8375 -1630 8395
rect -1610 8375 -1590 8395
rect -1570 8375 -1550 8395
rect -1530 8375 -1510 8395
rect -1490 8375 -1470 8395
rect -1450 8375 -1430 8395
rect -1410 8375 -1390 8395
rect -1370 8375 -1350 8395
rect -1330 8375 -1310 8395
rect -1290 8375 -1270 8395
rect -1250 8375 -1230 8395
rect -1210 8375 -1190 8395
rect -1170 8375 -1150 8395
rect -1130 8375 -1110 8395
rect -1090 8375 -1070 8395
rect -1050 8375 -1030 8395
rect -1010 8375 -990 8395
rect -970 8375 -950 8395
rect -930 8375 -910 8395
rect -890 8375 -870 8395
rect -850 8375 -830 8395
rect -810 8375 -790 8395
rect -770 8375 -750 8395
rect -730 8375 -710 8395
rect -690 8375 -670 8395
rect -650 8375 -630 8395
rect -610 8375 -590 8395
rect -570 8375 -550 8395
rect -530 8375 -510 8395
rect -490 8375 -470 8395
rect -450 8375 -430 8395
rect -410 8375 -390 8395
rect -370 8375 -350 8395
rect -330 8375 -310 8395
rect -290 8375 -270 8395
rect -250 8375 -230 8395
rect -210 8375 -190 8395
rect -170 8375 -150 8395
rect -130 8375 -110 8395
rect -90 8375 -70 8395
rect -50 8375 -30 8395
rect -10 8375 10 8395
rect 30 8375 50 8395
rect 70 8375 90 8395
rect 110 8375 130 8395
rect 150 8375 170 8395
rect 190 8375 210 8395
rect 230 8375 250 8395
rect 270 8375 290 8395
rect 310 8375 330 8395
rect 350 8375 370 8395
rect 390 8375 410 8395
rect 430 8375 450 8395
rect 470 8375 490 8395
rect 510 8375 525 8395
rect -1975 8360 525 8375
rect -1975 8313 525 8328
rect -1975 8293 -1950 8313
rect -1930 8293 -1910 8313
rect -1890 8293 -1870 8313
rect -1850 8293 -1830 8313
rect -1810 8293 -1790 8313
rect -1770 8293 -1750 8313
rect -1730 8293 -1710 8313
rect -1690 8293 -1670 8313
rect -1650 8293 -1630 8313
rect -1610 8293 -1590 8313
rect -1570 8293 -1550 8313
rect -1530 8293 -1510 8313
rect -1490 8293 -1470 8313
rect -1450 8293 -1430 8313
rect -1410 8293 -1390 8313
rect -1370 8293 -1350 8313
rect -1330 8293 -1310 8313
rect -1290 8293 -1270 8313
rect -1250 8293 -1230 8313
rect -1210 8293 -1190 8313
rect -1170 8293 -1150 8313
rect -1130 8293 -1110 8313
rect -1090 8293 -1070 8313
rect -1050 8293 -1030 8313
rect -1010 8293 -990 8313
rect -970 8293 -950 8313
rect -930 8293 -910 8313
rect -890 8293 -870 8313
rect -850 8293 -830 8313
rect -810 8293 -790 8313
rect -770 8293 -750 8313
rect -730 8293 -710 8313
rect -690 8293 -670 8313
rect -650 8293 -630 8313
rect -610 8293 -590 8313
rect -570 8293 -550 8313
rect -530 8293 -510 8313
rect -490 8293 -470 8313
rect -450 8293 -430 8313
rect -410 8293 -390 8313
rect -370 8293 -350 8313
rect -330 8293 -310 8313
rect -290 8293 -270 8313
rect -250 8293 -230 8313
rect -210 8293 -190 8313
rect -170 8293 -150 8313
rect -130 8293 -110 8313
rect -90 8293 -70 8313
rect -50 8293 -30 8313
rect -10 8293 10 8313
rect 30 8293 50 8313
rect 70 8293 90 8313
rect 110 8293 130 8313
rect 150 8293 170 8313
rect 190 8293 210 8313
rect 230 8293 250 8313
rect 270 8293 290 8313
rect 310 8293 330 8313
rect 350 8293 370 8313
rect 390 8293 410 8313
rect 430 8293 450 8313
rect 470 8293 490 8313
rect 510 8293 525 8313
rect -1975 8278 525 8293
rect -1975 8231 525 8246
rect -1975 8211 -1950 8231
rect -1930 8211 -1910 8231
rect -1890 8211 -1870 8231
rect -1850 8211 -1830 8231
rect -1810 8211 -1790 8231
rect -1770 8211 -1750 8231
rect -1730 8211 -1710 8231
rect -1690 8211 -1670 8231
rect -1650 8211 -1630 8231
rect -1610 8211 -1590 8231
rect -1570 8211 -1550 8231
rect -1530 8211 -1510 8231
rect -1490 8211 -1470 8231
rect -1450 8211 -1430 8231
rect -1410 8211 -1390 8231
rect -1370 8211 -1350 8231
rect -1330 8211 -1310 8231
rect -1290 8211 -1270 8231
rect -1250 8211 -1230 8231
rect -1210 8211 -1190 8231
rect -1170 8211 -1150 8231
rect -1130 8211 -1110 8231
rect -1090 8211 -1070 8231
rect -1050 8211 -1030 8231
rect -1010 8211 -990 8231
rect -970 8211 -950 8231
rect -930 8211 -910 8231
rect -890 8211 -870 8231
rect -850 8211 -830 8231
rect -810 8211 -790 8231
rect -770 8211 -750 8231
rect -730 8211 -710 8231
rect -690 8211 -670 8231
rect -650 8211 -630 8231
rect -610 8211 -590 8231
rect -570 8211 -550 8231
rect -530 8211 -510 8231
rect -490 8211 -470 8231
rect -450 8211 -430 8231
rect -410 8211 -390 8231
rect -370 8211 -350 8231
rect -330 8211 -310 8231
rect -290 8211 -270 8231
rect -250 8211 -230 8231
rect -210 8211 -190 8231
rect -170 8211 -150 8231
rect -130 8211 -110 8231
rect -90 8211 -70 8231
rect -50 8211 -30 8231
rect -10 8211 10 8231
rect 30 8211 50 8231
rect 70 8211 90 8231
rect 110 8211 130 8231
rect 150 8211 170 8231
rect 190 8211 210 8231
rect 230 8211 250 8231
rect 270 8211 290 8231
rect 310 8211 330 8231
rect 350 8211 370 8231
rect 390 8211 410 8231
rect 430 8211 450 8231
rect 470 8211 490 8231
rect 510 8211 525 8231
rect -1975 8196 525 8211
rect -1975 8149 525 8164
rect -1975 8129 -1950 8149
rect -1930 8129 -1910 8149
rect -1890 8129 -1870 8149
rect -1850 8129 -1830 8149
rect -1810 8129 -1790 8149
rect -1770 8129 -1750 8149
rect -1730 8129 -1710 8149
rect -1690 8129 -1670 8149
rect -1650 8129 -1630 8149
rect -1610 8129 -1590 8149
rect -1570 8129 -1550 8149
rect -1530 8129 -1510 8149
rect -1490 8129 -1470 8149
rect -1450 8129 -1430 8149
rect -1410 8129 -1390 8149
rect -1370 8129 -1350 8149
rect -1330 8129 -1310 8149
rect -1290 8129 -1270 8149
rect -1250 8129 -1230 8149
rect -1210 8129 -1190 8149
rect -1170 8129 -1150 8149
rect -1130 8129 -1110 8149
rect -1090 8129 -1070 8149
rect -1050 8129 -1030 8149
rect -1010 8129 -990 8149
rect -970 8129 -950 8149
rect -930 8129 -910 8149
rect -890 8129 -870 8149
rect -850 8129 -830 8149
rect -810 8129 -790 8149
rect -770 8129 -750 8149
rect -730 8129 -710 8149
rect -690 8129 -670 8149
rect -650 8129 -630 8149
rect -610 8129 -590 8149
rect -570 8129 -550 8149
rect -530 8129 -510 8149
rect -490 8129 -470 8149
rect -450 8129 -430 8149
rect -410 8129 -390 8149
rect -370 8129 -350 8149
rect -330 8129 -310 8149
rect -290 8129 -270 8149
rect -250 8129 -230 8149
rect -210 8129 -190 8149
rect -170 8129 -150 8149
rect -130 8129 -110 8149
rect -90 8129 -70 8149
rect -50 8129 -30 8149
rect -10 8129 10 8149
rect 30 8129 50 8149
rect 70 8129 90 8149
rect 110 8129 130 8149
rect 150 8129 170 8149
rect 190 8129 210 8149
rect 230 8129 250 8149
rect 270 8129 290 8149
rect 310 8129 330 8149
rect 350 8129 370 8149
rect 390 8129 410 8149
rect 430 8129 450 8149
rect 470 8129 490 8149
rect 510 8129 525 8149
rect -1975 8114 525 8129
rect -1975 8067 525 8082
rect -1975 8047 -1950 8067
rect -1930 8047 -1910 8067
rect -1890 8047 -1870 8067
rect -1850 8047 -1830 8067
rect -1810 8047 -1790 8067
rect -1770 8047 -1750 8067
rect -1730 8047 -1710 8067
rect -1690 8047 -1670 8067
rect -1650 8047 -1630 8067
rect -1610 8047 -1590 8067
rect -1570 8047 -1550 8067
rect -1530 8047 -1510 8067
rect -1490 8047 -1470 8067
rect -1450 8047 -1430 8067
rect -1410 8047 -1390 8067
rect -1370 8047 -1350 8067
rect -1330 8047 -1310 8067
rect -1290 8047 -1270 8067
rect -1250 8047 -1230 8067
rect -1210 8047 -1190 8067
rect -1170 8047 -1150 8067
rect -1130 8047 -1110 8067
rect -1090 8047 -1070 8067
rect -1050 8047 -1030 8067
rect -1010 8047 -990 8067
rect -970 8047 -950 8067
rect -930 8047 -910 8067
rect -890 8047 -870 8067
rect -850 8047 -830 8067
rect -810 8047 -790 8067
rect -770 8047 -750 8067
rect -730 8047 -710 8067
rect -690 8047 -670 8067
rect -650 8047 -630 8067
rect -610 8047 -590 8067
rect -570 8047 -550 8067
rect -530 8047 -510 8067
rect -490 8047 -470 8067
rect -450 8047 -430 8067
rect -410 8047 -390 8067
rect -370 8047 -350 8067
rect -330 8047 -310 8067
rect -290 8047 -270 8067
rect -250 8047 -230 8067
rect -210 8047 -190 8067
rect -170 8047 -150 8067
rect -130 8047 -110 8067
rect -90 8047 -70 8067
rect -50 8047 -30 8067
rect -10 8047 10 8067
rect 30 8047 50 8067
rect 70 8047 90 8067
rect 110 8047 130 8067
rect 150 8047 170 8067
rect 190 8047 210 8067
rect 230 8047 250 8067
rect 270 8047 290 8067
rect 310 8047 330 8067
rect 350 8047 370 8067
rect 390 8047 410 8067
rect 430 8047 450 8067
rect 470 8047 490 8067
rect 510 8047 525 8067
rect -1975 8032 525 8047
rect -1975 7985 525 8000
rect -1975 7965 -1950 7985
rect -1930 7965 -1910 7985
rect -1890 7965 -1870 7985
rect -1850 7965 -1830 7985
rect -1810 7965 -1790 7985
rect -1770 7965 -1750 7985
rect -1730 7965 -1710 7985
rect -1690 7965 -1670 7985
rect -1650 7965 -1630 7985
rect -1610 7965 -1590 7985
rect -1570 7965 -1550 7985
rect -1530 7965 -1510 7985
rect -1490 7965 -1470 7985
rect -1450 7965 -1430 7985
rect -1410 7965 -1390 7985
rect -1370 7965 -1350 7985
rect -1330 7965 -1310 7985
rect -1290 7965 -1270 7985
rect -1250 7965 -1230 7985
rect -1210 7965 -1190 7985
rect -1170 7965 -1150 7985
rect -1130 7965 -1110 7985
rect -1090 7965 -1070 7985
rect -1050 7965 -1030 7985
rect -1010 7965 -990 7985
rect -970 7965 -950 7985
rect -930 7965 -910 7985
rect -890 7965 -870 7985
rect -850 7965 -830 7985
rect -810 7965 -790 7985
rect -770 7965 -750 7985
rect -730 7965 -710 7985
rect -690 7965 -670 7985
rect -650 7965 -630 7985
rect -610 7965 -590 7985
rect -570 7965 -550 7985
rect -530 7965 -510 7985
rect -490 7965 -470 7985
rect -450 7965 -430 7985
rect -410 7965 -390 7985
rect -370 7965 -350 7985
rect -330 7965 -310 7985
rect -290 7965 -270 7985
rect -250 7965 -230 7985
rect -210 7965 -190 7985
rect -170 7965 -150 7985
rect -130 7965 -110 7985
rect -90 7965 -70 7985
rect -50 7965 -30 7985
rect -10 7965 10 7985
rect 30 7965 50 7985
rect 70 7965 90 7985
rect 110 7965 130 7985
rect 150 7965 170 7985
rect 190 7965 210 7985
rect 230 7965 250 7985
rect 270 7965 290 7985
rect 310 7965 330 7985
rect 350 7965 370 7985
rect 390 7965 410 7985
rect 430 7965 450 7985
rect 470 7965 490 7985
rect 510 7965 525 7985
rect -1975 7950 525 7965
rect -1975 7903 525 7918
rect -1975 7883 -1950 7903
rect -1930 7883 -1910 7903
rect -1890 7883 -1870 7903
rect -1850 7883 -1830 7903
rect -1810 7883 -1790 7903
rect -1770 7883 -1750 7903
rect -1730 7883 -1710 7903
rect -1690 7883 -1670 7903
rect -1650 7883 -1630 7903
rect -1610 7883 -1590 7903
rect -1570 7883 -1550 7903
rect -1530 7883 -1510 7903
rect -1490 7883 -1470 7903
rect -1450 7883 -1430 7903
rect -1410 7883 -1390 7903
rect -1370 7883 -1350 7903
rect -1330 7883 -1310 7903
rect -1290 7883 -1270 7903
rect -1250 7883 -1230 7903
rect -1210 7883 -1190 7903
rect -1170 7883 -1150 7903
rect -1130 7883 -1110 7903
rect -1090 7883 -1070 7903
rect -1050 7883 -1030 7903
rect -1010 7883 -990 7903
rect -970 7883 -950 7903
rect -930 7883 -910 7903
rect -890 7883 -870 7903
rect -850 7883 -830 7903
rect -810 7883 -790 7903
rect -770 7883 -750 7903
rect -730 7883 -710 7903
rect -690 7883 -670 7903
rect -650 7883 -630 7903
rect -610 7883 -590 7903
rect -570 7883 -550 7903
rect -530 7883 -510 7903
rect -490 7883 -470 7903
rect -450 7883 -430 7903
rect -410 7883 -390 7903
rect -370 7883 -350 7903
rect -330 7883 -310 7903
rect -290 7883 -270 7903
rect -250 7883 -230 7903
rect -210 7883 -190 7903
rect -170 7883 -150 7903
rect -130 7883 -110 7903
rect -90 7883 -70 7903
rect -50 7883 -30 7903
rect -10 7883 10 7903
rect 30 7883 50 7903
rect 70 7883 90 7903
rect 110 7883 130 7903
rect 150 7883 170 7903
rect 190 7883 210 7903
rect 230 7883 250 7903
rect 270 7883 290 7903
rect 310 7883 330 7903
rect 350 7883 370 7903
rect 390 7883 410 7903
rect 430 7883 450 7903
rect 470 7883 490 7903
rect 510 7883 525 7903
rect -1975 7868 525 7883
rect -1975 7821 525 7836
rect -1975 7801 -1950 7821
rect -1930 7801 -1910 7821
rect -1890 7801 -1870 7821
rect -1850 7801 -1830 7821
rect -1810 7801 -1790 7821
rect -1770 7801 -1750 7821
rect -1730 7801 -1710 7821
rect -1690 7801 -1670 7821
rect -1650 7801 -1630 7821
rect -1610 7801 -1590 7821
rect -1570 7801 -1550 7821
rect -1530 7801 -1510 7821
rect -1490 7801 -1470 7821
rect -1450 7801 -1430 7821
rect -1410 7801 -1390 7821
rect -1370 7801 -1350 7821
rect -1330 7801 -1310 7821
rect -1290 7801 -1270 7821
rect -1250 7801 -1230 7821
rect -1210 7801 -1190 7821
rect -1170 7801 -1150 7821
rect -1130 7801 -1110 7821
rect -1090 7801 -1070 7821
rect -1050 7801 -1030 7821
rect -1010 7801 -990 7821
rect -970 7801 -950 7821
rect -930 7801 -910 7821
rect -890 7801 -870 7821
rect -850 7801 -830 7821
rect -810 7801 -790 7821
rect -770 7801 -750 7821
rect -730 7801 -710 7821
rect -690 7801 -670 7821
rect -650 7801 -630 7821
rect -610 7801 -590 7821
rect -570 7801 -550 7821
rect -530 7801 -510 7821
rect -490 7801 -470 7821
rect -450 7801 -430 7821
rect -410 7801 -390 7821
rect -370 7801 -350 7821
rect -330 7801 -310 7821
rect -290 7801 -270 7821
rect -250 7801 -230 7821
rect -210 7801 -190 7821
rect -170 7801 -150 7821
rect -130 7801 -110 7821
rect -90 7801 -70 7821
rect -50 7801 -30 7821
rect -10 7801 10 7821
rect 30 7801 50 7821
rect 70 7801 90 7821
rect 110 7801 130 7821
rect 150 7801 170 7821
rect 190 7801 210 7821
rect 230 7801 250 7821
rect 270 7801 290 7821
rect 310 7801 330 7821
rect 350 7801 370 7821
rect 390 7801 410 7821
rect 430 7801 450 7821
rect 470 7801 490 7821
rect 510 7801 525 7821
rect -1975 7786 525 7801
rect -1975 7739 525 7754
rect -1975 7719 -1950 7739
rect -1930 7719 -1910 7739
rect -1890 7719 -1870 7739
rect -1850 7719 -1830 7739
rect -1810 7719 -1790 7739
rect -1770 7719 -1750 7739
rect -1730 7719 -1710 7739
rect -1690 7719 -1670 7739
rect -1650 7719 -1630 7739
rect -1610 7719 -1590 7739
rect -1570 7719 -1550 7739
rect -1530 7719 -1510 7739
rect -1490 7719 -1470 7739
rect -1450 7719 -1430 7739
rect -1410 7719 -1390 7739
rect -1370 7719 -1350 7739
rect -1330 7719 -1310 7739
rect -1290 7719 -1270 7739
rect -1250 7719 -1230 7739
rect -1210 7719 -1190 7739
rect -1170 7719 -1150 7739
rect -1130 7719 -1110 7739
rect -1090 7719 -1070 7739
rect -1050 7719 -1030 7739
rect -1010 7719 -990 7739
rect -970 7719 -950 7739
rect -930 7719 -910 7739
rect -890 7719 -870 7739
rect -850 7719 -830 7739
rect -810 7719 -790 7739
rect -770 7719 -750 7739
rect -730 7719 -710 7739
rect -690 7719 -670 7739
rect -650 7719 -630 7739
rect -610 7719 -590 7739
rect -570 7719 -550 7739
rect -530 7719 -510 7739
rect -490 7719 -470 7739
rect -450 7719 -430 7739
rect -410 7719 -390 7739
rect -370 7719 -350 7739
rect -330 7719 -310 7739
rect -290 7719 -270 7739
rect -250 7719 -230 7739
rect -210 7719 -190 7739
rect -170 7719 -150 7739
rect -130 7719 -110 7739
rect -90 7719 -70 7739
rect -50 7719 -30 7739
rect -10 7719 10 7739
rect 30 7719 50 7739
rect 70 7719 90 7739
rect 110 7719 130 7739
rect 150 7719 170 7739
rect 190 7719 210 7739
rect 230 7719 250 7739
rect 270 7719 290 7739
rect 310 7719 330 7739
rect 350 7719 370 7739
rect 390 7719 410 7739
rect 430 7719 450 7739
rect 470 7719 490 7739
rect 510 7719 525 7739
rect -1975 7704 525 7719
rect -1975 7657 525 7672
rect -1975 7637 -1950 7657
rect -1930 7637 -1910 7657
rect -1890 7637 -1870 7657
rect -1850 7637 -1830 7657
rect -1810 7637 -1790 7657
rect -1770 7637 -1750 7657
rect -1730 7637 -1710 7657
rect -1690 7637 -1670 7657
rect -1650 7637 -1630 7657
rect -1610 7637 -1590 7657
rect -1570 7637 -1550 7657
rect -1530 7637 -1510 7657
rect -1490 7637 -1470 7657
rect -1450 7637 -1430 7657
rect -1410 7637 -1390 7657
rect -1370 7637 -1350 7657
rect -1330 7637 -1310 7657
rect -1290 7637 -1270 7657
rect -1250 7637 -1230 7657
rect -1210 7637 -1190 7657
rect -1170 7637 -1150 7657
rect -1130 7637 -1110 7657
rect -1090 7637 -1070 7657
rect -1050 7637 -1030 7657
rect -1010 7637 -990 7657
rect -970 7637 -950 7657
rect -930 7637 -910 7657
rect -890 7637 -870 7657
rect -850 7637 -830 7657
rect -810 7637 -790 7657
rect -770 7637 -750 7657
rect -730 7637 -710 7657
rect -690 7637 -670 7657
rect -650 7637 -630 7657
rect -610 7637 -590 7657
rect -570 7637 -550 7657
rect -530 7637 -510 7657
rect -490 7637 -470 7657
rect -450 7637 -430 7657
rect -410 7637 -390 7657
rect -370 7637 -350 7657
rect -330 7637 -310 7657
rect -290 7637 -270 7657
rect -250 7637 -230 7657
rect -210 7637 -190 7657
rect -170 7637 -150 7657
rect -130 7637 -110 7657
rect -90 7637 -70 7657
rect -50 7637 -30 7657
rect -10 7637 10 7657
rect 30 7637 50 7657
rect 70 7637 90 7657
rect 110 7637 130 7657
rect 150 7637 170 7657
rect 190 7637 210 7657
rect 230 7637 250 7657
rect 270 7637 290 7657
rect 310 7637 330 7657
rect 350 7637 370 7657
rect 390 7637 410 7657
rect 430 7637 450 7657
rect 470 7637 490 7657
rect 510 7637 525 7657
rect -1975 7622 525 7637
rect -1975 7575 525 7590
rect -1975 7555 -1950 7575
rect -1930 7555 -1910 7575
rect -1890 7555 -1870 7575
rect -1850 7555 -1830 7575
rect -1810 7555 -1790 7575
rect -1770 7555 -1750 7575
rect -1730 7555 -1710 7575
rect -1690 7555 -1670 7575
rect -1650 7555 -1630 7575
rect -1610 7555 -1590 7575
rect -1570 7555 -1550 7575
rect -1530 7555 -1510 7575
rect -1490 7555 -1470 7575
rect -1450 7555 -1430 7575
rect -1410 7555 -1390 7575
rect -1370 7555 -1350 7575
rect -1330 7555 -1310 7575
rect -1290 7555 -1270 7575
rect -1250 7555 -1230 7575
rect -1210 7555 -1190 7575
rect -1170 7555 -1150 7575
rect -1130 7555 -1110 7575
rect -1090 7555 -1070 7575
rect -1050 7555 -1030 7575
rect -1010 7555 -990 7575
rect -970 7555 -950 7575
rect -930 7555 -910 7575
rect -890 7555 -870 7575
rect -850 7555 -830 7575
rect -810 7555 -790 7575
rect -770 7555 -750 7575
rect -730 7555 -710 7575
rect -690 7555 -670 7575
rect -650 7555 -630 7575
rect -610 7555 -590 7575
rect -570 7555 -550 7575
rect -530 7555 -510 7575
rect -490 7555 -470 7575
rect -450 7555 -430 7575
rect -410 7555 -390 7575
rect -370 7555 -350 7575
rect -330 7555 -310 7575
rect -290 7555 -270 7575
rect -250 7555 -230 7575
rect -210 7555 -190 7575
rect -170 7555 -150 7575
rect -130 7555 -110 7575
rect -90 7555 -70 7575
rect -50 7555 -30 7575
rect -10 7555 10 7575
rect 30 7555 50 7575
rect 70 7555 90 7575
rect 110 7555 130 7575
rect 150 7555 170 7575
rect 190 7555 210 7575
rect 230 7555 250 7575
rect 270 7555 290 7575
rect 310 7555 330 7575
rect 350 7555 370 7575
rect 390 7555 410 7575
rect 430 7555 450 7575
rect 470 7555 490 7575
rect 510 7555 525 7575
rect -1975 7540 525 7555
rect -1975 7493 525 7508
rect -1975 7473 -1950 7493
rect -1930 7473 -1910 7493
rect -1890 7473 -1870 7493
rect -1850 7473 -1830 7493
rect -1810 7473 -1790 7493
rect -1770 7473 -1750 7493
rect -1730 7473 -1710 7493
rect -1690 7473 -1670 7493
rect -1650 7473 -1630 7493
rect -1610 7473 -1590 7493
rect -1570 7473 -1550 7493
rect -1530 7473 -1510 7493
rect -1490 7473 -1470 7493
rect -1450 7473 -1430 7493
rect -1410 7473 -1390 7493
rect -1370 7473 -1350 7493
rect -1330 7473 -1310 7493
rect -1290 7473 -1270 7493
rect -1250 7473 -1230 7493
rect -1210 7473 -1190 7493
rect -1170 7473 -1150 7493
rect -1130 7473 -1110 7493
rect -1090 7473 -1070 7493
rect -1050 7473 -1030 7493
rect -1010 7473 -990 7493
rect -970 7473 -950 7493
rect -930 7473 -910 7493
rect -890 7473 -870 7493
rect -850 7473 -830 7493
rect -810 7473 -790 7493
rect -770 7473 -750 7493
rect -730 7473 -710 7493
rect -690 7473 -670 7493
rect -650 7473 -630 7493
rect -610 7473 -590 7493
rect -570 7473 -550 7493
rect -530 7473 -510 7493
rect -490 7473 -470 7493
rect -450 7473 -430 7493
rect -410 7473 -390 7493
rect -370 7473 -350 7493
rect -330 7473 -310 7493
rect -290 7473 -270 7493
rect -250 7473 -230 7493
rect -210 7473 -190 7493
rect -170 7473 -150 7493
rect -130 7473 -110 7493
rect -90 7473 -70 7493
rect -50 7473 -30 7493
rect -10 7473 10 7493
rect 30 7473 50 7493
rect 70 7473 90 7493
rect 110 7473 130 7493
rect 150 7473 170 7493
rect 190 7473 210 7493
rect 230 7473 250 7493
rect 270 7473 290 7493
rect 310 7473 330 7493
rect 350 7473 370 7493
rect 390 7473 410 7493
rect 430 7473 450 7493
rect 470 7473 490 7493
rect 510 7473 525 7493
rect -1975 7458 525 7473
rect -1975 7411 525 7426
rect -1975 7391 -1950 7411
rect -1930 7391 -1910 7411
rect -1890 7391 -1870 7411
rect -1850 7391 -1830 7411
rect -1810 7391 -1790 7411
rect -1770 7391 -1750 7411
rect -1730 7391 -1710 7411
rect -1690 7391 -1670 7411
rect -1650 7391 -1630 7411
rect -1610 7391 -1590 7411
rect -1570 7391 -1550 7411
rect -1530 7391 -1510 7411
rect -1490 7391 -1470 7411
rect -1450 7391 -1430 7411
rect -1410 7391 -1390 7411
rect -1370 7391 -1350 7411
rect -1330 7391 -1310 7411
rect -1290 7391 -1270 7411
rect -1250 7391 -1230 7411
rect -1210 7391 -1190 7411
rect -1170 7391 -1150 7411
rect -1130 7391 -1110 7411
rect -1090 7391 -1070 7411
rect -1050 7391 -1030 7411
rect -1010 7391 -990 7411
rect -970 7391 -950 7411
rect -930 7391 -910 7411
rect -890 7391 -870 7411
rect -850 7391 -830 7411
rect -810 7391 -790 7411
rect -770 7391 -750 7411
rect -730 7391 -710 7411
rect -690 7391 -670 7411
rect -650 7391 -630 7411
rect -610 7391 -590 7411
rect -570 7391 -550 7411
rect -530 7391 -510 7411
rect -490 7391 -470 7411
rect -450 7391 -430 7411
rect -410 7391 -390 7411
rect -370 7391 -350 7411
rect -330 7391 -310 7411
rect -290 7391 -270 7411
rect -250 7391 -230 7411
rect -210 7391 -190 7411
rect -170 7391 -150 7411
rect -130 7391 -110 7411
rect -90 7391 -70 7411
rect -50 7391 -30 7411
rect -10 7391 10 7411
rect 30 7391 50 7411
rect 70 7391 90 7411
rect 110 7391 130 7411
rect 150 7391 170 7411
rect 190 7391 210 7411
rect 230 7391 250 7411
rect 270 7391 290 7411
rect 310 7391 330 7411
rect 350 7391 370 7411
rect 390 7391 410 7411
rect 430 7391 450 7411
rect 470 7391 490 7411
rect 510 7391 525 7411
rect -1975 7376 525 7391
rect -1975 7329 525 7344
rect -1975 7309 -1950 7329
rect -1930 7309 -1910 7329
rect -1890 7309 -1870 7329
rect -1850 7309 -1830 7329
rect -1810 7309 -1790 7329
rect -1770 7309 -1750 7329
rect -1730 7309 -1710 7329
rect -1690 7309 -1670 7329
rect -1650 7309 -1630 7329
rect -1610 7309 -1590 7329
rect -1570 7309 -1550 7329
rect -1530 7309 -1510 7329
rect -1490 7309 -1470 7329
rect -1450 7309 -1430 7329
rect -1410 7309 -1390 7329
rect -1370 7309 -1350 7329
rect -1330 7309 -1310 7329
rect -1290 7309 -1270 7329
rect -1250 7309 -1230 7329
rect -1210 7309 -1190 7329
rect -1170 7309 -1150 7329
rect -1130 7309 -1110 7329
rect -1090 7309 -1070 7329
rect -1050 7309 -1030 7329
rect -1010 7309 -990 7329
rect -970 7309 -950 7329
rect -930 7309 -910 7329
rect -890 7309 -870 7329
rect -850 7309 -830 7329
rect -810 7309 -790 7329
rect -770 7309 -750 7329
rect -730 7309 -710 7329
rect -690 7309 -670 7329
rect -650 7309 -630 7329
rect -610 7309 -590 7329
rect -570 7309 -550 7329
rect -530 7309 -510 7329
rect -490 7309 -470 7329
rect -450 7309 -430 7329
rect -410 7309 -390 7329
rect -370 7309 -350 7329
rect -330 7309 -310 7329
rect -290 7309 -270 7329
rect -250 7309 -230 7329
rect -210 7309 -190 7329
rect -170 7309 -150 7329
rect -130 7309 -110 7329
rect -90 7309 -70 7329
rect -50 7309 -30 7329
rect -10 7309 10 7329
rect 30 7309 50 7329
rect 70 7309 90 7329
rect 110 7309 130 7329
rect 150 7309 170 7329
rect 190 7309 210 7329
rect 230 7309 250 7329
rect 270 7309 290 7329
rect 310 7309 330 7329
rect 350 7309 370 7329
rect 390 7309 410 7329
rect 430 7309 450 7329
rect 470 7309 490 7329
rect 510 7309 525 7329
rect -1975 7294 525 7309
rect -1975 7247 525 7262
rect -1975 7227 -1950 7247
rect -1930 7227 -1910 7247
rect -1890 7227 -1870 7247
rect -1850 7227 -1830 7247
rect -1810 7227 -1790 7247
rect -1770 7227 -1750 7247
rect -1730 7227 -1710 7247
rect -1690 7227 -1670 7247
rect -1650 7227 -1630 7247
rect -1610 7227 -1590 7247
rect -1570 7227 -1550 7247
rect -1530 7227 -1510 7247
rect -1490 7227 -1470 7247
rect -1450 7227 -1430 7247
rect -1410 7227 -1390 7247
rect -1370 7227 -1350 7247
rect -1330 7227 -1310 7247
rect -1290 7227 -1270 7247
rect -1250 7227 -1230 7247
rect -1210 7227 -1190 7247
rect -1170 7227 -1150 7247
rect -1130 7227 -1110 7247
rect -1090 7227 -1070 7247
rect -1050 7227 -1030 7247
rect -1010 7227 -990 7247
rect -970 7227 -950 7247
rect -930 7227 -910 7247
rect -890 7227 -870 7247
rect -850 7227 -830 7247
rect -810 7227 -790 7247
rect -770 7227 -750 7247
rect -730 7227 -710 7247
rect -690 7227 -670 7247
rect -650 7227 -630 7247
rect -610 7227 -590 7247
rect -570 7227 -550 7247
rect -530 7227 -510 7247
rect -490 7227 -470 7247
rect -450 7227 -430 7247
rect -410 7227 -390 7247
rect -370 7227 -350 7247
rect -330 7227 -310 7247
rect -290 7227 -270 7247
rect -250 7227 -230 7247
rect -210 7227 -190 7247
rect -170 7227 -150 7247
rect -130 7227 -110 7247
rect -90 7227 -70 7247
rect -50 7227 -30 7247
rect -10 7227 10 7247
rect 30 7227 50 7247
rect 70 7227 90 7247
rect 110 7227 130 7247
rect 150 7227 170 7247
rect 190 7227 210 7247
rect 230 7227 250 7247
rect 270 7227 290 7247
rect 310 7227 330 7247
rect 350 7227 370 7247
rect 390 7227 410 7247
rect 430 7227 450 7247
rect 470 7227 490 7247
rect 510 7227 525 7247
rect -1975 7212 525 7227
rect -1975 7165 525 7180
rect -1975 7145 -1950 7165
rect -1930 7145 -1910 7165
rect -1890 7145 -1870 7165
rect -1850 7145 -1830 7165
rect -1810 7145 -1790 7165
rect -1770 7145 -1750 7165
rect -1730 7145 -1710 7165
rect -1690 7145 -1670 7165
rect -1650 7145 -1630 7165
rect -1610 7145 -1590 7165
rect -1570 7145 -1550 7165
rect -1530 7145 -1510 7165
rect -1490 7145 -1470 7165
rect -1450 7145 -1430 7165
rect -1410 7145 -1390 7165
rect -1370 7145 -1350 7165
rect -1330 7145 -1310 7165
rect -1290 7145 -1270 7165
rect -1250 7145 -1230 7165
rect -1210 7145 -1190 7165
rect -1170 7145 -1150 7165
rect -1130 7145 -1110 7165
rect -1090 7145 -1070 7165
rect -1050 7145 -1030 7165
rect -1010 7145 -990 7165
rect -970 7145 -950 7165
rect -930 7145 -910 7165
rect -890 7145 -870 7165
rect -850 7145 -830 7165
rect -810 7145 -790 7165
rect -770 7145 -750 7165
rect -730 7145 -710 7165
rect -690 7145 -670 7165
rect -650 7145 -630 7165
rect -610 7145 -590 7165
rect -570 7145 -550 7165
rect -530 7145 -510 7165
rect -490 7145 -470 7165
rect -450 7145 -430 7165
rect -410 7145 -390 7165
rect -370 7145 -350 7165
rect -330 7145 -310 7165
rect -290 7145 -270 7165
rect -250 7145 -230 7165
rect -210 7145 -190 7165
rect -170 7145 -150 7165
rect -130 7145 -110 7165
rect -90 7145 -70 7165
rect -50 7145 -30 7165
rect -10 7145 10 7165
rect 30 7145 50 7165
rect 70 7145 90 7165
rect 110 7145 130 7165
rect 150 7145 170 7165
rect 190 7145 210 7165
rect 230 7145 250 7165
rect 270 7145 290 7165
rect 310 7145 330 7165
rect 350 7145 370 7165
rect 390 7145 410 7165
rect 430 7145 450 7165
rect 470 7145 490 7165
rect 510 7145 525 7165
rect -1975 7130 525 7145
rect -1975 7083 525 7098
rect -1975 7063 -1950 7083
rect -1930 7063 -1910 7083
rect -1890 7063 -1870 7083
rect -1850 7063 -1830 7083
rect -1810 7063 -1790 7083
rect -1770 7063 -1750 7083
rect -1730 7063 -1710 7083
rect -1690 7063 -1670 7083
rect -1650 7063 -1630 7083
rect -1610 7063 -1590 7083
rect -1570 7063 -1550 7083
rect -1530 7063 -1510 7083
rect -1490 7063 -1470 7083
rect -1450 7063 -1430 7083
rect -1410 7063 -1390 7083
rect -1370 7063 -1350 7083
rect -1330 7063 -1310 7083
rect -1290 7063 -1270 7083
rect -1250 7063 -1230 7083
rect -1210 7063 -1190 7083
rect -1170 7063 -1150 7083
rect -1130 7063 -1110 7083
rect -1090 7063 -1070 7083
rect -1050 7063 -1030 7083
rect -1010 7063 -990 7083
rect -970 7063 -950 7083
rect -930 7063 -910 7083
rect -890 7063 -870 7083
rect -850 7063 -830 7083
rect -810 7063 -790 7083
rect -770 7063 -750 7083
rect -730 7063 -710 7083
rect -690 7063 -670 7083
rect -650 7063 -630 7083
rect -610 7063 -590 7083
rect -570 7063 -550 7083
rect -530 7063 -510 7083
rect -490 7063 -470 7083
rect -450 7063 -430 7083
rect -410 7063 -390 7083
rect -370 7063 -350 7083
rect -330 7063 -310 7083
rect -290 7063 -270 7083
rect -250 7063 -230 7083
rect -210 7063 -190 7083
rect -170 7063 -150 7083
rect -130 7063 -110 7083
rect -90 7063 -70 7083
rect -50 7063 -30 7083
rect -10 7063 10 7083
rect 30 7063 50 7083
rect 70 7063 90 7083
rect 110 7063 130 7083
rect 150 7063 170 7083
rect 190 7063 210 7083
rect 230 7063 250 7083
rect 270 7063 290 7083
rect 310 7063 330 7083
rect 350 7063 370 7083
rect 390 7063 410 7083
rect 430 7063 450 7083
rect 470 7063 490 7083
rect 510 7063 525 7083
rect -1975 7048 525 7063
rect -1975 7001 525 7016
rect -1975 6981 -1950 7001
rect -1930 6981 -1910 7001
rect -1890 6981 -1870 7001
rect -1850 6981 -1830 7001
rect -1810 6981 -1790 7001
rect -1770 6981 -1750 7001
rect -1730 6981 -1710 7001
rect -1690 6981 -1670 7001
rect -1650 6981 -1630 7001
rect -1610 6981 -1590 7001
rect -1570 6981 -1550 7001
rect -1530 6981 -1510 7001
rect -1490 6981 -1470 7001
rect -1450 6981 -1430 7001
rect -1410 6981 -1390 7001
rect -1370 6981 -1350 7001
rect -1330 6981 -1310 7001
rect -1290 6981 -1270 7001
rect -1250 6981 -1230 7001
rect -1210 6981 -1190 7001
rect -1170 6981 -1150 7001
rect -1130 6981 -1110 7001
rect -1090 6981 -1070 7001
rect -1050 6981 -1030 7001
rect -1010 6981 -990 7001
rect -970 6981 -950 7001
rect -930 6981 -910 7001
rect -890 6981 -870 7001
rect -850 6981 -830 7001
rect -810 6981 -790 7001
rect -770 6981 -750 7001
rect -730 6981 -710 7001
rect -690 6981 -670 7001
rect -650 6981 -630 7001
rect -610 6981 -590 7001
rect -570 6981 -550 7001
rect -530 6981 -510 7001
rect -490 6981 -470 7001
rect -450 6981 -430 7001
rect -410 6981 -390 7001
rect -370 6981 -350 7001
rect -330 6981 -310 7001
rect -290 6981 -270 7001
rect -250 6981 -230 7001
rect -210 6981 -190 7001
rect -170 6981 -150 7001
rect -130 6981 -110 7001
rect -90 6981 -70 7001
rect -50 6981 -30 7001
rect -10 6981 10 7001
rect 30 6981 50 7001
rect 70 6981 90 7001
rect 110 6981 130 7001
rect 150 6981 170 7001
rect 190 6981 210 7001
rect 230 6981 250 7001
rect 270 6981 290 7001
rect 310 6981 330 7001
rect 350 6981 370 7001
rect 390 6981 410 7001
rect 430 6981 450 7001
rect 470 6981 490 7001
rect 510 6981 525 7001
rect -1975 6966 525 6981
rect -1975 6919 525 6934
rect -1975 6899 -1950 6919
rect -1930 6899 -1910 6919
rect -1890 6899 -1870 6919
rect -1850 6899 -1830 6919
rect -1810 6899 -1790 6919
rect -1770 6899 -1750 6919
rect -1730 6899 -1710 6919
rect -1690 6899 -1670 6919
rect -1650 6899 -1630 6919
rect -1610 6899 -1590 6919
rect -1570 6899 -1550 6919
rect -1530 6899 -1510 6919
rect -1490 6899 -1470 6919
rect -1450 6899 -1430 6919
rect -1410 6899 -1390 6919
rect -1370 6899 -1350 6919
rect -1330 6899 -1310 6919
rect -1290 6899 -1270 6919
rect -1250 6899 -1230 6919
rect -1210 6899 -1190 6919
rect -1170 6899 -1150 6919
rect -1130 6899 -1110 6919
rect -1090 6899 -1070 6919
rect -1050 6899 -1030 6919
rect -1010 6899 -990 6919
rect -970 6899 -950 6919
rect -930 6899 -910 6919
rect -890 6899 -870 6919
rect -850 6899 -830 6919
rect -810 6899 -790 6919
rect -770 6899 -750 6919
rect -730 6899 -710 6919
rect -690 6899 -670 6919
rect -650 6899 -630 6919
rect -610 6899 -590 6919
rect -570 6899 -550 6919
rect -530 6899 -510 6919
rect -490 6899 -470 6919
rect -450 6899 -430 6919
rect -410 6899 -390 6919
rect -370 6899 -350 6919
rect -330 6899 -310 6919
rect -290 6899 -270 6919
rect -250 6899 -230 6919
rect -210 6899 -190 6919
rect -170 6899 -150 6919
rect -130 6899 -110 6919
rect -90 6899 -70 6919
rect -50 6899 -30 6919
rect -10 6899 10 6919
rect 30 6899 50 6919
rect 70 6899 90 6919
rect 110 6899 130 6919
rect 150 6899 170 6919
rect 190 6899 210 6919
rect 230 6899 250 6919
rect 270 6899 290 6919
rect 310 6899 330 6919
rect 350 6899 370 6919
rect 390 6899 410 6919
rect 430 6899 450 6919
rect 470 6899 490 6919
rect 510 6899 525 6919
rect -1975 6884 525 6899
rect -1975 6837 525 6852
rect -1975 6817 -1950 6837
rect -1930 6817 -1910 6837
rect -1890 6817 -1870 6837
rect -1850 6817 -1830 6837
rect -1810 6817 -1790 6837
rect -1770 6817 -1750 6837
rect -1730 6817 -1710 6837
rect -1690 6817 -1670 6837
rect -1650 6817 -1630 6837
rect -1610 6817 -1590 6837
rect -1570 6817 -1550 6837
rect -1530 6817 -1510 6837
rect -1490 6817 -1470 6837
rect -1450 6817 -1430 6837
rect -1410 6817 -1390 6837
rect -1370 6817 -1350 6837
rect -1330 6817 -1310 6837
rect -1290 6817 -1270 6837
rect -1250 6817 -1230 6837
rect -1210 6817 -1190 6837
rect -1170 6817 -1150 6837
rect -1130 6817 -1110 6837
rect -1090 6817 -1070 6837
rect -1050 6817 -1030 6837
rect -1010 6817 -990 6837
rect -970 6817 -950 6837
rect -930 6817 -910 6837
rect -890 6817 -870 6837
rect -850 6817 -830 6837
rect -810 6817 -790 6837
rect -770 6817 -750 6837
rect -730 6817 -710 6837
rect -690 6817 -670 6837
rect -650 6817 -630 6837
rect -610 6817 -590 6837
rect -570 6817 -550 6837
rect -530 6817 -510 6837
rect -490 6817 -470 6837
rect -450 6817 -430 6837
rect -410 6817 -390 6837
rect -370 6817 -350 6837
rect -330 6817 -310 6837
rect -290 6817 -270 6837
rect -250 6817 -230 6837
rect -210 6817 -190 6837
rect -170 6817 -150 6837
rect -130 6817 -110 6837
rect -90 6817 -70 6837
rect -50 6817 -30 6837
rect -10 6817 10 6837
rect 30 6817 50 6837
rect 70 6817 90 6837
rect 110 6817 130 6837
rect 150 6817 170 6837
rect 190 6817 210 6837
rect 230 6817 250 6837
rect 270 6817 290 6837
rect 310 6817 330 6837
rect 350 6817 370 6837
rect 390 6817 410 6837
rect 430 6817 450 6837
rect 470 6817 490 6837
rect 510 6817 525 6837
rect -1975 6802 525 6817
rect -1975 6755 525 6770
rect -1975 6735 -1950 6755
rect -1930 6735 -1910 6755
rect -1890 6735 -1870 6755
rect -1850 6735 -1830 6755
rect -1810 6735 -1790 6755
rect -1770 6735 -1750 6755
rect -1730 6735 -1710 6755
rect -1690 6735 -1670 6755
rect -1650 6735 -1630 6755
rect -1610 6735 -1590 6755
rect -1570 6735 -1550 6755
rect -1530 6735 -1510 6755
rect -1490 6735 -1470 6755
rect -1450 6735 -1430 6755
rect -1410 6735 -1390 6755
rect -1370 6735 -1350 6755
rect -1330 6735 -1310 6755
rect -1290 6735 -1270 6755
rect -1250 6735 -1230 6755
rect -1210 6735 -1190 6755
rect -1170 6735 -1150 6755
rect -1130 6735 -1110 6755
rect -1090 6735 -1070 6755
rect -1050 6735 -1030 6755
rect -1010 6735 -990 6755
rect -970 6735 -950 6755
rect -930 6735 -910 6755
rect -890 6735 -870 6755
rect -850 6735 -830 6755
rect -810 6735 -790 6755
rect -770 6735 -750 6755
rect -730 6735 -710 6755
rect -690 6735 -670 6755
rect -650 6735 -630 6755
rect -610 6735 -590 6755
rect -570 6735 -550 6755
rect -530 6735 -510 6755
rect -490 6735 -470 6755
rect -450 6735 -430 6755
rect -410 6735 -390 6755
rect -370 6735 -350 6755
rect -330 6735 -310 6755
rect -290 6735 -270 6755
rect -250 6735 -230 6755
rect -210 6735 -190 6755
rect -170 6735 -150 6755
rect -130 6735 -110 6755
rect -90 6735 -70 6755
rect -50 6735 -30 6755
rect -10 6735 10 6755
rect 30 6735 50 6755
rect 70 6735 90 6755
rect 110 6735 130 6755
rect 150 6735 170 6755
rect 190 6735 210 6755
rect 230 6735 250 6755
rect 270 6735 290 6755
rect 310 6735 330 6755
rect 350 6735 370 6755
rect 390 6735 410 6755
rect 430 6735 450 6755
rect 470 6735 490 6755
rect 510 6735 525 6755
rect -1975 6720 525 6735
rect -1975 6673 525 6688
rect -1975 6653 -1950 6673
rect -1930 6653 -1910 6673
rect -1890 6653 -1870 6673
rect -1850 6653 -1830 6673
rect -1810 6653 -1790 6673
rect -1770 6653 -1750 6673
rect -1730 6653 -1710 6673
rect -1690 6653 -1670 6673
rect -1650 6653 -1630 6673
rect -1610 6653 -1590 6673
rect -1570 6653 -1550 6673
rect -1530 6653 -1510 6673
rect -1490 6653 -1470 6673
rect -1450 6653 -1430 6673
rect -1410 6653 -1390 6673
rect -1370 6653 -1350 6673
rect -1330 6653 -1310 6673
rect -1290 6653 -1270 6673
rect -1250 6653 -1230 6673
rect -1210 6653 -1190 6673
rect -1170 6653 -1150 6673
rect -1130 6653 -1110 6673
rect -1090 6653 -1070 6673
rect -1050 6653 -1030 6673
rect -1010 6653 -990 6673
rect -970 6653 -950 6673
rect -930 6653 -910 6673
rect -890 6653 -870 6673
rect -850 6653 -830 6673
rect -810 6653 -790 6673
rect -770 6653 -750 6673
rect -730 6653 -710 6673
rect -690 6653 -670 6673
rect -650 6653 -630 6673
rect -610 6653 -590 6673
rect -570 6653 -550 6673
rect -530 6653 -510 6673
rect -490 6653 -470 6673
rect -450 6653 -430 6673
rect -410 6653 -390 6673
rect -370 6653 -350 6673
rect -330 6653 -310 6673
rect -290 6653 -270 6673
rect -250 6653 -230 6673
rect -210 6653 -190 6673
rect -170 6653 -150 6673
rect -130 6653 -110 6673
rect -90 6653 -70 6673
rect -50 6653 -30 6673
rect -10 6653 10 6673
rect 30 6653 50 6673
rect 70 6653 90 6673
rect 110 6653 130 6673
rect 150 6653 170 6673
rect 190 6653 210 6673
rect 230 6653 250 6673
rect 270 6653 290 6673
rect 310 6653 330 6673
rect 350 6653 370 6673
rect 390 6653 410 6673
rect 430 6653 450 6673
rect 470 6653 490 6673
rect 510 6653 525 6673
rect -1975 6638 525 6653
rect -1975 6591 525 6606
rect -1975 6571 -1950 6591
rect -1930 6571 -1910 6591
rect -1890 6571 -1870 6591
rect -1850 6571 -1830 6591
rect -1810 6571 -1790 6591
rect -1770 6571 -1750 6591
rect -1730 6571 -1710 6591
rect -1690 6571 -1670 6591
rect -1650 6571 -1630 6591
rect -1610 6571 -1590 6591
rect -1570 6571 -1550 6591
rect -1530 6571 -1510 6591
rect -1490 6571 -1470 6591
rect -1450 6571 -1430 6591
rect -1410 6571 -1390 6591
rect -1370 6571 -1350 6591
rect -1330 6571 -1310 6591
rect -1290 6571 -1270 6591
rect -1250 6571 -1230 6591
rect -1210 6571 -1190 6591
rect -1170 6571 -1150 6591
rect -1130 6571 -1110 6591
rect -1090 6571 -1070 6591
rect -1050 6571 -1030 6591
rect -1010 6571 -990 6591
rect -970 6571 -950 6591
rect -930 6571 -910 6591
rect -890 6571 -870 6591
rect -850 6571 -830 6591
rect -810 6571 -790 6591
rect -770 6571 -750 6591
rect -730 6571 -710 6591
rect -690 6571 -670 6591
rect -650 6571 -630 6591
rect -610 6571 -590 6591
rect -570 6571 -550 6591
rect -530 6571 -510 6591
rect -490 6571 -470 6591
rect -450 6571 -430 6591
rect -410 6571 -390 6591
rect -370 6571 -350 6591
rect -330 6571 -310 6591
rect -290 6571 -270 6591
rect -250 6571 -230 6591
rect -210 6571 -190 6591
rect -170 6571 -150 6591
rect -130 6571 -110 6591
rect -90 6571 -70 6591
rect -50 6571 -30 6591
rect -10 6571 10 6591
rect 30 6571 50 6591
rect 70 6571 90 6591
rect 110 6571 130 6591
rect 150 6571 170 6591
rect 190 6571 210 6591
rect 230 6571 250 6591
rect 270 6571 290 6591
rect 310 6571 330 6591
rect 350 6571 370 6591
rect 390 6571 410 6591
rect 430 6571 450 6591
rect 470 6571 490 6591
rect 510 6571 525 6591
rect -1975 6556 525 6571
rect -1975 6509 525 6524
rect -1975 6489 -1950 6509
rect -1930 6489 -1910 6509
rect -1890 6489 -1870 6509
rect -1850 6489 -1830 6509
rect -1810 6489 -1790 6509
rect -1770 6489 -1750 6509
rect -1730 6489 -1710 6509
rect -1690 6489 -1670 6509
rect -1650 6489 -1630 6509
rect -1610 6489 -1590 6509
rect -1570 6489 -1550 6509
rect -1530 6489 -1510 6509
rect -1490 6489 -1470 6509
rect -1450 6489 -1430 6509
rect -1410 6489 -1390 6509
rect -1370 6489 -1350 6509
rect -1330 6489 -1310 6509
rect -1290 6489 -1270 6509
rect -1250 6489 -1230 6509
rect -1210 6489 -1190 6509
rect -1170 6489 -1150 6509
rect -1130 6489 -1110 6509
rect -1090 6489 -1070 6509
rect -1050 6489 -1030 6509
rect -1010 6489 -990 6509
rect -970 6489 -950 6509
rect -930 6489 -910 6509
rect -890 6489 -870 6509
rect -850 6489 -830 6509
rect -810 6489 -790 6509
rect -770 6489 -750 6509
rect -730 6489 -710 6509
rect -690 6489 -670 6509
rect -650 6489 -630 6509
rect -610 6489 -590 6509
rect -570 6489 -550 6509
rect -530 6489 -510 6509
rect -490 6489 -470 6509
rect -450 6489 -430 6509
rect -410 6489 -390 6509
rect -370 6489 -350 6509
rect -330 6489 -310 6509
rect -290 6489 -270 6509
rect -250 6489 -230 6509
rect -210 6489 -190 6509
rect -170 6489 -150 6509
rect -130 6489 -110 6509
rect -90 6489 -70 6509
rect -50 6489 -30 6509
rect -10 6489 10 6509
rect 30 6489 50 6509
rect 70 6489 90 6509
rect 110 6489 130 6509
rect 150 6489 170 6509
rect 190 6489 210 6509
rect 230 6489 250 6509
rect 270 6489 290 6509
rect 310 6489 330 6509
rect 350 6489 370 6509
rect 390 6489 410 6509
rect 430 6489 450 6509
rect 470 6489 490 6509
rect 510 6489 525 6509
rect -1975 6474 525 6489
rect -1975 6427 525 6442
rect -1975 6407 -1950 6427
rect -1930 6407 -1910 6427
rect -1890 6407 -1870 6427
rect -1850 6407 -1830 6427
rect -1810 6407 -1790 6427
rect -1770 6407 -1750 6427
rect -1730 6407 -1710 6427
rect -1690 6407 -1670 6427
rect -1650 6407 -1630 6427
rect -1610 6407 -1590 6427
rect -1570 6407 -1550 6427
rect -1530 6407 -1510 6427
rect -1490 6407 -1470 6427
rect -1450 6407 -1430 6427
rect -1410 6407 -1390 6427
rect -1370 6407 -1350 6427
rect -1330 6407 -1310 6427
rect -1290 6407 -1270 6427
rect -1250 6407 -1230 6427
rect -1210 6407 -1190 6427
rect -1170 6407 -1150 6427
rect -1130 6407 -1110 6427
rect -1090 6407 -1070 6427
rect -1050 6407 -1030 6427
rect -1010 6407 -990 6427
rect -970 6407 -950 6427
rect -930 6407 -910 6427
rect -890 6407 -870 6427
rect -850 6407 -830 6427
rect -810 6407 -790 6427
rect -770 6407 -750 6427
rect -730 6407 -710 6427
rect -690 6407 -670 6427
rect -650 6407 -630 6427
rect -610 6407 -590 6427
rect -570 6407 -550 6427
rect -530 6407 -510 6427
rect -490 6407 -470 6427
rect -450 6407 -430 6427
rect -410 6407 -390 6427
rect -370 6407 -350 6427
rect -330 6407 -310 6427
rect -290 6407 -270 6427
rect -250 6407 -230 6427
rect -210 6407 -190 6427
rect -170 6407 -150 6427
rect -130 6407 -110 6427
rect -90 6407 -70 6427
rect -50 6407 -30 6427
rect -10 6407 10 6427
rect 30 6407 50 6427
rect 70 6407 90 6427
rect 110 6407 130 6427
rect 150 6407 170 6427
rect 190 6407 210 6427
rect 230 6407 250 6427
rect 270 6407 290 6427
rect 310 6407 330 6427
rect 350 6407 370 6427
rect 390 6407 410 6427
rect 430 6407 450 6427
rect 470 6407 490 6427
rect 510 6407 525 6427
rect -1975 6392 525 6407
rect -1975 6345 525 6360
rect -1975 6325 -1950 6345
rect -1930 6325 -1910 6345
rect -1890 6325 -1870 6345
rect -1850 6325 -1830 6345
rect -1810 6325 -1790 6345
rect -1770 6325 -1750 6345
rect -1730 6325 -1710 6345
rect -1690 6325 -1670 6345
rect -1650 6325 -1630 6345
rect -1610 6325 -1590 6345
rect -1570 6325 -1550 6345
rect -1530 6325 -1510 6345
rect -1490 6325 -1470 6345
rect -1450 6325 -1430 6345
rect -1410 6325 -1390 6345
rect -1370 6325 -1350 6345
rect -1330 6325 -1310 6345
rect -1290 6325 -1270 6345
rect -1250 6325 -1230 6345
rect -1210 6325 -1190 6345
rect -1170 6325 -1150 6345
rect -1130 6325 -1110 6345
rect -1090 6325 -1070 6345
rect -1050 6325 -1030 6345
rect -1010 6325 -990 6345
rect -970 6325 -950 6345
rect -930 6325 -910 6345
rect -890 6325 -870 6345
rect -850 6325 -830 6345
rect -810 6325 -790 6345
rect -770 6325 -750 6345
rect -730 6325 -710 6345
rect -690 6325 -670 6345
rect -650 6325 -630 6345
rect -610 6325 -590 6345
rect -570 6325 -550 6345
rect -530 6325 -510 6345
rect -490 6325 -470 6345
rect -450 6325 -430 6345
rect -410 6325 -390 6345
rect -370 6325 -350 6345
rect -330 6325 -310 6345
rect -290 6325 -270 6345
rect -250 6325 -230 6345
rect -210 6325 -190 6345
rect -170 6325 -150 6345
rect -130 6325 -110 6345
rect -90 6325 -70 6345
rect -50 6325 -30 6345
rect -10 6325 10 6345
rect 30 6325 50 6345
rect 70 6325 90 6345
rect 110 6325 130 6345
rect 150 6325 170 6345
rect 190 6325 210 6345
rect 230 6325 250 6345
rect 270 6325 290 6345
rect 310 6325 330 6345
rect 350 6325 370 6345
rect 390 6325 410 6345
rect 430 6325 450 6345
rect 470 6325 490 6345
rect 510 6325 525 6345
rect -1975 6315 525 6325
rect -5595 6045 -3095 6055
rect -5595 6025 -5580 6045
rect -5550 6025 -5530 6045
rect -5510 6025 -5490 6045
rect -5470 6025 -5450 6045
rect -5430 6025 -5410 6045
rect -5390 6025 -5370 6045
rect -5350 6025 -5330 6045
rect -5310 6025 -5290 6045
rect -5270 6025 -5250 6045
rect -5230 6025 -5210 6045
rect -5190 6025 -5170 6045
rect -5150 6025 -5130 6045
rect -5110 6025 -5090 6045
rect -5070 6025 -5050 6045
rect -5030 6025 -5010 6045
rect -4990 6025 -4970 6045
rect -4950 6025 -4930 6045
rect -4910 6025 -4890 6045
rect -4870 6025 -4850 6045
rect -4830 6025 -4810 6045
rect -4790 6025 -4770 6045
rect -4750 6025 -4730 6045
rect -4710 6025 -4690 6045
rect -4670 6025 -4650 6045
rect -4630 6025 -4610 6045
rect -4590 6025 -4570 6045
rect -4550 6025 -4530 6045
rect -4510 6025 -4490 6045
rect -4470 6025 -4450 6045
rect -4430 6025 -4410 6045
rect -4390 6025 -4370 6045
rect -4350 6025 -4330 6045
rect -4310 6025 -4290 6045
rect -4270 6025 -4250 6045
rect -4230 6025 -4210 6045
rect -4190 6025 -4170 6045
rect -4150 6025 -4130 6045
rect -4110 6025 -4090 6045
rect -4070 6025 -4050 6045
rect -4030 6025 -4010 6045
rect -3990 6025 -3970 6045
rect -3950 6025 -3930 6045
rect -3910 6025 -3890 6045
rect -3870 6025 -3850 6045
rect -3830 6025 -3810 6045
rect -3790 6025 -3770 6045
rect -3750 6025 -3730 6045
rect -3710 6025 -3690 6045
rect -3670 6025 -3650 6045
rect -3630 6025 -3610 6045
rect -3590 6025 -3570 6045
rect -3550 6025 -3530 6045
rect -3510 6025 -3490 6045
rect -3470 6025 -3450 6045
rect -3430 6025 -3410 6045
rect -3390 6025 -3370 6045
rect -3350 6025 -3330 6045
rect -3310 6025 -3290 6045
rect -3270 6025 -3250 6045
rect -3230 6025 -3210 6045
rect -3190 6025 -3170 6045
rect -3150 6025 -3130 6045
rect -3110 6025 -3095 6045
rect -5595 6010 -3095 6025
rect -2045 6045 455 6055
rect -2045 6025 -2030 6045
rect -2010 6025 -1990 6045
rect -1970 6025 -1950 6045
rect -1930 6025 -1910 6045
rect -1890 6025 -1870 6045
rect -1850 6025 -1830 6045
rect -1810 6025 -1790 6045
rect -1770 6025 -1750 6045
rect -1730 6025 -1710 6045
rect -1690 6025 -1670 6045
rect -1650 6025 -1630 6045
rect -1610 6025 -1590 6045
rect -1570 6025 -1550 6045
rect -1530 6025 -1510 6045
rect -1490 6025 -1470 6045
rect -1450 6025 -1430 6045
rect -1410 6025 -1390 6045
rect -1370 6025 -1350 6045
rect -1330 6025 -1310 6045
rect -1290 6025 -1270 6045
rect -1250 6025 -1230 6045
rect -1210 6025 -1190 6045
rect -1170 6025 -1150 6045
rect -1130 6025 -1110 6045
rect -1090 6025 -1070 6045
rect -1050 6025 -1030 6045
rect -1010 6025 -990 6045
rect -970 6025 -950 6045
rect -930 6025 -910 6045
rect -890 6025 -870 6045
rect -850 6025 -830 6045
rect -810 6025 -790 6045
rect -770 6025 -750 6045
rect -730 6025 -710 6045
rect -690 6025 -670 6045
rect -650 6025 -630 6045
rect -610 6025 -590 6045
rect -570 6025 -550 6045
rect -530 6025 -510 6045
rect -490 6025 -470 6045
rect -450 6025 -430 6045
rect -410 6025 -390 6045
rect -370 6025 -350 6045
rect -330 6025 -310 6045
rect -290 6025 -270 6045
rect -250 6025 -230 6045
rect -210 6025 -190 6045
rect -170 6025 -150 6045
rect -130 6025 -110 6045
rect -90 6025 -70 6045
rect -50 6025 -30 6045
rect -10 6025 10 6045
rect 30 6025 50 6045
rect 70 6025 90 6045
rect 110 6025 130 6045
rect 150 6025 170 6045
rect 190 6025 210 6045
rect 230 6025 250 6045
rect 270 6025 290 6045
rect 310 6025 330 6045
rect 350 6025 370 6045
rect 390 6025 410 6045
rect 440 6025 455 6045
rect -2045 6010 455 6025
rect -5595 5950 -3095 5965
rect -5595 5930 -5580 5950
rect -5550 5930 -5530 5950
rect -5510 5930 -5490 5950
rect -5470 5930 -5450 5950
rect -5430 5930 -5410 5950
rect -5390 5930 -5370 5950
rect -5350 5930 -5330 5950
rect -5310 5930 -5290 5950
rect -5270 5930 -5250 5950
rect -5230 5930 -5210 5950
rect -5190 5930 -5170 5950
rect -5150 5930 -5130 5950
rect -5110 5930 -5090 5950
rect -5070 5930 -5050 5950
rect -5030 5930 -5010 5950
rect -4990 5930 -4970 5950
rect -4950 5930 -4930 5950
rect -4910 5930 -4890 5950
rect -4870 5930 -4850 5950
rect -4830 5930 -4810 5950
rect -4790 5930 -4770 5950
rect -4750 5930 -4730 5950
rect -4710 5930 -4690 5950
rect -4670 5930 -4650 5950
rect -4630 5930 -4610 5950
rect -4590 5930 -4570 5950
rect -4550 5930 -4530 5950
rect -4510 5930 -4490 5950
rect -4470 5930 -4450 5950
rect -4430 5930 -4410 5950
rect -4390 5930 -4370 5950
rect -4350 5930 -4330 5950
rect -4310 5930 -4290 5950
rect -4270 5930 -4250 5950
rect -4230 5930 -4210 5950
rect -4190 5930 -4170 5950
rect -4150 5930 -4130 5950
rect -4110 5930 -4090 5950
rect -4070 5930 -4050 5950
rect -4030 5930 -4010 5950
rect -3990 5930 -3970 5950
rect -3950 5930 -3930 5950
rect -3910 5930 -3890 5950
rect -3870 5930 -3850 5950
rect -3830 5930 -3810 5950
rect -3790 5930 -3770 5950
rect -3750 5930 -3730 5950
rect -3710 5930 -3690 5950
rect -3670 5930 -3650 5950
rect -3630 5930 -3610 5950
rect -3590 5930 -3570 5950
rect -3550 5930 -3530 5950
rect -3510 5930 -3490 5950
rect -3470 5930 -3450 5950
rect -3430 5930 -3410 5950
rect -3390 5930 -3370 5950
rect -3350 5930 -3330 5950
rect -3310 5930 -3290 5950
rect -3270 5930 -3250 5950
rect -3230 5930 -3210 5950
rect -3190 5930 -3170 5950
rect -3150 5930 -3130 5950
rect -3110 5930 -3095 5950
rect -5595 5915 -3095 5930
rect -2045 5950 455 5965
rect -2045 5930 -2030 5950
rect -2010 5930 -1990 5950
rect -1970 5930 -1950 5950
rect -1930 5930 -1910 5950
rect -1890 5930 -1870 5950
rect -1850 5930 -1830 5950
rect -1810 5930 -1790 5950
rect -1770 5930 -1750 5950
rect -1730 5930 -1710 5950
rect -1690 5930 -1670 5950
rect -1650 5930 -1630 5950
rect -1610 5930 -1590 5950
rect -1570 5930 -1550 5950
rect -1530 5930 -1510 5950
rect -1490 5930 -1470 5950
rect -1450 5930 -1430 5950
rect -1410 5930 -1390 5950
rect -1370 5930 -1350 5950
rect -1330 5930 -1310 5950
rect -1290 5930 -1270 5950
rect -1250 5930 -1230 5950
rect -1210 5930 -1190 5950
rect -1170 5930 -1150 5950
rect -1130 5930 -1110 5950
rect -1090 5930 -1070 5950
rect -1050 5930 -1030 5950
rect -1010 5930 -990 5950
rect -970 5930 -950 5950
rect -930 5930 -910 5950
rect -890 5930 -870 5950
rect -850 5930 -830 5950
rect -810 5930 -790 5950
rect -770 5930 -750 5950
rect -730 5930 -710 5950
rect -690 5930 -670 5950
rect -650 5930 -630 5950
rect -610 5930 -590 5950
rect -570 5930 -550 5950
rect -530 5930 -510 5950
rect -490 5930 -470 5950
rect -450 5930 -430 5950
rect -410 5930 -390 5950
rect -370 5930 -350 5950
rect -330 5930 -310 5950
rect -290 5930 -270 5950
rect -250 5930 -230 5950
rect -210 5930 -190 5950
rect -170 5930 -150 5950
rect -130 5930 -110 5950
rect -90 5930 -70 5950
rect -50 5930 -30 5950
rect -10 5930 10 5950
rect 30 5930 50 5950
rect 70 5930 90 5950
rect 110 5930 130 5950
rect 150 5930 170 5950
rect 190 5930 210 5950
rect 230 5930 250 5950
rect 270 5930 290 5950
rect 310 5930 330 5950
rect 350 5930 370 5950
rect 390 5930 410 5950
rect 440 5930 455 5950
rect -2045 5915 455 5930
rect -5595 5855 -3095 5870
rect -5595 5835 -5580 5855
rect -5550 5835 -5530 5855
rect -5510 5835 -5490 5855
rect -5470 5835 -5450 5855
rect -5430 5835 -5410 5855
rect -5390 5835 -5370 5855
rect -5350 5835 -5330 5855
rect -5310 5835 -5290 5855
rect -5270 5835 -5250 5855
rect -5230 5835 -5210 5855
rect -5190 5835 -5170 5855
rect -5150 5835 -5130 5855
rect -5110 5835 -5090 5855
rect -5070 5835 -5050 5855
rect -5030 5835 -5010 5855
rect -4990 5835 -4970 5855
rect -4950 5835 -4930 5855
rect -4910 5835 -4890 5855
rect -4870 5835 -4850 5855
rect -4830 5835 -4810 5855
rect -4790 5835 -4770 5855
rect -4750 5835 -4730 5855
rect -4710 5835 -4690 5855
rect -4670 5835 -4650 5855
rect -4630 5835 -4610 5855
rect -4590 5835 -4570 5855
rect -4550 5835 -4530 5855
rect -4510 5835 -4490 5855
rect -4470 5835 -4450 5855
rect -4430 5835 -4410 5855
rect -4390 5835 -4370 5855
rect -4350 5835 -4330 5855
rect -4310 5835 -4290 5855
rect -4270 5835 -4250 5855
rect -4230 5835 -4210 5855
rect -4190 5835 -4170 5855
rect -4150 5835 -4130 5855
rect -4110 5835 -4090 5855
rect -4070 5835 -4050 5855
rect -4030 5835 -4010 5855
rect -3990 5835 -3970 5855
rect -3950 5835 -3930 5855
rect -3910 5835 -3890 5855
rect -3870 5835 -3850 5855
rect -3830 5835 -3810 5855
rect -3790 5835 -3770 5855
rect -3750 5835 -3730 5855
rect -3710 5835 -3690 5855
rect -3670 5835 -3650 5855
rect -3630 5835 -3610 5855
rect -3590 5835 -3570 5855
rect -3550 5835 -3530 5855
rect -3510 5835 -3490 5855
rect -3470 5835 -3450 5855
rect -3430 5835 -3410 5855
rect -3390 5835 -3370 5855
rect -3350 5835 -3330 5855
rect -3310 5835 -3290 5855
rect -3270 5835 -3250 5855
rect -3230 5835 -3210 5855
rect -3190 5835 -3170 5855
rect -3150 5835 -3130 5855
rect -3110 5835 -3095 5855
rect -5595 5820 -3095 5835
rect -2045 5855 455 5870
rect -2045 5835 -2030 5855
rect -2010 5835 -1990 5855
rect -1970 5835 -1950 5855
rect -1930 5835 -1910 5855
rect -1890 5835 -1870 5855
rect -1850 5835 -1830 5855
rect -1810 5835 -1790 5855
rect -1770 5835 -1750 5855
rect -1730 5835 -1710 5855
rect -1690 5835 -1670 5855
rect -1650 5835 -1630 5855
rect -1610 5835 -1590 5855
rect -1570 5835 -1550 5855
rect -1530 5835 -1510 5855
rect -1490 5835 -1470 5855
rect -1450 5835 -1430 5855
rect -1410 5835 -1390 5855
rect -1370 5835 -1350 5855
rect -1330 5835 -1310 5855
rect -1290 5835 -1270 5855
rect -1250 5835 -1230 5855
rect -1210 5835 -1190 5855
rect -1170 5835 -1150 5855
rect -1130 5835 -1110 5855
rect -1090 5835 -1070 5855
rect -1050 5835 -1030 5855
rect -1010 5835 -990 5855
rect -970 5835 -950 5855
rect -930 5835 -910 5855
rect -890 5835 -870 5855
rect -850 5835 -830 5855
rect -810 5835 -790 5855
rect -770 5835 -750 5855
rect -730 5835 -710 5855
rect -690 5835 -670 5855
rect -650 5835 -630 5855
rect -610 5835 -590 5855
rect -570 5835 -550 5855
rect -530 5835 -510 5855
rect -490 5835 -470 5855
rect -450 5835 -430 5855
rect -410 5835 -390 5855
rect -370 5835 -350 5855
rect -330 5835 -310 5855
rect -290 5835 -270 5855
rect -250 5835 -230 5855
rect -210 5835 -190 5855
rect -170 5835 -150 5855
rect -130 5835 -110 5855
rect -90 5835 -70 5855
rect -50 5835 -30 5855
rect -10 5835 10 5855
rect 30 5835 50 5855
rect 70 5835 90 5855
rect 110 5835 130 5855
rect 150 5835 170 5855
rect 190 5835 210 5855
rect 230 5835 250 5855
rect 270 5835 290 5855
rect 310 5835 330 5855
rect 350 5835 370 5855
rect 390 5835 410 5855
rect 440 5835 455 5855
rect -2045 5820 455 5835
rect -5595 5760 -3095 5775
rect -5595 5740 -5580 5760
rect -5550 5740 -5530 5760
rect -5510 5740 -5490 5760
rect -5470 5740 -5450 5760
rect -5430 5740 -5410 5760
rect -5390 5740 -5370 5760
rect -5350 5740 -5330 5760
rect -5310 5740 -5290 5760
rect -5270 5740 -5250 5760
rect -5230 5740 -5210 5760
rect -5190 5740 -5170 5760
rect -5150 5740 -5130 5760
rect -5110 5740 -5090 5760
rect -5070 5740 -5050 5760
rect -5030 5740 -5010 5760
rect -4990 5740 -4970 5760
rect -4950 5740 -4930 5760
rect -4910 5740 -4890 5760
rect -4870 5740 -4850 5760
rect -4830 5740 -4810 5760
rect -4790 5740 -4770 5760
rect -4750 5740 -4730 5760
rect -4710 5740 -4690 5760
rect -4670 5740 -4650 5760
rect -4630 5740 -4610 5760
rect -4590 5740 -4570 5760
rect -4550 5740 -4530 5760
rect -4510 5740 -4490 5760
rect -4470 5740 -4450 5760
rect -4430 5740 -4410 5760
rect -4390 5740 -4370 5760
rect -4350 5740 -4330 5760
rect -4310 5740 -4290 5760
rect -4270 5740 -4250 5760
rect -4230 5740 -4210 5760
rect -4190 5740 -4170 5760
rect -4150 5740 -4130 5760
rect -4110 5740 -4090 5760
rect -4070 5740 -4050 5760
rect -4030 5740 -4010 5760
rect -3990 5740 -3970 5760
rect -3950 5740 -3930 5760
rect -3910 5740 -3890 5760
rect -3870 5740 -3850 5760
rect -3830 5740 -3810 5760
rect -3790 5740 -3770 5760
rect -3750 5740 -3730 5760
rect -3710 5740 -3690 5760
rect -3670 5740 -3650 5760
rect -3630 5740 -3610 5760
rect -3590 5740 -3570 5760
rect -3550 5740 -3530 5760
rect -3510 5740 -3490 5760
rect -3470 5740 -3450 5760
rect -3430 5740 -3410 5760
rect -3390 5740 -3370 5760
rect -3350 5740 -3330 5760
rect -3310 5740 -3290 5760
rect -3270 5740 -3250 5760
rect -3230 5740 -3210 5760
rect -3190 5740 -3170 5760
rect -3150 5740 -3130 5760
rect -3110 5740 -3095 5760
rect -5595 5725 -3095 5740
rect -2045 5760 455 5775
rect -2045 5740 -2030 5760
rect -2010 5740 -1990 5760
rect -1970 5740 -1950 5760
rect -1930 5740 -1910 5760
rect -1890 5740 -1870 5760
rect -1850 5740 -1830 5760
rect -1810 5740 -1790 5760
rect -1770 5740 -1750 5760
rect -1730 5740 -1710 5760
rect -1690 5740 -1670 5760
rect -1650 5740 -1630 5760
rect -1610 5740 -1590 5760
rect -1570 5740 -1550 5760
rect -1530 5740 -1510 5760
rect -1490 5740 -1470 5760
rect -1450 5740 -1430 5760
rect -1410 5740 -1390 5760
rect -1370 5740 -1350 5760
rect -1330 5740 -1310 5760
rect -1290 5740 -1270 5760
rect -1250 5740 -1230 5760
rect -1210 5740 -1190 5760
rect -1170 5740 -1150 5760
rect -1130 5740 -1110 5760
rect -1090 5740 -1070 5760
rect -1050 5740 -1030 5760
rect -1010 5740 -990 5760
rect -970 5740 -950 5760
rect -930 5740 -910 5760
rect -890 5740 -870 5760
rect -850 5740 -830 5760
rect -810 5740 -790 5760
rect -770 5740 -750 5760
rect -730 5740 -710 5760
rect -690 5740 -670 5760
rect -650 5740 -630 5760
rect -610 5740 -590 5760
rect -570 5740 -550 5760
rect -530 5740 -510 5760
rect -490 5740 -470 5760
rect -450 5740 -430 5760
rect -410 5740 -390 5760
rect -370 5740 -350 5760
rect -330 5740 -310 5760
rect -290 5740 -270 5760
rect -250 5740 -230 5760
rect -210 5740 -190 5760
rect -170 5740 -150 5760
rect -130 5740 -110 5760
rect -90 5740 -70 5760
rect -50 5740 -30 5760
rect -10 5740 10 5760
rect 30 5740 50 5760
rect 70 5740 90 5760
rect 110 5740 130 5760
rect 150 5740 170 5760
rect 190 5740 210 5760
rect 230 5740 250 5760
rect 270 5740 290 5760
rect 310 5740 330 5760
rect 350 5740 370 5760
rect 390 5740 410 5760
rect 440 5740 455 5760
rect -2045 5725 455 5740
rect -5595 5665 -3095 5680
rect -5595 5645 -5580 5665
rect -5550 5645 -5530 5665
rect -5510 5645 -5490 5665
rect -5470 5645 -5450 5665
rect -5430 5645 -5410 5665
rect -5390 5645 -5370 5665
rect -5350 5645 -5330 5665
rect -5310 5645 -5290 5665
rect -5270 5645 -5250 5665
rect -5230 5645 -5210 5665
rect -5190 5645 -5170 5665
rect -5150 5645 -5130 5665
rect -5110 5645 -5090 5665
rect -5070 5645 -5050 5665
rect -5030 5645 -5010 5665
rect -4990 5645 -4970 5665
rect -4950 5645 -4930 5665
rect -4910 5645 -4890 5665
rect -4870 5645 -4850 5665
rect -4830 5645 -4810 5665
rect -4790 5645 -4770 5665
rect -4750 5645 -4730 5665
rect -4710 5645 -4690 5665
rect -4670 5645 -4650 5665
rect -4630 5645 -4610 5665
rect -4590 5645 -4570 5665
rect -4550 5645 -4530 5665
rect -4510 5645 -4490 5665
rect -4470 5645 -4450 5665
rect -4430 5645 -4410 5665
rect -4390 5645 -4370 5665
rect -4350 5645 -4330 5665
rect -4310 5645 -4290 5665
rect -4270 5645 -4250 5665
rect -4230 5645 -4210 5665
rect -4190 5645 -4170 5665
rect -4150 5645 -4130 5665
rect -4110 5645 -4090 5665
rect -4070 5645 -4050 5665
rect -4030 5645 -4010 5665
rect -3990 5645 -3970 5665
rect -3950 5645 -3930 5665
rect -3910 5645 -3890 5665
rect -3870 5645 -3850 5665
rect -3830 5645 -3810 5665
rect -3790 5645 -3770 5665
rect -3750 5645 -3730 5665
rect -3710 5645 -3690 5665
rect -3670 5645 -3650 5665
rect -3630 5645 -3610 5665
rect -3590 5645 -3570 5665
rect -3550 5645 -3530 5665
rect -3510 5645 -3490 5665
rect -3470 5645 -3450 5665
rect -3430 5645 -3410 5665
rect -3390 5645 -3370 5665
rect -3350 5645 -3330 5665
rect -3310 5645 -3290 5665
rect -3270 5645 -3250 5665
rect -3230 5645 -3210 5665
rect -3190 5645 -3170 5665
rect -3150 5645 -3130 5665
rect -3110 5645 -3095 5665
rect -5595 5630 -3095 5645
rect -2045 5665 455 5680
rect -2045 5645 -2030 5665
rect -2010 5645 -1990 5665
rect -1970 5645 -1950 5665
rect -1930 5645 -1910 5665
rect -1890 5645 -1870 5665
rect -1850 5645 -1830 5665
rect -1810 5645 -1790 5665
rect -1770 5645 -1750 5665
rect -1730 5645 -1710 5665
rect -1690 5645 -1670 5665
rect -1650 5645 -1630 5665
rect -1610 5645 -1590 5665
rect -1570 5645 -1550 5665
rect -1530 5645 -1510 5665
rect -1490 5645 -1470 5665
rect -1450 5645 -1430 5665
rect -1410 5645 -1390 5665
rect -1370 5645 -1350 5665
rect -1330 5645 -1310 5665
rect -1290 5645 -1270 5665
rect -1250 5645 -1230 5665
rect -1210 5645 -1190 5665
rect -1170 5645 -1150 5665
rect -1130 5645 -1110 5665
rect -1090 5645 -1070 5665
rect -1050 5645 -1030 5665
rect -1010 5645 -990 5665
rect -970 5645 -950 5665
rect -930 5645 -910 5665
rect -890 5645 -870 5665
rect -850 5645 -830 5665
rect -810 5645 -790 5665
rect -770 5645 -750 5665
rect -730 5645 -710 5665
rect -690 5645 -670 5665
rect -650 5645 -630 5665
rect -610 5645 -590 5665
rect -570 5645 -550 5665
rect -530 5645 -510 5665
rect -490 5645 -470 5665
rect -450 5645 -430 5665
rect -410 5645 -390 5665
rect -370 5645 -350 5665
rect -330 5645 -310 5665
rect -290 5645 -270 5665
rect -250 5645 -230 5665
rect -210 5645 -190 5665
rect -170 5645 -150 5665
rect -130 5645 -110 5665
rect -90 5645 -70 5665
rect -50 5645 -30 5665
rect -10 5645 10 5665
rect 30 5645 50 5665
rect 70 5645 90 5665
rect 110 5645 130 5665
rect 150 5645 170 5665
rect 190 5645 210 5665
rect 230 5645 250 5665
rect 270 5645 290 5665
rect 310 5645 330 5665
rect 350 5645 370 5665
rect 390 5645 410 5665
rect 440 5645 455 5665
rect -2045 5630 455 5645
rect -5595 5570 -3095 5585
rect -5595 5550 -5580 5570
rect -5550 5550 -5530 5570
rect -5510 5550 -5490 5570
rect -5470 5550 -5450 5570
rect -5430 5550 -5410 5570
rect -5390 5550 -5370 5570
rect -5350 5550 -5330 5570
rect -5310 5550 -5290 5570
rect -5270 5550 -5250 5570
rect -5230 5550 -5210 5570
rect -5190 5550 -5170 5570
rect -5150 5550 -5130 5570
rect -5110 5550 -5090 5570
rect -5070 5550 -5050 5570
rect -5030 5550 -5010 5570
rect -4990 5550 -4970 5570
rect -4950 5550 -4930 5570
rect -4910 5550 -4890 5570
rect -4870 5550 -4850 5570
rect -4830 5550 -4810 5570
rect -4790 5550 -4770 5570
rect -4750 5550 -4730 5570
rect -4710 5550 -4690 5570
rect -4670 5550 -4650 5570
rect -4630 5550 -4610 5570
rect -4590 5550 -4570 5570
rect -4550 5550 -4530 5570
rect -4510 5550 -4490 5570
rect -4470 5550 -4450 5570
rect -4430 5550 -4410 5570
rect -4390 5550 -4370 5570
rect -4350 5550 -4330 5570
rect -4310 5550 -4290 5570
rect -4270 5550 -4250 5570
rect -4230 5550 -4210 5570
rect -4190 5550 -4170 5570
rect -4150 5550 -4130 5570
rect -4110 5550 -4090 5570
rect -4070 5550 -4050 5570
rect -4030 5550 -4010 5570
rect -3990 5550 -3970 5570
rect -3950 5550 -3930 5570
rect -3910 5550 -3890 5570
rect -3870 5550 -3850 5570
rect -3830 5550 -3810 5570
rect -3790 5550 -3770 5570
rect -3750 5550 -3730 5570
rect -3710 5550 -3690 5570
rect -3670 5550 -3650 5570
rect -3630 5550 -3610 5570
rect -3590 5550 -3570 5570
rect -3550 5550 -3530 5570
rect -3510 5550 -3490 5570
rect -3470 5550 -3450 5570
rect -3430 5550 -3410 5570
rect -3390 5550 -3370 5570
rect -3350 5550 -3330 5570
rect -3310 5550 -3290 5570
rect -3270 5550 -3250 5570
rect -3230 5550 -3210 5570
rect -3190 5550 -3170 5570
rect -3150 5550 -3130 5570
rect -3110 5550 -3095 5570
rect -5595 5535 -3095 5550
rect -2045 5570 455 5585
rect -2045 5550 -2030 5570
rect -2010 5550 -1990 5570
rect -1970 5550 -1950 5570
rect -1930 5550 -1910 5570
rect -1890 5550 -1870 5570
rect -1850 5550 -1830 5570
rect -1810 5550 -1790 5570
rect -1770 5550 -1750 5570
rect -1730 5550 -1710 5570
rect -1690 5550 -1670 5570
rect -1650 5550 -1630 5570
rect -1610 5550 -1590 5570
rect -1570 5550 -1550 5570
rect -1530 5550 -1510 5570
rect -1490 5550 -1470 5570
rect -1450 5550 -1430 5570
rect -1410 5550 -1390 5570
rect -1370 5550 -1350 5570
rect -1330 5550 -1310 5570
rect -1290 5550 -1270 5570
rect -1250 5550 -1230 5570
rect -1210 5550 -1190 5570
rect -1170 5550 -1150 5570
rect -1130 5550 -1110 5570
rect -1090 5550 -1070 5570
rect -1050 5550 -1030 5570
rect -1010 5550 -990 5570
rect -970 5550 -950 5570
rect -930 5550 -910 5570
rect -890 5550 -870 5570
rect -850 5550 -830 5570
rect -810 5550 -790 5570
rect -770 5550 -750 5570
rect -730 5550 -710 5570
rect -690 5550 -670 5570
rect -650 5550 -630 5570
rect -610 5550 -590 5570
rect -570 5550 -550 5570
rect -530 5550 -510 5570
rect -490 5550 -470 5570
rect -450 5550 -430 5570
rect -410 5550 -390 5570
rect -370 5550 -350 5570
rect -330 5550 -310 5570
rect -290 5550 -270 5570
rect -250 5550 -230 5570
rect -210 5550 -190 5570
rect -170 5550 -150 5570
rect -130 5550 -110 5570
rect -90 5550 -70 5570
rect -50 5550 -30 5570
rect -10 5550 10 5570
rect 30 5550 50 5570
rect 70 5550 90 5570
rect 110 5550 130 5570
rect 150 5550 170 5570
rect 190 5550 210 5570
rect 230 5550 250 5570
rect 270 5550 290 5570
rect 310 5550 330 5570
rect 350 5550 370 5570
rect 390 5550 410 5570
rect 440 5550 455 5570
rect -2045 5535 455 5550
rect -5595 5475 -3095 5490
rect -5595 5455 -5580 5475
rect -5550 5455 -5530 5475
rect -5510 5455 -5490 5475
rect -5470 5455 -5450 5475
rect -5430 5455 -5410 5475
rect -5390 5455 -5370 5475
rect -5350 5455 -5330 5475
rect -5310 5455 -5290 5475
rect -5270 5455 -5250 5475
rect -5230 5455 -5210 5475
rect -5190 5455 -5170 5475
rect -5150 5455 -5130 5475
rect -5110 5455 -5090 5475
rect -5070 5455 -5050 5475
rect -5030 5455 -5010 5475
rect -4990 5455 -4970 5475
rect -4950 5455 -4930 5475
rect -4910 5455 -4890 5475
rect -4870 5455 -4850 5475
rect -4830 5455 -4810 5475
rect -4790 5455 -4770 5475
rect -4750 5455 -4730 5475
rect -4710 5455 -4690 5475
rect -4670 5455 -4650 5475
rect -4630 5455 -4610 5475
rect -4590 5455 -4570 5475
rect -4550 5455 -4530 5475
rect -4510 5455 -4490 5475
rect -4470 5455 -4450 5475
rect -4430 5455 -4410 5475
rect -4390 5455 -4370 5475
rect -4350 5455 -4330 5475
rect -4310 5455 -4290 5475
rect -4270 5455 -4250 5475
rect -4230 5455 -4210 5475
rect -4190 5455 -4170 5475
rect -4150 5455 -4130 5475
rect -4110 5455 -4090 5475
rect -4070 5455 -4050 5475
rect -4030 5455 -4010 5475
rect -3990 5455 -3970 5475
rect -3950 5455 -3930 5475
rect -3910 5455 -3890 5475
rect -3870 5455 -3850 5475
rect -3830 5455 -3810 5475
rect -3790 5455 -3770 5475
rect -3750 5455 -3730 5475
rect -3710 5455 -3690 5475
rect -3670 5455 -3650 5475
rect -3630 5455 -3610 5475
rect -3590 5455 -3570 5475
rect -3550 5455 -3530 5475
rect -3510 5455 -3490 5475
rect -3470 5455 -3450 5475
rect -3430 5455 -3410 5475
rect -3390 5455 -3370 5475
rect -3350 5455 -3330 5475
rect -3310 5455 -3290 5475
rect -3270 5455 -3250 5475
rect -3230 5455 -3210 5475
rect -3190 5455 -3170 5475
rect -3150 5455 -3130 5475
rect -3110 5455 -3095 5475
rect -5595 5440 -3095 5455
rect -2045 5475 455 5490
rect -2045 5455 -2030 5475
rect -2010 5455 -1990 5475
rect -1970 5455 -1950 5475
rect -1930 5455 -1910 5475
rect -1890 5455 -1870 5475
rect -1850 5455 -1830 5475
rect -1810 5455 -1790 5475
rect -1770 5455 -1750 5475
rect -1730 5455 -1710 5475
rect -1690 5455 -1670 5475
rect -1650 5455 -1630 5475
rect -1610 5455 -1590 5475
rect -1570 5455 -1550 5475
rect -1530 5455 -1510 5475
rect -1490 5455 -1470 5475
rect -1450 5455 -1430 5475
rect -1410 5455 -1390 5475
rect -1370 5455 -1350 5475
rect -1330 5455 -1310 5475
rect -1290 5455 -1270 5475
rect -1250 5455 -1230 5475
rect -1210 5455 -1190 5475
rect -1170 5455 -1150 5475
rect -1130 5455 -1110 5475
rect -1090 5455 -1070 5475
rect -1050 5455 -1030 5475
rect -1010 5455 -990 5475
rect -970 5455 -950 5475
rect -930 5455 -910 5475
rect -890 5455 -870 5475
rect -850 5455 -830 5475
rect -810 5455 -790 5475
rect -770 5455 -750 5475
rect -730 5455 -710 5475
rect -690 5455 -670 5475
rect -650 5455 -630 5475
rect -610 5455 -590 5475
rect -570 5455 -550 5475
rect -530 5455 -510 5475
rect -490 5455 -470 5475
rect -450 5455 -430 5475
rect -410 5455 -390 5475
rect -370 5455 -350 5475
rect -330 5455 -310 5475
rect -290 5455 -270 5475
rect -250 5455 -230 5475
rect -210 5455 -190 5475
rect -170 5455 -150 5475
rect -130 5455 -110 5475
rect -90 5455 -70 5475
rect -50 5455 -30 5475
rect -10 5455 10 5475
rect 30 5455 50 5475
rect 70 5455 90 5475
rect 110 5455 130 5475
rect 150 5455 170 5475
rect 190 5455 210 5475
rect 230 5455 250 5475
rect 270 5455 290 5475
rect 310 5455 330 5475
rect 350 5455 370 5475
rect 390 5455 410 5475
rect 440 5455 455 5475
rect -2045 5440 455 5455
rect -5595 5380 -3095 5395
rect -5595 5360 -5580 5380
rect -5550 5360 -5530 5380
rect -5510 5360 -5490 5380
rect -5470 5360 -5450 5380
rect -5430 5360 -5410 5380
rect -5390 5360 -5370 5380
rect -5350 5360 -5330 5380
rect -5310 5360 -5290 5380
rect -5270 5360 -5250 5380
rect -5230 5360 -5210 5380
rect -5190 5360 -5170 5380
rect -5150 5360 -5130 5380
rect -5110 5360 -5090 5380
rect -5070 5360 -5050 5380
rect -5030 5360 -5010 5380
rect -4990 5360 -4970 5380
rect -4950 5360 -4930 5380
rect -4910 5360 -4890 5380
rect -4870 5360 -4850 5380
rect -4830 5360 -4810 5380
rect -4790 5360 -4770 5380
rect -4750 5360 -4730 5380
rect -4710 5360 -4690 5380
rect -4670 5360 -4650 5380
rect -4630 5360 -4610 5380
rect -4590 5360 -4570 5380
rect -4550 5360 -4530 5380
rect -4510 5360 -4490 5380
rect -4470 5360 -4450 5380
rect -4430 5360 -4410 5380
rect -4390 5360 -4370 5380
rect -4350 5360 -4330 5380
rect -4310 5360 -4290 5380
rect -4270 5360 -4250 5380
rect -4230 5360 -4210 5380
rect -4190 5360 -4170 5380
rect -4150 5360 -4130 5380
rect -4110 5360 -4090 5380
rect -4070 5360 -4050 5380
rect -4030 5360 -4010 5380
rect -3990 5360 -3970 5380
rect -3950 5360 -3930 5380
rect -3910 5360 -3890 5380
rect -3870 5360 -3850 5380
rect -3830 5360 -3810 5380
rect -3790 5360 -3770 5380
rect -3750 5360 -3730 5380
rect -3710 5360 -3690 5380
rect -3670 5360 -3650 5380
rect -3630 5360 -3610 5380
rect -3590 5360 -3570 5380
rect -3550 5360 -3530 5380
rect -3510 5360 -3490 5380
rect -3470 5360 -3450 5380
rect -3430 5360 -3410 5380
rect -3390 5360 -3370 5380
rect -3350 5360 -3330 5380
rect -3310 5360 -3290 5380
rect -3270 5360 -3250 5380
rect -3230 5360 -3210 5380
rect -3190 5360 -3170 5380
rect -3150 5360 -3130 5380
rect -3110 5360 -3095 5380
rect -5595 5345 -3095 5360
rect -2045 5380 455 5395
rect -2045 5360 -2030 5380
rect -2010 5360 -1990 5380
rect -1970 5360 -1950 5380
rect -1930 5360 -1910 5380
rect -1890 5360 -1870 5380
rect -1850 5360 -1830 5380
rect -1810 5360 -1790 5380
rect -1770 5360 -1750 5380
rect -1730 5360 -1710 5380
rect -1690 5360 -1670 5380
rect -1650 5360 -1630 5380
rect -1610 5360 -1590 5380
rect -1570 5360 -1550 5380
rect -1530 5360 -1510 5380
rect -1490 5360 -1470 5380
rect -1450 5360 -1430 5380
rect -1410 5360 -1390 5380
rect -1370 5360 -1350 5380
rect -1330 5360 -1310 5380
rect -1290 5360 -1270 5380
rect -1250 5360 -1230 5380
rect -1210 5360 -1190 5380
rect -1170 5360 -1150 5380
rect -1130 5360 -1110 5380
rect -1090 5360 -1070 5380
rect -1050 5360 -1030 5380
rect -1010 5360 -990 5380
rect -970 5360 -950 5380
rect -930 5360 -910 5380
rect -890 5360 -870 5380
rect -850 5360 -830 5380
rect -810 5360 -790 5380
rect -770 5360 -750 5380
rect -730 5360 -710 5380
rect -690 5360 -670 5380
rect -650 5360 -630 5380
rect -610 5360 -590 5380
rect -570 5360 -550 5380
rect -530 5360 -510 5380
rect -490 5360 -470 5380
rect -450 5360 -430 5380
rect -410 5360 -390 5380
rect -370 5360 -350 5380
rect -330 5360 -310 5380
rect -290 5360 -270 5380
rect -250 5360 -230 5380
rect -210 5360 -190 5380
rect -170 5360 -150 5380
rect -130 5360 -110 5380
rect -90 5360 -70 5380
rect -50 5360 -30 5380
rect -10 5360 10 5380
rect 30 5360 50 5380
rect 70 5360 90 5380
rect 110 5360 130 5380
rect 150 5360 170 5380
rect 190 5360 210 5380
rect 230 5360 250 5380
rect 270 5360 290 5380
rect 310 5360 330 5380
rect 350 5360 370 5380
rect 390 5360 410 5380
rect 440 5360 455 5380
rect -2045 5345 455 5360
rect -5595 5285 -3095 5300
rect -5595 5265 -5580 5285
rect -5550 5265 -5530 5285
rect -5510 5265 -5490 5285
rect -5470 5265 -5450 5285
rect -5430 5265 -5410 5285
rect -5390 5265 -5370 5285
rect -5350 5265 -5330 5285
rect -5310 5265 -5290 5285
rect -5270 5265 -5250 5285
rect -5230 5265 -5210 5285
rect -5190 5265 -5170 5285
rect -5150 5265 -5130 5285
rect -5110 5265 -5090 5285
rect -5070 5265 -5050 5285
rect -5030 5265 -5010 5285
rect -4990 5265 -4970 5285
rect -4950 5265 -4930 5285
rect -4910 5265 -4890 5285
rect -4870 5265 -4850 5285
rect -4830 5265 -4810 5285
rect -4790 5265 -4770 5285
rect -4750 5265 -4730 5285
rect -4710 5265 -4690 5285
rect -4670 5265 -4650 5285
rect -4630 5265 -4610 5285
rect -4590 5265 -4570 5285
rect -4550 5265 -4530 5285
rect -4510 5265 -4490 5285
rect -4470 5265 -4450 5285
rect -4430 5265 -4410 5285
rect -4390 5265 -4370 5285
rect -4350 5265 -4330 5285
rect -4310 5265 -4290 5285
rect -4270 5265 -4250 5285
rect -4230 5265 -4210 5285
rect -4190 5265 -4170 5285
rect -4150 5265 -4130 5285
rect -4110 5265 -4090 5285
rect -4070 5265 -4050 5285
rect -4030 5265 -4010 5285
rect -3990 5265 -3970 5285
rect -3950 5265 -3930 5285
rect -3910 5265 -3890 5285
rect -3870 5265 -3850 5285
rect -3830 5265 -3810 5285
rect -3790 5265 -3770 5285
rect -3750 5265 -3730 5285
rect -3710 5265 -3690 5285
rect -3670 5265 -3650 5285
rect -3630 5265 -3610 5285
rect -3590 5265 -3570 5285
rect -3550 5265 -3530 5285
rect -3510 5265 -3490 5285
rect -3470 5265 -3450 5285
rect -3430 5265 -3410 5285
rect -3390 5265 -3370 5285
rect -3350 5265 -3330 5285
rect -3310 5265 -3290 5285
rect -3270 5265 -3250 5285
rect -3230 5265 -3210 5285
rect -3190 5265 -3170 5285
rect -3150 5265 -3130 5285
rect -3110 5265 -3095 5285
rect -5595 5250 -3095 5265
rect -2045 5285 455 5300
rect -2045 5265 -2030 5285
rect -2010 5265 -1990 5285
rect -1970 5265 -1950 5285
rect -1930 5265 -1910 5285
rect -1890 5265 -1870 5285
rect -1850 5265 -1830 5285
rect -1810 5265 -1790 5285
rect -1770 5265 -1750 5285
rect -1730 5265 -1710 5285
rect -1690 5265 -1670 5285
rect -1650 5265 -1630 5285
rect -1610 5265 -1590 5285
rect -1570 5265 -1550 5285
rect -1530 5265 -1510 5285
rect -1490 5265 -1470 5285
rect -1450 5265 -1430 5285
rect -1410 5265 -1390 5285
rect -1370 5265 -1350 5285
rect -1330 5265 -1310 5285
rect -1290 5265 -1270 5285
rect -1250 5265 -1230 5285
rect -1210 5265 -1190 5285
rect -1170 5265 -1150 5285
rect -1130 5265 -1110 5285
rect -1090 5265 -1070 5285
rect -1050 5265 -1030 5285
rect -1010 5265 -990 5285
rect -970 5265 -950 5285
rect -930 5265 -910 5285
rect -890 5265 -870 5285
rect -850 5265 -830 5285
rect -810 5265 -790 5285
rect -770 5265 -750 5285
rect -730 5265 -710 5285
rect -690 5265 -670 5285
rect -650 5265 -630 5285
rect -610 5265 -590 5285
rect -570 5265 -550 5285
rect -530 5265 -510 5285
rect -490 5265 -470 5285
rect -450 5265 -430 5285
rect -410 5265 -390 5285
rect -370 5265 -350 5285
rect -330 5265 -310 5285
rect -290 5265 -270 5285
rect -250 5265 -230 5285
rect -210 5265 -190 5285
rect -170 5265 -150 5285
rect -130 5265 -110 5285
rect -90 5265 -70 5285
rect -50 5265 -30 5285
rect -10 5265 10 5285
rect 30 5265 50 5285
rect 70 5265 90 5285
rect 110 5265 130 5285
rect 150 5265 170 5285
rect 190 5265 210 5285
rect 230 5265 250 5285
rect 270 5265 290 5285
rect 310 5265 330 5285
rect 350 5265 370 5285
rect 390 5265 410 5285
rect 440 5265 455 5285
rect -2045 5250 455 5265
rect -5595 5190 -3095 5205
rect -5595 5170 -5580 5190
rect -5550 5170 -5530 5190
rect -5510 5170 -5490 5190
rect -5470 5170 -5450 5190
rect -5430 5170 -5410 5190
rect -5390 5170 -5370 5190
rect -5350 5170 -5330 5190
rect -5310 5170 -5290 5190
rect -5270 5170 -5250 5190
rect -5230 5170 -5210 5190
rect -5190 5170 -5170 5190
rect -5150 5170 -5130 5190
rect -5110 5170 -5090 5190
rect -5070 5170 -5050 5190
rect -5030 5170 -5010 5190
rect -4990 5170 -4970 5190
rect -4950 5170 -4930 5190
rect -4910 5170 -4890 5190
rect -4870 5170 -4850 5190
rect -4830 5170 -4810 5190
rect -4790 5170 -4770 5190
rect -4750 5170 -4730 5190
rect -4710 5170 -4690 5190
rect -4670 5170 -4650 5190
rect -4630 5170 -4610 5190
rect -4590 5170 -4570 5190
rect -4550 5170 -4530 5190
rect -4510 5170 -4490 5190
rect -4470 5170 -4450 5190
rect -4430 5170 -4410 5190
rect -4390 5170 -4370 5190
rect -4350 5170 -4330 5190
rect -4310 5170 -4290 5190
rect -4270 5170 -4250 5190
rect -4230 5170 -4210 5190
rect -4190 5170 -4170 5190
rect -4150 5170 -4130 5190
rect -4110 5170 -4090 5190
rect -4070 5170 -4050 5190
rect -4030 5170 -4010 5190
rect -3990 5170 -3970 5190
rect -3950 5170 -3930 5190
rect -3910 5170 -3890 5190
rect -3870 5170 -3850 5190
rect -3830 5170 -3810 5190
rect -3790 5170 -3770 5190
rect -3750 5170 -3730 5190
rect -3710 5170 -3690 5190
rect -3670 5170 -3650 5190
rect -3630 5170 -3610 5190
rect -3590 5170 -3570 5190
rect -3550 5170 -3530 5190
rect -3510 5170 -3490 5190
rect -3470 5170 -3450 5190
rect -3430 5170 -3410 5190
rect -3390 5170 -3370 5190
rect -3350 5170 -3330 5190
rect -3310 5170 -3290 5190
rect -3270 5170 -3250 5190
rect -3230 5170 -3210 5190
rect -3190 5170 -3170 5190
rect -3150 5170 -3130 5190
rect -3110 5170 -3095 5190
rect -5595 5155 -3095 5170
rect -2045 5190 455 5205
rect -2045 5170 -2030 5190
rect -2010 5170 -1990 5190
rect -1970 5170 -1950 5190
rect -1930 5170 -1910 5190
rect -1890 5170 -1870 5190
rect -1850 5170 -1830 5190
rect -1810 5170 -1790 5190
rect -1770 5170 -1750 5190
rect -1730 5170 -1710 5190
rect -1690 5170 -1670 5190
rect -1650 5170 -1630 5190
rect -1610 5170 -1590 5190
rect -1570 5170 -1550 5190
rect -1530 5170 -1510 5190
rect -1490 5170 -1470 5190
rect -1450 5170 -1430 5190
rect -1410 5170 -1390 5190
rect -1370 5170 -1350 5190
rect -1330 5170 -1310 5190
rect -1290 5170 -1270 5190
rect -1250 5170 -1230 5190
rect -1210 5170 -1190 5190
rect -1170 5170 -1150 5190
rect -1130 5170 -1110 5190
rect -1090 5170 -1070 5190
rect -1050 5170 -1030 5190
rect -1010 5170 -990 5190
rect -970 5170 -950 5190
rect -930 5170 -910 5190
rect -890 5170 -870 5190
rect -850 5170 -830 5190
rect -810 5170 -790 5190
rect -770 5170 -750 5190
rect -730 5170 -710 5190
rect -690 5170 -670 5190
rect -650 5170 -630 5190
rect -610 5170 -590 5190
rect -570 5170 -550 5190
rect -530 5170 -510 5190
rect -490 5170 -470 5190
rect -450 5170 -430 5190
rect -410 5170 -390 5190
rect -370 5170 -350 5190
rect -330 5170 -310 5190
rect -290 5170 -270 5190
rect -250 5170 -230 5190
rect -210 5170 -190 5190
rect -170 5170 -150 5190
rect -130 5170 -110 5190
rect -90 5170 -70 5190
rect -50 5170 -30 5190
rect -10 5170 10 5190
rect 30 5170 50 5190
rect 70 5170 90 5190
rect 110 5170 130 5190
rect 150 5170 170 5190
rect 190 5170 210 5190
rect 230 5170 250 5190
rect 270 5170 290 5190
rect 310 5170 330 5190
rect 350 5170 370 5190
rect 390 5170 410 5190
rect 440 5170 455 5190
rect -2045 5155 455 5170
rect -5595 5095 -3095 5110
rect -5595 5075 -5580 5095
rect -5550 5075 -5530 5095
rect -5510 5075 -5490 5095
rect -5470 5075 -5450 5095
rect -5430 5075 -5410 5095
rect -5390 5075 -5370 5095
rect -5350 5075 -5330 5095
rect -5310 5075 -5290 5095
rect -5270 5075 -5250 5095
rect -5230 5075 -5210 5095
rect -5190 5075 -5170 5095
rect -5150 5075 -5130 5095
rect -5110 5075 -5090 5095
rect -5070 5075 -5050 5095
rect -5030 5075 -5010 5095
rect -4990 5075 -4970 5095
rect -4950 5075 -4930 5095
rect -4910 5075 -4890 5095
rect -4870 5075 -4850 5095
rect -4830 5075 -4810 5095
rect -4790 5075 -4770 5095
rect -4750 5075 -4730 5095
rect -4710 5075 -4690 5095
rect -4670 5075 -4650 5095
rect -4630 5075 -4610 5095
rect -4590 5075 -4570 5095
rect -4550 5075 -4530 5095
rect -4510 5075 -4490 5095
rect -4470 5075 -4450 5095
rect -4430 5075 -4410 5095
rect -4390 5075 -4370 5095
rect -4350 5075 -4330 5095
rect -4310 5075 -4290 5095
rect -4270 5075 -4250 5095
rect -4230 5075 -4210 5095
rect -4190 5075 -4170 5095
rect -4150 5075 -4130 5095
rect -4110 5075 -4090 5095
rect -4070 5075 -4050 5095
rect -4030 5075 -4010 5095
rect -3990 5075 -3970 5095
rect -3950 5075 -3930 5095
rect -3910 5075 -3890 5095
rect -3870 5075 -3850 5095
rect -3830 5075 -3810 5095
rect -3790 5075 -3770 5095
rect -3750 5075 -3730 5095
rect -3710 5075 -3690 5095
rect -3670 5075 -3650 5095
rect -3630 5075 -3610 5095
rect -3590 5075 -3570 5095
rect -3550 5075 -3530 5095
rect -3510 5075 -3490 5095
rect -3470 5075 -3450 5095
rect -3430 5075 -3410 5095
rect -3390 5075 -3370 5095
rect -3350 5075 -3330 5095
rect -3310 5075 -3290 5095
rect -3270 5075 -3250 5095
rect -3230 5075 -3210 5095
rect -3190 5075 -3170 5095
rect -3150 5075 -3130 5095
rect -3110 5075 -3095 5095
rect -5595 5060 -3095 5075
rect -2045 5095 455 5110
rect -2045 5075 -2030 5095
rect -2010 5075 -1990 5095
rect -1970 5075 -1950 5095
rect -1930 5075 -1910 5095
rect -1890 5075 -1870 5095
rect -1850 5075 -1830 5095
rect -1810 5075 -1790 5095
rect -1770 5075 -1750 5095
rect -1730 5075 -1710 5095
rect -1690 5075 -1670 5095
rect -1650 5075 -1630 5095
rect -1610 5075 -1590 5095
rect -1570 5075 -1550 5095
rect -1530 5075 -1510 5095
rect -1490 5075 -1470 5095
rect -1450 5075 -1430 5095
rect -1410 5075 -1390 5095
rect -1370 5075 -1350 5095
rect -1330 5075 -1310 5095
rect -1290 5075 -1270 5095
rect -1250 5075 -1230 5095
rect -1210 5075 -1190 5095
rect -1170 5075 -1150 5095
rect -1130 5075 -1110 5095
rect -1090 5075 -1070 5095
rect -1050 5075 -1030 5095
rect -1010 5075 -990 5095
rect -970 5075 -950 5095
rect -930 5075 -910 5095
rect -890 5075 -870 5095
rect -850 5075 -830 5095
rect -810 5075 -790 5095
rect -770 5075 -750 5095
rect -730 5075 -710 5095
rect -690 5075 -670 5095
rect -650 5075 -630 5095
rect -610 5075 -590 5095
rect -570 5075 -550 5095
rect -530 5075 -510 5095
rect -490 5075 -470 5095
rect -450 5075 -430 5095
rect -410 5075 -390 5095
rect -370 5075 -350 5095
rect -330 5075 -310 5095
rect -290 5075 -270 5095
rect -250 5075 -230 5095
rect -210 5075 -190 5095
rect -170 5075 -150 5095
rect -130 5075 -110 5095
rect -90 5075 -70 5095
rect -50 5075 -30 5095
rect -10 5075 10 5095
rect 30 5075 50 5095
rect 70 5075 90 5095
rect 110 5075 130 5095
rect 150 5075 170 5095
rect 190 5075 210 5095
rect 230 5075 250 5095
rect 270 5075 290 5095
rect 310 5075 330 5095
rect 350 5075 370 5095
rect 390 5075 410 5095
rect 440 5075 455 5095
rect -2045 5060 455 5075
rect -5595 5000 -3095 5015
rect -5595 4980 -5580 5000
rect -5550 4980 -5530 5000
rect -5510 4980 -5490 5000
rect -5470 4980 -5450 5000
rect -5430 4980 -5410 5000
rect -5390 4980 -5370 5000
rect -5350 4980 -5330 5000
rect -5310 4980 -5290 5000
rect -5270 4980 -5250 5000
rect -5230 4980 -5210 5000
rect -5190 4980 -5170 5000
rect -5150 4980 -5130 5000
rect -5110 4980 -5090 5000
rect -5070 4980 -5050 5000
rect -5030 4980 -5010 5000
rect -4990 4980 -4970 5000
rect -4950 4980 -4930 5000
rect -4910 4980 -4890 5000
rect -4870 4980 -4850 5000
rect -4830 4980 -4810 5000
rect -4790 4980 -4770 5000
rect -4750 4980 -4730 5000
rect -4710 4980 -4690 5000
rect -4670 4980 -4650 5000
rect -4630 4980 -4610 5000
rect -4590 4980 -4570 5000
rect -4550 4980 -4530 5000
rect -4510 4980 -4490 5000
rect -4470 4980 -4450 5000
rect -4430 4980 -4410 5000
rect -4390 4980 -4370 5000
rect -4350 4980 -4330 5000
rect -4310 4980 -4290 5000
rect -4270 4980 -4250 5000
rect -4230 4980 -4210 5000
rect -4190 4980 -4170 5000
rect -4150 4980 -4130 5000
rect -4110 4980 -4090 5000
rect -4070 4980 -4050 5000
rect -4030 4980 -4010 5000
rect -3990 4980 -3970 5000
rect -3950 4980 -3930 5000
rect -3910 4980 -3890 5000
rect -3870 4980 -3850 5000
rect -3830 4980 -3810 5000
rect -3790 4980 -3770 5000
rect -3750 4980 -3730 5000
rect -3710 4980 -3690 5000
rect -3670 4980 -3650 5000
rect -3630 4980 -3610 5000
rect -3590 4980 -3570 5000
rect -3550 4980 -3530 5000
rect -3510 4980 -3490 5000
rect -3470 4980 -3450 5000
rect -3430 4980 -3410 5000
rect -3390 4980 -3370 5000
rect -3350 4980 -3330 5000
rect -3310 4980 -3290 5000
rect -3270 4980 -3250 5000
rect -3230 4980 -3210 5000
rect -3190 4980 -3170 5000
rect -3150 4980 -3130 5000
rect -3110 4980 -3095 5000
rect -5595 4965 -3095 4980
rect -2045 5000 455 5015
rect -2045 4980 -2030 5000
rect -2010 4980 -1990 5000
rect -1970 4980 -1950 5000
rect -1930 4980 -1910 5000
rect -1890 4980 -1870 5000
rect -1850 4980 -1830 5000
rect -1810 4980 -1790 5000
rect -1770 4980 -1750 5000
rect -1730 4980 -1710 5000
rect -1690 4980 -1670 5000
rect -1650 4980 -1630 5000
rect -1610 4980 -1590 5000
rect -1570 4980 -1550 5000
rect -1530 4980 -1510 5000
rect -1490 4980 -1470 5000
rect -1450 4980 -1430 5000
rect -1410 4980 -1390 5000
rect -1370 4980 -1350 5000
rect -1330 4980 -1310 5000
rect -1290 4980 -1270 5000
rect -1250 4980 -1230 5000
rect -1210 4980 -1190 5000
rect -1170 4980 -1150 5000
rect -1130 4980 -1110 5000
rect -1090 4980 -1070 5000
rect -1050 4980 -1030 5000
rect -1010 4980 -990 5000
rect -970 4980 -950 5000
rect -930 4980 -910 5000
rect -890 4980 -870 5000
rect -850 4980 -830 5000
rect -810 4980 -790 5000
rect -770 4980 -750 5000
rect -730 4980 -710 5000
rect -690 4980 -670 5000
rect -650 4980 -630 5000
rect -610 4980 -590 5000
rect -570 4980 -550 5000
rect -530 4980 -510 5000
rect -490 4980 -470 5000
rect -450 4980 -430 5000
rect -410 4980 -390 5000
rect -370 4980 -350 5000
rect -330 4980 -310 5000
rect -290 4980 -270 5000
rect -250 4980 -230 5000
rect -210 4980 -190 5000
rect -170 4980 -150 5000
rect -130 4980 -110 5000
rect -90 4980 -70 5000
rect -50 4980 -30 5000
rect -10 4980 10 5000
rect 30 4980 50 5000
rect 70 4980 90 5000
rect 110 4980 130 5000
rect 150 4980 170 5000
rect 190 4980 210 5000
rect 230 4980 250 5000
rect 270 4980 290 5000
rect 310 4980 330 5000
rect 350 4980 370 5000
rect 390 4980 410 5000
rect 440 4980 455 5000
rect -2045 4965 455 4980
rect -5595 4905 -3095 4920
rect -5595 4885 -5580 4905
rect -5550 4885 -5530 4905
rect -5510 4885 -5490 4905
rect -5470 4885 -5450 4905
rect -5430 4885 -5410 4905
rect -5390 4885 -5370 4905
rect -5350 4885 -5330 4905
rect -5310 4885 -5290 4905
rect -5270 4885 -5250 4905
rect -5230 4885 -5210 4905
rect -5190 4885 -5170 4905
rect -5150 4885 -5130 4905
rect -5110 4885 -5090 4905
rect -5070 4885 -5050 4905
rect -5030 4885 -5010 4905
rect -4990 4885 -4970 4905
rect -4950 4885 -4930 4905
rect -4910 4885 -4890 4905
rect -4870 4885 -4850 4905
rect -4830 4885 -4810 4905
rect -4790 4885 -4770 4905
rect -4750 4885 -4730 4905
rect -4710 4885 -4690 4905
rect -4670 4885 -4650 4905
rect -4630 4885 -4610 4905
rect -4590 4885 -4570 4905
rect -4550 4885 -4530 4905
rect -4510 4885 -4490 4905
rect -4470 4885 -4450 4905
rect -4430 4885 -4410 4905
rect -4390 4885 -4370 4905
rect -4350 4885 -4330 4905
rect -4310 4885 -4290 4905
rect -4270 4885 -4250 4905
rect -4230 4885 -4210 4905
rect -4190 4885 -4170 4905
rect -4150 4885 -4130 4905
rect -4110 4885 -4090 4905
rect -4070 4885 -4050 4905
rect -4030 4885 -4010 4905
rect -3990 4885 -3970 4905
rect -3950 4885 -3930 4905
rect -3910 4885 -3890 4905
rect -3870 4885 -3850 4905
rect -3830 4885 -3810 4905
rect -3790 4885 -3770 4905
rect -3750 4885 -3730 4905
rect -3710 4885 -3690 4905
rect -3670 4885 -3650 4905
rect -3630 4885 -3610 4905
rect -3590 4885 -3570 4905
rect -3550 4885 -3530 4905
rect -3510 4885 -3490 4905
rect -3470 4885 -3450 4905
rect -3430 4885 -3410 4905
rect -3390 4885 -3370 4905
rect -3350 4885 -3330 4905
rect -3310 4885 -3290 4905
rect -3270 4885 -3250 4905
rect -3230 4885 -3210 4905
rect -3190 4885 -3170 4905
rect -3150 4885 -3130 4905
rect -3110 4885 -3095 4905
rect -5595 4870 -3095 4885
rect -2045 4905 455 4920
rect -2045 4885 -2030 4905
rect -2010 4885 -1990 4905
rect -1970 4885 -1950 4905
rect -1930 4885 -1910 4905
rect -1890 4885 -1870 4905
rect -1850 4885 -1830 4905
rect -1810 4885 -1790 4905
rect -1770 4885 -1750 4905
rect -1730 4885 -1710 4905
rect -1690 4885 -1670 4905
rect -1650 4885 -1630 4905
rect -1610 4885 -1590 4905
rect -1570 4885 -1550 4905
rect -1530 4885 -1510 4905
rect -1490 4885 -1470 4905
rect -1450 4885 -1430 4905
rect -1410 4885 -1390 4905
rect -1370 4885 -1350 4905
rect -1330 4885 -1310 4905
rect -1290 4885 -1270 4905
rect -1250 4885 -1230 4905
rect -1210 4885 -1190 4905
rect -1170 4885 -1150 4905
rect -1130 4885 -1110 4905
rect -1090 4885 -1070 4905
rect -1050 4885 -1030 4905
rect -1010 4885 -990 4905
rect -970 4885 -950 4905
rect -930 4885 -910 4905
rect -890 4885 -870 4905
rect -850 4885 -830 4905
rect -810 4885 -790 4905
rect -770 4885 -750 4905
rect -730 4885 -710 4905
rect -690 4885 -670 4905
rect -650 4885 -630 4905
rect -610 4885 -590 4905
rect -570 4885 -550 4905
rect -530 4885 -510 4905
rect -490 4885 -470 4905
rect -450 4885 -430 4905
rect -410 4885 -390 4905
rect -370 4885 -350 4905
rect -330 4885 -310 4905
rect -290 4885 -270 4905
rect -250 4885 -230 4905
rect -210 4885 -190 4905
rect -170 4885 -150 4905
rect -130 4885 -110 4905
rect -90 4885 -70 4905
rect -50 4885 -30 4905
rect -10 4885 10 4905
rect 30 4885 50 4905
rect 70 4885 90 4905
rect 110 4885 130 4905
rect 150 4885 170 4905
rect 190 4885 210 4905
rect 230 4885 250 4905
rect 270 4885 290 4905
rect 310 4885 330 4905
rect 350 4885 370 4905
rect 390 4885 410 4905
rect 440 4885 455 4905
rect -2045 4870 455 4885
rect -5595 4810 -3095 4825
rect -5595 4790 -5580 4810
rect -5550 4790 -5530 4810
rect -5510 4790 -5490 4810
rect -5470 4790 -5450 4810
rect -5430 4790 -5410 4810
rect -5390 4790 -5370 4810
rect -5350 4790 -5330 4810
rect -5310 4790 -5290 4810
rect -5270 4790 -5250 4810
rect -5230 4790 -5210 4810
rect -5190 4790 -5170 4810
rect -5150 4790 -5130 4810
rect -5110 4790 -5090 4810
rect -5070 4790 -5050 4810
rect -5030 4790 -5010 4810
rect -4990 4790 -4970 4810
rect -4950 4790 -4930 4810
rect -4910 4790 -4890 4810
rect -4870 4790 -4850 4810
rect -4830 4790 -4810 4810
rect -4790 4790 -4770 4810
rect -4750 4790 -4730 4810
rect -4710 4790 -4690 4810
rect -4670 4790 -4650 4810
rect -4630 4790 -4610 4810
rect -4590 4790 -4570 4810
rect -4550 4790 -4530 4810
rect -4510 4790 -4490 4810
rect -4470 4790 -4450 4810
rect -4430 4790 -4410 4810
rect -4390 4790 -4370 4810
rect -4350 4790 -4330 4810
rect -4310 4790 -4290 4810
rect -4270 4790 -4250 4810
rect -4230 4790 -4210 4810
rect -4190 4790 -4170 4810
rect -4150 4790 -4130 4810
rect -4110 4790 -4090 4810
rect -4070 4790 -4050 4810
rect -4030 4790 -4010 4810
rect -3990 4790 -3970 4810
rect -3950 4790 -3930 4810
rect -3910 4790 -3890 4810
rect -3870 4790 -3850 4810
rect -3830 4790 -3810 4810
rect -3790 4790 -3770 4810
rect -3750 4790 -3730 4810
rect -3710 4790 -3690 4810
rect -3670 4790 -3650 4810
rect -3630 4790 -3610 4810
rect -3590 4790 -3570 4810
rect -3550 4790 -3530 4810
rect -3510 4790 -3490 4810
rect -3470 4790 -3450 4810
rect -3430 4790 -3410 4810
rect -3390 4790 -3370 4810
rect -3350 4790 -3330 4810
rect -3310 4790 -3290 4810
rect -3270 4790 -3250 4810
rect -3230 4790 -3210 4810
rect -3190 4790 -3170 4810
rect -3150 4790 -3130 4810
rect -3110 4790 -3095 4810
rect -5595 4775 -3095 4790
rect -2045 4810 455 4825
rect -2045 4790 -2030 4810
rect -2010 4790 -1990 4810
rect -1970 4790 -1950 4810
rect -1930 4790 -1910 4810
rect -1890 4790 -1870 4810
rect -1850 4790 -1830 4810
rect -1810 4790 -1790 4810
rect -1770 4790 -1750 4810
rect -1730 4790 -1710 4810
rect -1690 4790 -1670 4810
rect -1650 4790 -1630 4810
rect -1610 4790 -1590 4810
rect -1570 4790 -1550 4810
rect -1530 4790 -1510 4810
rect -1490 4790 -1470 4810
rect -1450 4790 -1430 4810
rect -1410 4790 -1390 4810
rect -1370 4790 -1350 4810
rect -1330 4790 -1310 4810
rect -1290 4790 -1270 4810
rect -1250 4790 -1230 4810
rect -1210 4790 -1190 4810
rect -1170 4790 -1150 4810
rect -1130 4790 -1110 4810
rect -1090 4790 -1070 4810
rect -1050 4790 -1030 4810
rect -1010 4790 -990 4810
rect -970 4790 -950 4810
rect -930 4790 -910 4810
rect -890 4790 -870 4810
rect -850 4790 -830 4810
rect -810 4790 -790 4810
rect -770 4790 -750 4810
rect -730 4790 -710 4810
rect -690 4790 -670 4810
rect -650 4790 -630 4810
rect -610 4790 -590 4810
rect -570 4790 -550 4810
rect -530 4790 -510 4810
rect -490 4790 -470 4810
rect -450 4790 -430 4810
rect -410 4790 -390 4810
rect -370 4790 -350 4810
rect -330 4790 -310 4810
rect -290 4790 -270 4810
rect -250 4790 -230 4810
rect -210 4790 -190 4810
rect -170 4790 -150 4810
rect -130 4790 -110 4810
rect -90 4790 -70 4810
rect -50 4790 -30 4810
rect -10 4790 10 4810
rect 30 4790 50 4810
rect 70 4790 90 4810
rect 110 4790 130 4810
rect 150 4790 170 4810
rect 190 4790 210 4810
rect 230 4790 250 4810
rect 270 4790 290 4810
rect 310 4790 330 4810
rect 350 4790 370 4810
rect 390 4790 410 4810
rect 440 4790 455 4810
rect -2045 4775 455 4790
rect -5595 4715 -3095 4730
rect -5595 4695 -5580 4715
rect -5550 4695 -5530 4715
rect -5510 4695 -5490 4715
rect -5470 4695 -5450 4715
rect -5430 4695 -5410 4715
rect -5390 4695 -5370 4715
rect -5350 4695 -5330 4715
rect -5310 4695 -5290 4715
rect -5270 4695 -5250 4715
rect -5230 4695 -5210 4715
rect -5190 4695 -5170 4715
rect -5150 4695 -5130 4715
rect -5110 4695 -5090 4715
rect -5070 4695 -5050 4715
rect -5030 4695 -5010 4715
rect -4990 4695 -4970 4715
rect -4950 4695 -4930 4715
rect -4910 4695 -4890 4715
rect -4870 4695 -4850 4715
rect -4830 4695 -4810 4715
rect -4790 4695 -4770 4715
rect -4750 4695 -4730 4715
rect -4710 4695 -4690 4715
rect -4670 4695 -4650 4715
rect -4630 4695 -4610 4715
rect -4590 4695 -4570 4715
rect -4550 4695 -4530 4715
rect -4510 4695 -4490 4715
rect -4470 4695 -4450 4715
rect -4430 4695 -4410 4715
rect -4390 4695 -4370 4715
rect -4350 4695 -4330 4715
rect -4310 4695 -4290 4715
rect -4270 4695 -4250 4715
rect -4230 4695 -4210 4715
rect -4190 4695 -4170 4715
rect -4150 4695 -4130 4715
rect -4110 4695 -4090 4715
rect -4070 4695 -4050 4715
rect -4030 4695 -4010 4715
rect -3990 4695 -3970 4715
rect -3950 4695 -3930 4715
rect -3910 4695 -3890 4715
rect -3870 4695 -3850 4715
rect -3830 4695 -3810 4715
rect -3790 4695 -3770 4715
rect -3750 4695 -3730 4715
rect -3710 4695 -3690 4715
rect -3670 4695 -3650 4715
rect -3630 4695 -3610 4715
rect -3590 4695 -3570 4715
rect -3550 4695 -3530 4715
rect -3510 4695 -3490 4715
rect -3470 4695 -3450 4715
rect -3430 4695 -3410 4715
rect -3390 4695 -3370 4715
rect -3350 4695 -3330 4715
rect -3310 4695 -3290 4715
rect -3270 4695 -3250 4715
rect -3230 4695 -3210 4715
rect -3190 4695 -3170 4715
rect -3150 4695 -3130 4715
rect -3110 4695 -3095 4715
rect -5595 4680 -3095 4695
rect -2045 4715 455 4730
rect -2045 4695 -2030 4715
rect -2010 4695 -1990 4715
rect -1970 4695 -1950 4715
rect -1930 4695 -1910 4715
rect -1890 4695 -1870 4715
rect -1850 4695 -1830 4715
rect -1810 4695 -1790 4715
rect -1770 4695 -1750 4715
rect -1730 4695 -1710 4715
rect -1690 4695 -1670 4715
rect -1650 4695 -1630 4715
rect -1610 4695 -1590 4715
rect -1570 4695 -1550 4715
rect -1530 4695 -1510 4715
rect -1490 4695 -1470 4715
rect -1450 4695 -1430 4715
rect -1410 4695 -1390 4715
rect -1370 4695 -1350 4715
rect -1330 4695 -1310 4715
rect -1290 4695 -1270 4715
rect -1250 4695 -1230 4715
rect -1210 4695 -1190 4715
rect -1170 4695 -1150 4715
rect -1130 4695 -1110 4715
rect -1090 4695 -1070 4715
rect -1050 4695 -1030 4715
rect -1010 4695 -990 4715
rect -970 4695 -950 4715
rect -930 4695 -910 4715
rect -890 4695 -870 4715
rect -850 4695 -830 4715
rect -810 4695 -790 4715
rect -770 4695 -750 4715
rect -730 4695 -710 4715
rect -690 4695 -670 4715
rect -650 4695 -630 4715
rect -610 4695 -590 4715
rect -570 4695 -550 4715
rect -530 4695 -510 4715
rect -490 4695 -470 4715
rect -450 4695 -430 4715
rect -410 4695 -390 4715
rect -370 4695 -350 4715
rect -330 4695 -310 4715
rect -290 4695 -270 4715
rect -250 4695 -230 4715
rect -210 4695 -190 4715
rect -170 4695 -150 4715
rect -130 4695 -110 4715
rect -90 4695 -70 4715
rect -50 4695 -30 4715
rect -10 4695 10 4715
rect 30 4695 50 4715
rect 70 4695 90 4715
rect 110 4695 130 4715
rect 150 4695 170 4715
rect 190 4695 210 4715
rect 230 4695 250 4715
rect 270 4695 290 4715
rect 310 4695 330 4715
rect 350 4695 370 4715
rect 390 4695 410 4715
rect 440 4695 455 4715
rect -2045 4680 455 4695
rect -5595 4620 -3095 4635
rect -5595 4600 -5580 4620
rect -5550 4600 -5530 4620
rect -5510 4600 -5490 4620
rect -5470 4600 -5450 4620
rect -5430 4600 -5410 4620
rect -5390 4600 -5370 4620
rect -5350 4600 -5330 4620
rect -5310 4600 -5290 4620
rect -5270 4600 -5250 4620
rect -5230 4600 -5210 4620
rect -5190 4600 -5170 4620
rect -5150 4600 -5130 4620
rect -5110 4600 -5090 4620
rect -5070 4600 -5050 4620
rect -5030 4600 -5010 4620
rect -4990 4600 -4970 4620
rect -4950 4600 -4930 4620
rect -4910 4600 -4890 4620
rect -4870 4600 -4850 4620
rect -4830 4600 -4810 4620
rect -4790 4600 -4770 4620
rect -4750 4600 -4730 4620
rect -4710 4600 -4690 4620
rect -4670 4600 -4650 4620
rect -4630 4600 -4610 4620
rect -4590 4600 -4570 4620
rect -4550 4600 -4530 4620
rect -4510 4600 -4490 4620
rect -4470 4600 -4450 4620
rect -4430 4600 -4410 4620
rect -4390 4600 -4370 4620
rect -4350 4600 -4330 4620
rect -4310 4600 -4290 4620
rect -4270 4600 -4250 4620
rect -4230 4600 -4210 4620
rect -4190 4600 -4170 4620
rect -4150 4600 -4130 4620
rect -4110 4600 -4090 4620
rect -4070 4600 -4050 4620
rect -4030 4600 -4010 4620
rect -3990 4600 -3970 4620
rect -3950 4600 -3930 4620
rect -3910 4600 -3890 4620
rect -3870 4600 -3850 4620
rect -3830 4600 -3810 4620
rect -3790 4600 -3770 4620
rect -3750 4600 -3730 4620
rect -3710 4600 -3690 4620
rect -3670 4600 -3650 4620
rect -3630 4600 -3610 4620
rect -3590 4600 -3570 4620
rect -3550 4600 -3530 4620
rect -3510 4600 -3490 4620
rect -3470 4600 -3450 4620
rect -3430 4600 -3410 4620
rect -3390 4600 -3370 4620
rect -3350 4600 -3330 4620
rect -3310 4600 -3290 4620
rect -3270 4600 -3250 4620
rect -3230 4600 -3210 4620
rect -3190 4600 -3170 4620
rect -3150 4600 -3130 4620
rect -3110 4600 -3095 4620
rect -5595 4585 -3095 4600
rect -2045 4620 455 4635
rect -2045 4600 -2030 4620
rect -2010 4600 -1990 4620
rect -1970 4600 -1950 4620
rect -1930 4600 -1910 4620
rect -1890 4600 -1870 4620
rect -1850 4600 -1830 4620
rect -1810 4600 -1790 4620
rect -1770 4600 -1750 4620
rect -1730 4600 -1710 4620
rect -1690 4600 -1670 4620
rect -1650 4600 -1630 4620
rect -1610 4600 -1590 4620
rect -1570 4600 -1550 4620
rect -1530 4600 -1510 4620
rect -1490 4600 -1470 4620
rect -1450 4600 -1430 4620
rect -1410 4600 -1390 4620
rect -1370 4600 -1350 4620
rect -1330 4600 -1310 4620
rect -1290 4600 -1270 4620
rect -1250 4600 -1230 4620
rect -1210 4600 -1190 4620
rect -1170 4600 -1150 4620
rect -1130 4600 -1110 4620
rect -1090 4600 -1070 4620
rect -1050 4600 -1030 4620
rect -1010 4600 -990 4620
rect -970 4600 -950 4620
rect -930 4600 -910 4620
rect -890 4600 -870 4620
rect -850 4600 -830 4620
rect -810 4600 -790 4620
rect -770 4600 -750 4620
rect -730 4600 -710 4620
rect -690 4600 -670 4620
rect -650 4600 -630 4620
rect -610 4600 -590 4620
rect -570 4600 -550 4620
rect -530 4600 -510 4620
rect -490 4600 -470 4620
rect -450 4600 -430 4620
rect -410 4600 -390 4620
rect -370 4600 -350 4620
rect -330 4600 -310 4620
rect -290 4600 -270 4620
rect -250 4600 -230 4620
rect -210 4600 -190 4620
rect -170 4600 -150 4620
rect -130 4600 -110 4620
rect -90 4600 -70 4620
rect -50 4600 -30 4620
rect -10 4600 10 4620
rect 30 4600 50 4620
rect 70 4600 90 4620
rect 110 4600 130 4620
rect 150 4600 170 4620
rect 190 4600 210 4620
rect 230 4600 250 4620
rect 270 4600 290 4620
rect 310 4600 330 4620
rect 350 4600 370 4620
rect 390 4600 410 4620
rect 440 4600 455 4620
rect -2045 4585 455 4600
rect -5595 4525 -3095 4540
rect -5595 4505 -5580 4525
rect -5550 4505 -5530 4525
rect -5510 4505 -5490 4525
rect -5470 4505 -5450 4525
rect -5430 4505 -5410 4525
rect -5390 4505 -5370 4525
rect -5350 4505 -5330 4525
rect -5310 4505 -5290 4525
rect -5270 4505 -5250 4525
rect -5230 4505 -5210 4525
rect -5190 4505 -5170 4525
rect -5150 4505 -5130 4525
rect -5110 4505 -5090 4525
rect -5070 4505 -5050 4525
rect -5030 4505 -5010 4525
rect -4990 4505 -4970 4525
rect -4950 4505 -4930 4525
rect -4910 4505 -4890 4525
rect -4870 4505 -4850 4525
rect -4830 4505 -4810 4525
rect -4790 4505 -4770 4525
rect -4750 4505 -4730 4525
rect -4710 4505 -4690 4525
rect -4670 4505 -4650 4525
rect -4630 4505 -4610 4525
rect -4590 4505 -4570 4525
rect -4550 4505 -4530 4525
rect -4510 4505 -4490 4525
rect -4470 4505 -4450 4525
rect -4430 4505 -4410 4525
rect -4390 4505 -4370 4525
rect -4350 4505 -4330 4525
rect -4310 4505 -4290 4525
rect -4270 4505 -4250 4525
rect -4230 4505 -4210 4525
rect -4190 4505 -4170 4525
rect -4150 4505 -4130 4525
rect -4110 4505 -4090 4525
rect -4070 4505 -4050 4525
rect -4030 4505 -4010 4525
rect -3990 4505 -3970 4525
rect -3950 4505 -3930 4525
rect -3910 4505 -3890 4525
rect -3870 4505 -3850 4525
rect -3830 4505 -3810 4525
rect -3790 4505 -3770 4525
rect -3750 4505 -3730 4525
rect -3710 4505 -3690 4525
rect -3670 4505 -3650 4525
rect -3630 4505 -3610 4525
rect -3590 4505 -3570 4525
rect -3550 4505 -3530 4525
rect -3510 4505 -3490 4525
rect -3470 4505 -3450 4525
rect -3430 4505 -3410 4525
rect -3390 4505 -3370 4525
rect -3350 4505 -3330 4525
rect -3310 4505 -3290 4525
rect -3270 4505 -3250 4525
rect -3230 4505 -3210 4525
rect -3190 4505 -3170 4525
rect -3150 4505 -3130 4525
rect -3110 4505 -3095 4525
rect -5595 4490 -3095 4505
rect -2045 4525 455 4540
rect -2045 4505 -2030 4525
rect -2010 4505 -1990 4525
rect -1970 4505 -1950 4525
rect -1930 4505 -1910 4525
rect -1890 4505 -1870 4525
rect -1850 4505 -1830 4525
rect -1810 4505 -1790 4525
rect -1770 4505 -1750 4525
rect -1730 4505 -1710 4525
rect -1690 4505 -1670 4525
rect -1650 4505 -1630 4525
rect -1610 4505 -1590 4525
rect -1570 4505 -1550 4525
rect -1530 4505 -1510 4525
rect -1490 4505 -1470 4525
rect -1450 4505 -1430 4525
rect -1410 4505 -1390 4525
rect -1370 4505 -1350 4525
rect -1330 4505 -1310 4525
rect -1290 4505 -1270 4525
rect -1250 4505 -1230 4525
rect -1210 4505 -1190 4525
rect -1170 4505 -1150 4525
rect -1130 4505 -1110 4525
rect -1090 4505 -1070 4525
rect -1050 4505 -1030 4525
rect -1010 4505 -990 4525
rect -970 4505 -950 4525
rect -930 4505 -910 4525
rect -890 4505 -870 4525
rect -850 4505 -830 4525
rect -810 4505 -790 4525
rect -770 4505 -750 4525
rect -730 4505 -710 4525
rect -690 4505 -670 4525
rect -650 4505 -630 4525
rect -610 4505 -590 4525
rect -570 4505 -550 4525
rect -530 4505 -510 4525
rect -490 4505 -470 4525
rect -450 4505 -430 4525
rect -410 4505 -390 4525
rect -370 4505 -350 4525
rect -330 4505 -310 4525
rect -290 4505 -270 4525
rect -250 4505 -230 4525
rect -210 4505 -190 4525
rect -170 4505 -150 4525
rect -130 4505 -110 4525
rect -90 4505 -70 4525
rect -50 4505 -30 4525
rect -10 4505 10 4525
rect 30 4505 50 4525
rect 70 4505 90 4525
rect 110 4505 130 4525
rect 150 4505 170 4525
rect 190 4505 210 4525
rect 230 4505 250 4525
rect 270 4505 290 4525
rect 310 4505 330 4525
rect 350 4505 370 4525
rect 390 4505 410 4525
rect 440 4505 455 4525
rect -2045 4490 455 4505
rect -5595 4430 -3095 4445
rect -5595 4410 -5580 4430
rect -5550 4410 -5530 4430
rect -5510 4410 -5490 4430
rect -5470 4410 -5450 4430
rect -5430 4410 -5410 4430
rect -5390 4410 -5370 4430
rect -5350 4410 -5330 4430
rect -5310 4410 -5290 4430
rect -5270 4410 -5250 4430
rect -5230 4410 -5210 4430
rect -5190 4410 -5170 4430
rect -5150 4410 -5130 4430
rect -5110 4410 -5090 4430
rect -5070 4410 -5050 4430
rect -5030 4410 -5010 4430
rect -4990 4410 -4970 4430
rect -4950 4410 -4930 4430
rect -4910 4410 -4890 4430
rect -4870 4410 -4850 4430
rect -4830 4410 -4810 4430
rect -4790 4410 -4770 4430
rect -4750 4410 -4730 4430
rect -4710 4410 -4690 4430
rect -4670 4410 -4650 4430
rect -4630 4410 -4610 4430
rect -4590 4410 -4570 4430
rect -4550 4410 -4530 4430
rect -4510 4410 -4490 4430
rect -4470 4410 -4450 4430
rect -4430 4410 -4410 4430
rect -4390 4410 -4370 4430
rect -4350 4410 -4330 4430
rect -4310 4410 -4290 4430
rect -4270 4410 -4250 4430
rect -4230 4410 -4210 4430
rect -4190 4410 -4170 4430
rect -4150 4410 -4130 4430
rect -4110 4410 -4090 4430
rect -4070 4410 -4050 4430
rect -4030 4410 -4010 4430
rect -3990 4410 -3970 4430
rect -3950 4410 -3930 4430
rect -3910 4410 -3890 4430
rect -3870 4410 -3850 4430
rect -3830 4410 -3810 4430
rect -3790 4410 -3770 4430
rect -3750 4410 -3730 4430
rect -3710 4410 -3690 4430
rect -3670 4410 -3650 4430
rect -3630 4410 -3610 4430
rect -3590 4410 -3570 4430
rect -3550 4410 -3530 4430
rect -3510 4410 -3490 4430
rect -3470 4410 -3450 4430
rect -3430 4410 -3410 4430
rect -3390 4410 -3370 4430
rect -3350 4410 -3330 4430
rect -3310 4410 -3290 4430
rect -3270 4410 -3250 4430
rect -3230 4410 -3210 4430
rect -3190 4410 -3170 4430
rect -3150 4410 -3130 4430
rect -3110 4410 -3095 4430
rect -5595 4395 -3095 4410
rect -2045 4430 455 4445
rect -2045 4410 -2030 4430
rect -2010 4410 -1990 4430
rect -1970 4410 -1950 4430
rect -1930 4410 -1910 4430
rect -1890 4410 -1870 4430
rect -1850 4410 -1830 4430
rect -1810 4410 -1790 4430
rect -1770 4410 -1750 4430
rect -1730 4410 -1710 4430
rect -1690 4410 -1670 4430
rect -1650 4410 -1630 4430
rect -1610 4410 -1590 4430
rect -1570 4410 -1550 4430
rect -1530 4410 -1510 4430
rect -1490 4410 -1470 4430
rect -1450 4410 -1430 4430
rect -1410 4410 -1390 4430
rect -1370 4410 -1350 4430
rect -1330 4410 -1310 4430
rect -1290 4410 -1270 4430
rect -1250 4410 -1230 4430
rect -1210 4410 -1190 4430
rect -1170 4410 -1150 4430
rect -1130 4410 -1110 4430
rect -1090 4410 -1070 4430
rect -1050 4410 -1030 4430
rect -1010 4410 -990 4430
rect -970 4410 -950 4430
rect -930 4410 -910 4430
rect -890 4410 -870 4430
rect -850 4410 -830 4430
rect -810 4410 -790 4430
rect -770 4410 -750 4430
rect -730 4410 -710 4430
rect -690 4410 -670 4430
rect -650 4410 -630 4430
rect -610 4410 -590 4430
rect -570 4410 -550 4430
rect -530 4410 -510 4430
rect -490 4410 -470 4430
rect -450 4410 -430 4430
rect -410 4410 -390 4430
rect -370 4410 -350 4430
rect -330 4410 -310 4430
rect -290 4410 -270 4430
rect -250 4410 -230 4430
rect -210 4410 -190 4430
rect -170 4410 -150 4430
rect -130 4410 -110 4430
rect -90 4410 -70 4430
rect -50 4410 -30 4430
rect -10 4410 10 4430
rect 30 4410 50 4430
rect 70 4410 90 4430
rect 110 4410 130 4430
rect 150 4410 170 4430
rect 190 4410 210 4430
rect 230 4410 250 4430
rect 270 4410 290 4430
rect 310 4410 330 4430
rect 350 4410 370 4430
rect 390 4410 410 4430
rect 440 4410 455 4430
rect -2045 4395 455 4410
rect -5595 4335 -3095 4350
rect -5595 4315 -5580 4335
rect -5550 4315 -5530 4335
rect -5510 4315 -5490 4335
rect -5470 4315 -5450 4335
rect -5430 4315 -5410 4335
rect -5390 4315 -5370 4335
rect -5350 4315 -5330 4335
rect -5310 4315 -5290 4335
rect -5270 4315 -5250 4335
rect -5230 4315 -5210 4335
rect -5190 4315 -5170 4335
rect -5150 4315 -5130 4335
rect -5110 4315 -5090 4335
rect -5070 4315 -5050 4335
rect -5030 4315 -5010 4335
rect -4990 4315 -4970 4335
rect -4950 4315 -4930 4335
rect -4910 4315 -4890 4335
rect -4870 4315 -4850 4335
rect -4830 4315 -4810 4335
rect -4790 4315 -4770 4335
rect -4750 4315 -4730 4335
rect -4710 4315 -4690 4335
rect -4670 4315 -4650 4335
rect -4630 4315 -4610 4335
rect -4590 4315 -4570 4335
rect -4550 4315 -4530 4335
rect -4510 4315 -4490 4335
rect -4470 4315 -4450 4335
rect -4430 4315 -4410 4335
rect -4390 4315 -4370 4335
rect -4350 4315 -4330 4335
rect -4310 4315 -4290 4335
rect -4270 4315 -4250 4335
rect -4230 4315 -4210 4335
rect -4190 4315 -4170 4335
rect -4150 4315 -4130 4335
rect -4110 4315 -4090 4335
rect -4070 4315 -4050 4335
rect -4030 4315 -4010 4335
rect -3990 4315 -3970 4335
rect -3950 4315 -3930 4335
rect -3910 4315 -3890 4335
rect -3870 4315 -3850 4335
rect -3830 4315 -3810 4335
rect -3790 4315 -3770 4335
rect -3750 4315 -3730 4335
rect -3710 4315 -3690 4335
rect -3670 4315 -3650 4335
rect -3630 4315 -3610 4335
rect -3590 4315 -3570 4335
rect -3550 4315 -3530 4335
rect -3510 4315 -3490 4335
rect -3470 4315 -3450 4335
rect -3430 4315 -3410 4335
rect -3390 4315 -3370 4335
rect -3350 4315 -3330 4335
rect -3310 4315 -3290 4335
rect -3270 4315 -3250 4335
rect -3230 4315 -3210 4335
rect -3190 4315 -3170 4335
rect -3150 4315 -3130 4335
rect -3110 4315 -3095 4335
rect -5595 4300 -3095 4315
rect -2045 4335 455 4350
rect -2045 4315 -2030 4335
rect -2010 4315 -1990 4335
rect -1970 4315 -1950 4335
rect -1930 4315 -1910 4335
rect -1890 4315 -1870 4335
rect -1850 4315 -1830 4335
rect -1810 4315 -1790 4335
rect -1770 4315 -1750 4335
rect -1730 4315 -1710 4335
rect -1690 4315 -1670 4335
rect -1650 4315 -1630 4335
rect -1610 4315 -1590 4335
rect -1570 4315 -1550 4335
rect -1530 4315 -1510 4335
rect -1490 4315 -1470 4335
rect -1450 4315 -1430 4335
rect -1410 4315 -1390 4335
rect -1370 4315 -1350 4335
rect -1330 4315 -1310 4335
rect -1290 4315 -1270 4335
rect -1250 4315 -1230 4335
rect -1210 4315 -1190 4335
rect -1170 4315 -1150 4335
rect -1130 4315 -1110 4335
rect -1090 4315 -1070 4335
rect -1050 4315 -1030 4335
rect -1010 4315 -990 4335
rect -970 4315 -950 4335
rect -930 4315 -910 4335
rect -890 4315 -870 4335
rect -850 4315 -830 4335
rect -810 4315 -790 4335
rect -770 4315 -750 4335
rect -730 4315 -710 4335
rect -690 4315 -670 4335
rect -650 4315 -630 4335
rect -610 4315 -590 4335
rect -570 4315 -550 4335
rect -530 4315 -510 4335
rect -490 4315 -470 4335
rect -450 4315 -430 4335
rect -410 4315 -390 4335
rect -370 4315 -350 4335
rect -330 4315 -310 4335
rect -290 4315 -270 4335
rect -250 4315 -230 4335
rect -210 4315 -190 4335
rect -170 4315 -150 4335
rect -130 4315 -110 4335
rect -90 4315 -70 4335
rect -50 4315 -30 4335
rect -10 4315 10 4335
rect 30 4315 50 4335
rect 70 4315 90 4335
rect 110 4315 130 4335
rect 150 4315 170 4335
rect 190 4315 210 4335
rect 230 4315 250 4335
rect 270 4315 290 4335
rect 310 4315 330 4335
rect 350 4315 370 4335
rect 390 4315 410 4335
rect 440 4315 455 4335
rect -2045 4300 455 4315
rect -5595 4240 -3095 4255
rect -5595 4220 -5580 4240
rect -5550 4220 -5530 4240
rect -5510 4220 -5490 4240
rect -5470 4220 -5450 4240
rect -5430 4220 -5410 4240
rect -5390 4220 -5370 4240
rect -5350 4220 -5330 4240
rect -5310 4220 -5290 4240
rect -5270 4220 -5250 4240
rect -5230 4220 -5210 4240
rect -5190 4220 -5170 4240
rect -5150 4220 -5130 4240
rect -5110 4220 -5090 4240
rect -5070 4220 -5050 4240
rect -5030 4220 -5010 4240
rect -4990 4220 -4970 4240
rect -4950 4220 -4930 4240
rect -4910 4220 -4890 4240
rect -4870 4220 -4850 4240
rect -4830 4220 -4810 4240
rect -4790 4220 -4770 4240
rect -4750 4220 -4730 4240
rect -4710 4220 -4690 4240
rect -4670 4220 -4650 4240
rect -4630 4220 -4610 4240
rect -4590 4220 -4570 4240
rect -4550 4220 -4530 4240
rect -4510 4220 -4490 4240
rect -4470 4220 -4450 4240
rect -4430 4220 -4410 4240
rect -4390 4220 -4370 4240
rect -4350 4220 -4330 4240
rect -4310 4220 -4290 4240
rect -4270 4220 -4250 4240
rect -4230 4220 -4210 4240
rect -4190 4220 -4170 4240
rect -4150 4220 -4130 4240
rect -4110 4220 -4090 4240
rect -4070 4220 -4050 4240
rect -4030 4220 -4010 4240
rect -3990 4220 -3970 4240
rect -3950 4220 -3930 4240
rect -3910 4220 -3890 4240
rect -3870 4220 -3850 4240
rect -3830 4220 -3810 4240
rect -3790 4220 -3770 4240
rect -3750 4220 -3730 4240
rect -3710 4220 -3690 4240
rect -3670 4220 -3650 4240
rect -3630 4220 -3610 4240
rect -3590 4220 -3570 4240
rect -3550 4220 -3530 4240
rect -3510 4220 -3490 4240
rect -3470 4220 -3450 4240
rect -3430 4220 -3410 4240
rect -3390 4220 -3370 4240
rect -3350 4220 -3330 4240
rect -3310 4220 -3290 4240
rect -3270 4220 -3250 4240
rect -3230 4220 -3210 4240
rect -3190 4220 -3170 4240
rect -3150 4220 -3130 4240
rect -3110 4220 -3095 4240
rect -5595 4205 -3095 4220
rect -2045 4240 455 4255
rect -2045 4220 -2030 4240
rect -2010 4220 -1990 4240
rect -1970 4220 -1950 4240
rect -1930 4220 -1910 4240
rect -1890 4220 -1870 4240
rect -1850 4220 -1830 4240
rect -1810 4220 -1790 4240
rect -1770 4220 -1750 4240
rect -1730 4220 -1710 4240
rect -1690 4220 -1670 4240
rect -1650 4220 -1630 4240
rect -1610 4220 -1590 4240
rect -1570 4220 -1550 4240
rect -1530 4220 -1510 4240
rect -1490 4220 -1470 4240
rect -1450 4220 -1430 4240
rect -1410 4220 -1390 4240
rect -1370 4220 -1350 4240
rect -1330 4220 -1310 4240
rect -1290 4220 -1270 4240
rect -1250 4220 -1230 4240
rect -1210 4220 -1190 4240
rect -1170 4220 -1150 4240
rect -1130 4220 -1110 4240
rect -1090 4220 -1070 4240
rect -1050 4220 -1030 4240
rect -1010 4220 -990 4240
rect -970 4220 -950 4240
rect -930 4220 -910 4240
rect -890 4220 -870 4240
rect -850 4220 -830 4240
rect -810 4220 -790 4240
rect -770 4220 -750 4240
rect -730 4220 -710 4240
rect -690 4220 -670 4240
rect -650 4220 -630 4240
rect -610 4220 -590 4240
rect -570 4220 -550 4240
rect -530 4220 -510 4240
rect -490 4220 -470 4240
rect -450 4220 -430 4240
rect -410 4220 -390 4240
rect -370 4220 -350 4240
rect -330 4220 -310 4240
rect -290 4220 -270 4240
rect -250 4220 -230 4240
rect -210 4220 -190 4240
rect -170 4220 -150 4240
rect -130 4220 -110 4240
rect -90 4220 -70 4240
rect -50 4220 -30 4240
rect -10 4220 10 4240
rect 30 4220 50 4240
rect 70 4220 90 4240
rect 110 4220 130 4240
rect 150 4220 170 4240
rect 190 4220 210 4240
rect 230 4220 250 4240
rect 270 4220 290 4240
rect 310 4220 330 4240
rect 350 4220 370 4240
rect 390 4220 410 4240
rect 440 4220 455 4240
rect -2045 4205 455 4220
rect -5595 4145 -3095 4160
rect -5595 4125 -5580 4145
rect -5550 4125 -5530 4145
rect -5510 4125 -5490 4145
rect -5470 4125 -5450 4145
rect -5430 4125 -5410 4145
rect -5390 4125 -5370 4145
rect -5350 4125 -5330 4145
rect -5310 4125 -5290 4145
rect -5270 4125 -5250 4145
rect -5230 4125 -5210 4145
rect -5190 4125 -5170 4145
rect -5150 4125 -5130 4145
rect -5110 4125 -5090 4145
rect -5070 4125 -5050 4145
rect -5030 4125 -5010 4145
rect -4990 4125 -4970 4145
rect -4950 4125 -4930 4145
rect -4910 4125 -4890 4145
rect -4870 4125 -4850 4145
rect -4830 4125 -4810 4145
rect -4790 4125 -4770 4145
rect -4750 4125 -4730 4145
rect -4710 4125 -4690 4145
rect -4670 4125 -4650 4145
rect -4630 4125 -4610 4145
rect -4590 4125 -4570 4145
rect -4550 4125 -4530 4145
rect -4510 4125 -4490 4145
rect -4470 4125 -4450 4145
rect -4430 4125 -4410 4145
rect -4390 4125 -4370 4145
rect -4350 4125 -4330 4145
rect -4310 4125 -4290 4145
rect -4270 4125 -4250 4145
rect -4230 4125 -4210 4145
rect -4190 4125 -4170 4145
rect -4150 4125 -4130 4145
rect -4110 4125 -4090 4145
rect -4070 4125 -4050 4145
rect -4030 4125 -4010 4145
rect -3990 4125 -3970 4145
rect -3950 4125 -3930 4145
rect -3910 4125 -3890 4145
rect -3870 4125 -3850 4145
rect -3830 4125 -3810 4145
rect -3790 4125 -3770 4145
rect -3750 4125 -3730 4145
rect -3710 4125 -3690 4145
rect -3670 4125 -3650 4145
rect -3630 4125 -3610 4145
rect -3590 4125 -3570 4145
rect -3550 4125 -3530 4145
rect -3510 4125 -3490 4145
rect -3470 4125 -3450 4145
rect -3430 4125 -3410 4145
rect -3390 4125 -3370 4145
rect -3350 4125 -3330 4145
rect -3310 4125 -3290 4145
rect -3270 4125 -3250 4145
rect -3230 4125 -3210 4145
rect -3190 4125 -3170 4145
rect -3150 4125 -3130 4145
rect -3110 4125 -3095 4145
rect -5595 4110 -3095 4125
rect -2045 4145 455 4160
rect -2045 4125 -2030 4145
rect -2010 4125 -1990 4145
rect -1970 4125 -1950 4145
rect -1930 4125 -1910 4145
rect -1890 4125 -1870 4145
rect -1850 4125 -1830 4145
rect -1810 4125 -1790 4145
rect -1770 4125 -1750 4145
rect -1730 4125 -1710 4145
rect -1690 4125 -1670 4145
rect -1650 4125 -1630 4145
rect -1610 4125 -1590 4145
rect -1570 4125 -1550 4145
rect -1530 4125 -1510 4145
rect -1490 4125 -1470 4145
rect -1450 4125 -1430 4145
rect -1410 4125 -1390 4145
rect -1370 4125 -1350 4145
rect -1330 4125 -1310 4145
rect -1290 4125 -1270 4145
rect -1250 4125 -1230 4145
rect -1210 4125 -1190 4145
rect -1170 4125 -1150 4145
rect -1130 4125 -1110 4145
rect -1090 4125 -1070 4145
rect -1050 4125 -1030 4145
rect -1010 4125 -990 4145
rect -970 4125 -950 4145
rect -930 4125 -910 4145
rect -890 4125 -870 4145
rect -850 4125 -830 4145
rect -810 4125 -790 4145
rect -770 4125 -750 4145
rect -730 4125 -710 4145
rect -690 4125 -670 4145
rect -650 4125 -630 4145
rect -610 4125 -590 4145
rect -570 4125 -550 4145
rect -530 4125 -510 4145
rect -490 4125 -470 4145
rect -450 4125 -430 4145
rect -410 4125 -390 4145
rect -370 4125 -350 4145
rect -330 4125 -310 4145
rect -290 4125 -270 4145
rect -250 4125 -230 4145
rect -210 4125 -190 4145
rect -170 4125 -150 4145
rect -130 4125 -110 4145
rect -90 4125 -70 4145
rect -50 4125 -30 4145
rect -10 4125 10 4145
rect 30 4125 50 4145
rect 70 4125 90 4145
rect 110 4125 130 4145
rect 150 4125 170 4145
rect 190 4125 210 4145
rect 230 4125 250 4145
rect 270 4125 290 4145
rect 310 4125 330 4145
rect 350 4125 370 4145
rect 390 4125 410 4145
rect 440 4125 455 4145
rect -2045 4110 455 4125
rect -5595 4050 -3095 4065
rect -5595 4030 -5580 4050
rect -5550 4030 -5530 4050
rect -5510 4030 -5490 4050
rect -5470 4030 -5450 4050
rect -5430 4030 -5410 4050
rect -5390 4030 -5370 4050
rect -5350 4030 -5330 4050
rect -5310 4030 -5290 4050
rect -5270 4030 -5250 4050
rect -5230 4030 -5210 4050
rect -5190 4030 -5170 4050
rect -5150 4030 -5130 4050
rect -5110 4030 -5090 4050
rect -5070 4030 -5050 4050
rect -5030 4030 -5010 4050
rect -4990 4030 -4970 4050
rect -4950 4030 -4930 4050
rect -4910 4030 -4890 4050
rect -4870 4030 -4850 4050
rect -4830 4030 -4810 4050
rect -4790 4030 -4770 4050
rect -4750 4030 -4730 4050
rect -4710 4030 -4690 4050
rect -4670 4030 -4650 4050
rect -4630 4030 -4610 4050
rect -4590 4030 -4570 4050
rect -4550 4030 -4530 4050
rect -4510 4030 -4490 4050
rect -4470 4030 -4450 4050
rect -4430 4030 -4410 4050
rect -4390 4030 -4370 4050
rect -4350 4030 -4330 4050
rect -4310 4030 -4290 4050
rect -4270 4030 -4250 4050
rect -4230 4030 -4210 4050
rect -4190 4030 -4170 4050
rect -4150 4030 -4130 4050
rect -4110 4030 -4090 4050
rect -4070 4030 -4050 4050
rect -4030 4030 -4010 4050
rect -3990 4030 -3970 4050
rect -3950 4030 -3930 4050
rect -3910 4030 -3890 4050
rect -3870 4030 -3850 4050
rect -3830 4030 -3810 4050
rect -3790 4030 -3770 4050
rect -3750 4030 -3730 4050
rect -3710 4030 -3690 4050
rect -3670 4030 -3650 4050
rect -3630 4030 -3610 4050
rect -3590 4030 -3570 4050
rect -3550 4030 -3530 4050
rect -3510 4030 -3490 4050
rect -3470 4030 -3450 4050
rect -3430 4030 -3410 4050
rect -3390 4030 -3370 4050
rect -3350 4030 -3330 4050
rect -3310 4030 -3290 4050
rect -3270 4030 -3250 4050
rect -3230 4030 -3210 4050
rect -3190 4030 -3170 4050
rect -3150 4030 -3130 4050
rect -3110 4030 -3095 4050
rect -5595 4015 -3095 4030
rect -2045 4050 455 4065
rect -2045 4030 -2030 4050
rect -2010 4030 -1990 4050
rect -1970 4030 -1950 4050
rect -1930 4030 -1910 4050
rect -1890 4030 -1870 4050
rect -1850 4030 -1830 4050
rect -1810 4030 -1790 4050
rect -1770 4030 -1750 4050
rect -1730 4030 -1710 4050
rect -1690 4030 -1670 4050
rect -1650 4030 -1630 4050
rect -1610 4030 -1590 4050
rect -1570 4030 -1550 4050
rect -1530 4030 -1510 4050
rect -1490 4030 -1470 4050
rect -1450 4030 -1430 4050
rect -1410 4030 -1390 4050
rect -1370 4030 -1350 4050
rect -1330 4030 -1310 4050
rect -1290 4030 -1270 4050
rect -1250 4030 -1230 4050
rect -1210 4030 -1190 4050
rect -1170 4030 -1150 4050
rect -1130 4030 -1110 4050
rect -1090 4030 -1070 4050
rect -1050 4030 -1030 4050
rect -1010 4030 -990 4050
rect -970 4030 -950 4050
rect -930 4030 -910 4050
rect -890 4030 -870 4050
rect -850 4030 -830 4050
rect -810 4030 -790 4050
rect -770 4030 -750 4050
rect -730 4030 -710 4050
rect -690 4030 -670 4050
rect -650 4030 -630 4050
rect -610 4030 -590 4050
rect -570 4030 -550 4050
rect -530 4030 -510 4050
rect -490 4030 -470 4050
rect -450 4030 -430 4050
rect -410 4030 -390 4050
rect -370 4030 -350 4050
rect -330 4030 -310 4050
rect -290 4030 -270 4050
rect -250 4030 -230 4050
rect -210 4030 -190 4050
rect -170 4030 -150 4050
rect -130 4030 -110 4050
rect -90 4030 -70 4050
rect -50 4030 -30 4050
rect -10 4030 10 4050
rect 30 4030 50 4050
rect 70 4030 90 4050
rect 110 4030 130 4050
rect 150 4030 170 4050
rect 190 4030 210 4050
rect 230 4030 250 4050
rect 270 4030 290 4050
rect 310 4030 330 4050
rect 350 4030 370 4050
rect 390 4030 410 4050
rect 440 4030 455 4050
rect -2045 4015 455 4030
rect -5595 3955 -3095 3970
rect -5595 3935 -5580 3955
rect -5550 3935 -5530 3955
rect -5510 3935 -5490 3955
rect -5470 3935 -5450 3955
rect -5430 3935 -5410 3955
rect -5390 3935 -5370 3955
rect -5350 3935 -5330 3955
rect -5310 3935 -5290 3955
rect -5270 3935 -5250 3955
rect -5230 3935 -5210 3955
rect -5190 3935 -5170 3955
rect -5150 3935 -5130 3955
rect -5110 3935 -5090 3955
rect -5070 3935 -5050 3955
rect -5030 3935 -5010 3955
rect -4990 3935 -4970 3955
rect -4950 3935 -4930 3955
rect -4910 3935 -4890 3955
rect -4870 3935 -4850 3955
rect -4830 3935 -4810 3955
rect -4790 3935 -4770 3955
rect -4750 3935 -4730 3955
rect -4710 3935 -4690 3955
rect -4670 3935 -4650 3955
rect -4630 3935 -4610 3955
rect -4590 3935 -4570 3955
rect -4550 3935 -4530 3955
rect -4510 3935 -4490 3955
rect -4470 3935 -4450 3955
rect -4430 3935 -4410 3955
rect -4390 3935 -4370 3955
rect -4350 3935 -4330 3955
rect -4310 3935 -4290 3955
rect -4270 3935 -4250 3955
rect -4230 3935 -4210 3955
rect -4190 3935 -4170 3955
rect -4150 3935 -4130 3955
rect -4110 3935 -4090 3955
rect -4070 3935 -4050 3955
rect -4030 3935 -4010 3955
rect -3990 3935 -3970 3955
rect -3950 3935 -3930 3955
rect -3910 3935 -3890 3955
rect -3870 3935 -3850 3955
rect -3830 3935 -3810 3955
rect -3790 3935 -3770 3955
rect -3750 3935 -3730 3955
rect -3710 3935 -3690 3955
rect -3670 3935 -3650 3955
rect -3630 3935 -3610 3955
rect -3590 3935 -3570 3955
rect -3550 3935 -3530 3955
rect -3510 3935 -3490 3955
rect -3470 3935 -3450 3955
rect -3430 3935 -3410 3955
rect -3390 3935 -3370 3955
rect -3350 3935 -3330 3955
rect -3310 3935 -3290 3955
rect -3270 3935 -3250 3955
rect -3230 3935 -3210 3955
rect -3190 3935 -3170 3955
rect -3150 3935 -3130 3955
rect -3110 3935 -3095 3955
rect -5595 3920 -3095 3935
rect -2045 3955 455 3970
rect -2045 3935 -2030 3955
rect -2010 3935 -1990 3955
rect -1970 3935 -1950 3955
rect -1930 3935 -1910 3955
rect -1890 3935 -1870 3955
rect -1850 3935 -1830 3955
rect -1810 3935 -1790 3955
rect -1770 3935 -1750 3955
rect -1730 3935 -1710 3955
rect -1690 3935 -1670 3955
rect -1650 3935 -1630 3955
rect -1610 3935 -1590 3955
rect -1570 3935 -1550 3955
rect -1530 3935 -1510 3955
rect -1490 3935 -1470 3955
rect -1450 3935 -1430 3955
rect -1410 3935 -1390 3955
rect -1370 3935 -1350 3955
rect -1330 3935 -1310 3955
rect -1290 3935 -1270 3955
rect -1250 3935 -1230 3955
rect -1210 3935 -1190 3955
rect -1170 3935 -1150 3955
rect -1130 3935 -1110 3955
rect -1090 3935 -1070 3955
rect -1050 3935 -1030 3955
rect -1010 3935 -990 3955
rect -970 3935 -950 3955
rect -930 3935 -910 3955
rect -890 3935 -870 3955
rect -850 3935 -830 3955
rect -810 3935 -790 3955
rect -770 3935 -750 3955
rect -730 3935 -710 3955
rect -690 3935 -670 3955
rect -650 3935 -630 3955
rect -610 3935 -590 3955
rect -570 3935 -550 3955
rect -530 3935 -510 3955
rect -490 3935 -470 3955
rect -450 3935 -430 3955
rect -410 3935 -390 3955
rect -370 3935 -350 3955
rect -330 3935 -310 3955
rect -290 3935 -270 3955
rect -250 3935 -230 3955
rect -210 3935 -190 3955
rect -170 3935 -150 3955
rect -130 3935 -110 3955
rect -90 3935 -70 3955
rect -50 3935 -30 3955
rect -10 3935 10 3955
rect 30 3935 50 3955
rect 70 3935 90 3955
rect 110 3935 130 3955
rect 150 3935 170 3955
rect 190 3935 210 3955
rect 230 3935 250 3955
rect 270 3935 290 3955
rect 310 3935 330 3955
rect 350 3935 370 3955
rect 390 3935 410 3955
rect 440 3935 455 3955
rect -2045 3920 455 3935
rect -5595 3860 -3095 3875
rect -5595 3840 -5580 3860
rect -5550 3840 -5530 3860
rect -5510 3840 -5490 3860
rect -5470 3840 -5450 3860
rect -5430 3840 -5410 3860
rect -5390 3840 -5370 3860
rect -5350 3840 -5330 3860
rect -5310 3840 -5290 3860
rect -5270 3840 -5250 3860
rect -5230 3840 -5210 3860
rect -5190 3840 -5170 3860
rect -5150 3840 -5130 3860
rect -5110 3840 -5090 3860
rect -5070 3840 -5050 3860
rect -5030 3840 -5010 3860
rect -4990 3840 -4970 3860
rect -4950 3840 -4930 3860
rect -4910 3840 -4890 3860
rect -4870 3840 -4850 3860
rect -4830 3840 -4810 3860
rect -4790 3840 -4770 3860
rect -4750 3840 -4730 3860
rect -4710 3840 -4690 3860
rect -4670 3840 -4650 3860
rect -4630 3840 -4610 3860
rect -4590 3840 -4570 3860
rect -4550 3840 -4530 3860
rect -4510 3840 -4490 3860
rect -4470 3840 -4450 3860
rect -4430 3840 -4410 3860
rect -4390 3840 -4370 3860
rect -4350 3840 -4330 3860
rect -4310 3840 -4290 3860
rect -4270 3840 -4250 3860
rect -4230 3840 -4210 3860
rect -4190 3840 -4170 3860
rect -4150 3840 -4130 3860
rect -4110 3840 -4090 3860
rect -4070 3840 -4050 3860
rect -4030 3840 -4010 3860
rect -3990 3840 -3970 3860
rect -3950 3840 -3930 3860
rect -3910 3840 -3890 3860
rect -3870 3840 -3850 3860
rect -3830 3840 -3810 3860
rect -3790 3840 -3770 3860
rect -3750 3840 -3730 3860
rect -3710 3840 -3690 3860
rect -3670 3840 -3650 3860
rect -3630 3840 -3610 3860
rect -3590 3840 -3570 3860
rect -3550 3840 -3530 3860
rect -3510 3840 -3490 3860
rect -3470 3840 -3450 3860
rect -3430 3840 -3410 3860
rect -3390 3840 -3370 3860
rect -3350 3840 -3330 3860
rect -3310 3840 -3290 3860
rect -3270 3840 -3250 3860
rect -3230 3840 -3210 3860
rect -3190 3840 -3170 3860
rect -3150 3840 -3130 3860
rect -3110 3840 -3095 3860
rect -5595 3825 -3095 3840
rect -2045 3860 455 3875
rect -2045 3840 -2030 3860
rect -2010 3840 -1990 3860
rect -1970 3840 -1950 3860
rect -1930 3840 -1910 3860
rect -1890 3840 -1870 3860
rect -1850 3840 -1830 3860
rect -1810 3840 -1790 3860
rect -1770 3840 -1750 3860
rect -1730 3840 -1710 3860
rect -1690 3840 -1670 3860
rect -1650 3840 -1630 3860
rect -1610 3840 -1590 3860
rect -1570 3840 -1550 3860
rect -1530 3840 -1510 3860
rect -1490 3840 -1470 3860
rect -1450 3840 -1430 3860
rect -1410 3840 -1390 3860
rect -1370 3840 -1350 3860
rect -1330 3840 -1310 3860
rect -1290 3840 -1270 3860
rect -1250 3840 -1230 3860
rect -1210 3840 -1190 3860
rect -1170 3840 -1150 3860
rect -1130 3840 -1110 3860
rect -1090 3840 -1070 3860
rect -1050 3840 -1030 3860
rect -1010 3840 -990 3860
rect -970 3840 -950 3860
rect -930 3840 -910 3860
rect -890 3840 -870 3860
rect -850 3840 -830 3860
rect -810 3840 -790 3860
rect -770 3840 -750 3860
rect -730 3840 -710 3860
rect -690 3840 -670 3860
rect -650 3840 -630 3860
rect -610 3840 -590 3860
rect -570 3840 -550 3860
rect -530 3840 -510 3860
rect -490 3840 -470 3860
rect -450 3840 -430 3860
rect -410 3840 -390 3860
rect -370 3840 -350 3860
rect -330 3840 -310 3860
rect -290 3840 -270 3860
rect -250 3840 -230 3860
rect -210 3840 -190 3860
rect -170 3840 -150 3860
rect -130 3840 -110 3860
rect -90 3840 -70 3860
rect -50 3840 -30 3860
rect -10 3840 10 3860
rect 30 3840 50 3860
rect 70 3840 90 3860
rect 110 3840 130 3860
rect 150 3840 170 3860
rect 190 3840 210 3860
rect 230 3840 250 3860
rect 270 3840 290 3860
rect 310 3840 330 3860
rect 350 3840 370 3860
rect 390 3840 410 3860
rect 440 3840 455 3860
rect -2045 3825 455 3840
rect -5595 3765 -3095 3780
rect -5595 3745 -5580 3765
rect -5550 3745 -5530 3765
rect -5510 3745 -5490 3765
rect -5470 3745 -5450 3765
rect -5430 3745 -5410 3765
rect -5390 3745 -5370 3765
rect -5350 3745 -5330 3765
rect -5310 3745 -5290 3765
rect -5270 3745 -5250 3765
rect -5230 3745 -5210 3765
rect -5190 3745 -5170 3765
rect -5150 3745 -5130 3765
rect -5110 3745 -5090 3765
rect -5070 3745 -5050 3765
rect -5030 3745 -5010 3765
rect -4990 3745 -4970 3765
rect -4950 3745 -4930 3765
rect -4910 3745 -4890 3765
rect -4870 3745 -4850 3765
rect -4830 3745 -4810 3765
rect -4790 3745 -4770 3765
rect -4750 3745 -4730 3765
rect -4710 3745 -4690 3765
rect -4670 3745 -4650 3765
rect -4630 3745 -4610 3765
rect -4590 3745 -4570 3765
rect -4550 3745 -4530 3765
rect -4510 3745 -4490 3765
rect -4470 3745 -4450 3765
rect -4430 3745 -4410 3765
rect -4390 3745 -4370 3765
rect -4350 3745 -4330 3765
rect -4310 3745 -4290 3765
rect -4270 3745 -4250 3765
rect -4230 3745 -4210 3765
rect -4190 3745 -4170 3765
rect -4150 3745 -4130 3765
rect -4110 3745 -4090 3765
rect -4070 3745 -4050 3765
rect -4030 3745 -4010 3765
rect -3990 3745 -3970 3765
rect -3950 3745 -3930 3765
rect -3910 3745 -3890 3765
rect -3870 3745 -3850 3765
rect -3830 3745 -3810 3765
rect -3790 3745 -3770 3765
rect -3750 3745 -3730 3765
rect -3710 3745 -3690 3765
rect -3670 3745 -3650 3765
rect -3630 3745 -3610 3765
rect -3590 3745 -3570 3765
rect -3550 3745 -3530 3765
rect -3510 3745 -3490 3765
rect -3470 3745 -3450 3765
rect -3430 3745 -3410 3765
rect -3390 3745 -3370 3765
rect -3350 3745 -3330 3765
rect -3310 3745 -3290 3765
rect -3270 3745 -3250 3765
rect -3230 3745 -3210 3765
rect -3190 3745 -3170 3765
rect -3150 3745 -3130 3765
rect -3110 3745 -3095 3765
rect -5595 3730 -3095 3745
rect -2045 3765 455 3780
rect -2045 3745 -2030 3765
rect -2010 3745 -1990 3765
rect -1970 3745 -1950 3765
rect -1930 3745 -1910 3765
rect -1890 3745 -1870 3765
rect -1850 3745 -1830 3765
rect -1810 3745 -1790 3765
rect -1770 3745 -1750 3765
rect -1730 3745 -1710 3765
rect -1690 3745 -1670 3765
rect -1650 3745 -1630 3765
rect -1610 3745 -1590 3765
rect -1570 3745 -1550 3765
rect -1530 3745 -1510 3765
rect -1490 3745 -1470 3765
rect -1450 3745 -1430 3765
rect -1410 3745 -1390 3765
rect -1370 3745 -1350 3765
rect -1330 3745 -1310 3765
rect -1290 3745 -1270 3765
rect -1250 3745 -1230 3765
rect -1210 3745 -1190 3765
rect -1170 3745 -1150 3765
rect -1130 3745 -1110 3765
rect -1090 3745 -1070 3765
rect -1050 3745 -1030 3765
rect -1010 3745 -990 3765
rect -970 3745 -950 3765
rect -930 3745 -910 3765
rect -890 3745 -870 3765
rect -850 3745 -830 3765
rect -810 3745 -790 3765
rect -770 3745 -750 3765
rect -730 3745 -710 3765
rect -690 3745 -670 3765
rect -650 3745 -630 3765
rect -610 3745 -590 3765
rect -570 3745 -550 3765
rect -530 3745 -510 3765
rect -490 3745 -470 3765
rect -450 3745 -430 3765
rect -410 3745 -390 3765
rect -370 3745 -350 3765
rect -330 3745 -310 3765
rect -290 3745 -270 3765
rect -250 3745 -230 3765
rect -210 3745 -190 3765
rect -170 3745 -150 3765
rect -130 3745 -110 3765
rect -90 3745 -70 3765
rect -50 3745 -30 3765
rect -10 3745 10 3765
rect 30 3745 50 3765
rect 70 3745 90 3765
rect 110 3745 130 3765
rect 150 3745 170 3765
rect 190 3745 210 3765
rect 230 3745 250 3765
rect 270 3745 290 3765
rect 310 3745 330 3765
rect 350 3745 370 3765
rect 390 3745 410 3765
rect 440 3745 455 3765
rect -2045 3730 455 3745
rect -5595 3670 -3095 3685
rect -5595 3650 -5580 3670
rect -5550 3650 -5530 3670
rect -5510 3650 -5490 3670
rect -5470 3650 -5450 3670
rect -5430 3650 -5410 3670
rect -5390 3650 -5370 3670
rect -5350 3650 -5330 3670
rect -5310 3650 -5290 3670
rect -5270 3650 -5250 3670
rect -5230 3650 -5210 3670
rect -5190 3650 -5170 3670
rect -5150 3650 -5130 3670
rect -5110 3650 -5090 3670
rect -5070 3650 -5050 3670
rect -5030 3650 -5010 3670
rect -4990 3650 -4970 3670
rect -4950 3650 -4930 3670
rect -4910 3650 -4890 3670
rect -4870 3650 -4850 3670
rect -4830 3650 -4810 3670
rect -4790 3650 -4770 3670
rect -4750 3650 -4730 3670
rect -4710 3650 -4690 3670
rect -4670 3650 -4650 3670
rect -4630 3650 -4610 3670
rect -4590 3650 -4570 3670
rect -4550 3650 -4530 3670
rect -4510 3650 -4490 3670
rect -4470 3650 -4450 3670
rect -4430 3650 -4410 3670
rect -4390 3650 -4370 3670
rect -4350 3650 -4330 3670
rect -4310 3650 -4290 3670
rect -4270 3650 -4250 3670
rect -4230 3650 -4210 3670
rect -4190 3650 -4170 3670
rect -4150 3650 -4130 3670
rect -4110 3650 -4090 3670
rect -4070 3650 -4050 3670
rect -4030 3650 -4010 3670
rect -3990 3650 -3970 3670
rect -3950 3650 -3930 3670
rect -3910 3650 -3890 3670
rect -3870 3650 -3850 3670
rect -3830 3650 -3810 3670
rect -3790 3650 -3770 3670
rect -3750 3650 -3730 3670
rect -3710 3650 -3690 3670
rect -3670 3650 -3650 3670
rect -3630 3650 -3610 3670
rect -3590 3650 -3570 3670
rect -3550 3650 -3530 3670
rect -3510 3650 -3490 3670
rect -3470 3650 -3450 3670
rect -3430 3650 -3410 3670
rect -3390 3650 -3370 3670
rect -3350 3650 -3330 3670
rect -3310 3650 -3290 3670
rect -3270 3650 -3250 3670
rect -3230 3650 -3210 3670
rect -3190 3650 -3170 3670
rect -3150 3650 -3130 3670
rect -3110 3650 -3095 3670
rect -5595 3635 -3095 3650
rect -2045 3670 455 3685
rect -2045 3650 -2030 3670
rect -2010 3650 -1990 3670
rect -1970 3650 -1950 3670
rect -1930 3650 -1910 3670
rect -1890 3650 -1870 3670
rect -1850 3650 -1830 3670
rect -1810 3650 -1790 3670
rect -1770 3650 -1750 3670
rect -1730 3650 -1710 3670
rect -1690 3650 -1670 3670
rect -1650 3650 -1630 3670
rect -1610 3650 -1590 3670
rect -1570 3650 -1550 3670
rect -1530 3650 -1510 3670
rect -1490 3650 -1470 3670
rect -1450 3650 -1430 3670
rect -1410 3650 -1390 3670
rect -1370 3650 -1350 3670
rect -1330 3650 -1310 3670
rect -1290 3650 -1270 3670
rect -1250 3650 -1230 3670
rect -1210 3650 -1190 3670
rect -1170 3650 -1150 3670
rect -1130 3650 -1110 3670
rect -1090 3650 -1070 3670
rect -1050 3650 -1030 3670
rect -1010 3650 -990 3670
rect -970 3650 -950 3670
rect -930 3650 -910 3670
rect -890 3650 -870 3670
rect -850 3650 -830 3670
rect -810 3650 -790 3670
rect -770 3650 -750 3670
rect -730 3650 -710 3670
rect -690 3650 -670 3670
rect -650 3650 -630 3670
rect -610 3650 -590 3670
rect -570 3650 -550 3670
rect -530 3650 -510 3670
rect -490 3650 -470 3670
rect -450 3650 -430 3670
rect -410 3650 -390 3670
rect -370 3650 -350 3670
rect -330 3650 -310 3670
rect -290 3650 -270 3670
rect -250 3650 -230 3670
rect -210 3650 -190 3670
rect -170 3650 -150 3670
rect -130 3650 -110 3670
rect -90 3650 -70 3670
rect -50 3650 -30 3670
rect -10 3650 10 3670
rect 30 3650 50 3670
rect 70 3650 90 3670
rect 110 3650 130 3670
rect 150 3650 170 3670
rect 190 3650 210 3670
rect 230 3650 250 3670
rect 270 3650 290 3670
rect 310 3650 330 3670
rect 350 3650 370 3670
rect 390 3650 410 3670
rect 440 3650 455 3670
rect -2045 3635 455 3650
rect -5595 3575 -3095 3590
rect -5595 3555 -5580 3575
rect -5550 3555 -5530 3575
rect -5510 3555 -5490 3575
rect -5470 3555 -5450 3575
rect -5430 3555 -5410 3575
rect -5390 3555 -5370 3575
rect -5350 3555 -5330 3575
rect -5310 3555 -5290 3575
rect -5270 3555 -5250 3575
rect -5230 3555 -5210 3575
rect -5190 3555 -5170 3575
rect -5150 3555 -5130 3575
rect -5110 3555 -5090 3575
rect -5070 3555 -5050 3575
rect -5030 3555 -5010 3575
rect -4990 3555 -4970 3575
rect -4950 3555 -4930 3575
rect -4910 3555 -4890 3575
rect -4870 3555 -4850 3575
rect -4830 3555 -4810 3575
rect -4790 3555 -4770 3575
rect -4750 3555 -4730 3575
rect -4710 3555 -4690 3575
rect -4670 3555 -4650 3575
rect -4630 3555 -4610 3575
rect -4590 3555 -4570 3575
rect -4550 3555 -4530 3575
rect -4510 3555 -4490 3575
rect -4470 3555 -4450 3575
rect -4430 3555 -4410 3575
rect -4390 3555 -4370 3575
rect -4350 3555 -4330 3575
rect -4310 3555 -4290 3575
rect -4270 3555 -4250 3575
rect -4230 3555 -4210 3575
rect -4190 3555 -4170 3575
rect -4150 3555 -4130 3575
rect -4110 3555 -4090 3575
rect -4070 3555 -4050 3575
rect -4030 3555 -4010 3575
rect -3990 3555 -3970 3575
rect -3950 3555 -3930 3575
rect -3910 3555 -3890 3575
rect -3870 3555 -3850 3575
rect -3830 3555 -3810 3575
rect -3790 3555 -3770 3575
rect -3750 3555 -3730 3575
rect -3710 3555 -3690 3575
rect -3670 3555 -3650 3575
rect -3630 3555 -3610 3575
rect -3590 3555 -3570 3575
rect -3550 3555 -3530 3575
rect -3510 3555 -3490 3575
rect -3470 3555 -3450 3575
rect -3430 3555 -3410 3575
rect -3390 3555 -3370 3575
rect -3350 3555 -3330 3575
rect -3310 3555 -3290 3575
rect -3270 3555 -3250 3575
rect -3230 3555 -3210 3575
rect -3190 3555 -3170 3575
rect -3150 3555 -3130 3575
rect -3110 3555 -3095 3575
rect -5595 3545 -3095 3555
rect -2045 3575 455 3590
rect -2045 3555 -2030 3575
rect -2010 3555 -1990 3575
rect -1970 3555 -1950 3575
rect -1930 3555 -1910 3575
rect -1890 3555 -1870 3575
rect -1850 3555 -1830 3575
rect -1810 3555 -1790 3575
rect -1770 3555 -1750 3575
rect -1730 3555 -1710 3575
rect -1690 3555 -1670 3575
rect -1650 3555 -1630 3575
rect -1610 3555 -1590 3575
rect -1570 3555 -1550 3575
rect -1530 3555 -1510 3575
rect -1490 3555 -1470 3575
rect -1450 3555 -1430 3575
rect -1410 3555 -1390 3575
rect -1370 3555 -1350 3575
rect -1330 3555 -1310 3575
rect -1290 3555 -1270 3575
rect -1250 3555 -1230 3575
rect -1210 3555 -1190 3575
rect -1170 3555 -1150 3575
rect -1130 3555 -1110 3575
rect -1090 3555 -1070 3575
rect -1050 3555 -1030 3575
rect -1010 3555 -990 3575
rect -970 3555 -950 3575
rect -930 3555 -910 3575
rect -890 3555 -870 3575
rect -850 3555 -830 3575
rect -810 3555 -790 3575
rect -770 3555 -750 3575
rect -730 3555 -710 3575
rect -690 3555 -670 3575
rect -650 3555 -630 3575
rect -610 3555 -590 3575
rect -570 3555 -550 3575
rect -530 3555 -510 3575
rect -490 3555 -470 3575
rect -450 3555 -430 3575
rect -410 3555 -390 3575
rect -370 3555 -350 3575
rect -330 3555 -310 3575
rect -290 3555 -270 3575
rect -250 3555 -230 3575
rect -210 3555 -190 3575
rect -170 3555 -150 3575
rect -130 3555 -110 3575
rect -90 3555 -70 3575
rect -50 3555 -30 3575
rect -10 3555 10 3575
rect 30 3555 50 3575
rect 70 3555 90 3575
rect 110 3555 130 3575
rect 150 3555 170 3575
rect 190 3555 210 3575
rect 230 3555 250 3575
rect 270 3555 290 3575
rect 310 3555 330 3575
rect 350 3555 370 3575
rect 390 3555 410 3575
rect 440 3555 455 3575
rect -2045 3545 455 3555
<< ndiffc >>
rect -5650 8457 -5630 8477
rect -5610 8457 -5590 8477
rect -5570 8457 -5550 8477
rect -5530 8457 -5510 8477
rect -5490 8457 -5470 8477
rect -5450 8457 -5430 8477
rect -5410 8457 -5390 8477
rect -5370 8457 -5350 8477
rect -5330 8457 -5310 8477
rect -5290 8457 -5270 8477
rect -5250 8457 -5230 8477
rect -5210 8457 -5190 8477
rect -5170 8457 -5150 8477
rect -5130 8457 -5110 8477
rect -5090 8457 -5070 8477
rect -5050 8457 -5030 8477
rect -5010 8457 -4990 8477
rect -4970 8457 -4950 8477
rect -4930 8457 -4910 8477
rect -4890 8457 -4870 8477
rect -4850 8457 -4830 8477
rect -4810 8457 -4790 8477
rect -4770 8457 -4750 8477
rect -4730 8457 -4710 8477
rect -4690 8457 -4670 8477
rect -4650 8457 -4630 8477
rect -4610 8457 -4590 8477
rect -4570 8457 -4550 8477
rect -4530 8457 -4510 8477
rect -4490 8457 -4470 8477
rect -4450 8457 -4430 8477
rect -4410 8457 -4390 8477
rect -4370 8457 -4350 8477
rect -4330 8457 -4310 8477
rect -4290 8457 -4270 8477
rect -4250 8457 -4230 8477
rect -4210 8457 -4190 8477
rect -4170 8457 -4150 8477
rect -4130 8457 -4110 8477
rect -4090 8457 -4070 8477
rect -4050 8457 -4030 8477
rect -4010 8457 -3990 8477
rect -3970 8457 -3950 8477
rect -3930 8457 -3910 8477
rect -3890 8457 -3870 8477
rect -3850 8457 -3830 8477
rect -3810 8457 -3790 8477
rect -3770 8457 -3750 8477
rect -3730 8457 -3710 8477
rect -3690 8457 -3670 8477
rect -3650 8457 -3630 8477
rect -3610 8457 -3590 8477
rect -3570 8457 -3550 8477
rect -3530 8457 -3510 8477
rect -3490 8457 -3470 8477
rect -3450 8457 -3430 8477
rect -3410 8457 -3390 8477
rect -3370 8457 -3350 8477
rect -3330 8457 -3310 8477
rect -3290 8457 -3270 8477
rect -3250 8457 -3230 8477
rect -3210 8457 -3190 8477
rect -5650 8375 -5630 8395
rect -5610 8375 -5590 8395
rect -5570 8375 -5550 8395
rect -5530 8375 -5510 8395
rect -5490 8375 -5470 8395
rect -5450 8375 -5430 8395
rect -5410 8375 -5390 8395
rect -5370 8375 -5350 8395
rect -5330 8375 -5310 8395
rect -5290 8375 -5270 8395
rect -5250 8375 -5230 8395
rect -5210 8375 -5190 8395
rect -5170 8375 -5150 8395
rect -5130 8375 -5110 8395
rect -5090 8375 -5070 8395
rect -5050 8375 -5030 8395
rect -5010 8375 -4990 8395
rect -4970 8375 -4950 8395
rect -4930 8375 -4910 8395
rect -4890 8375 -4870 8395
rect -4850 8375 -4830 8395
rect -4810 8375 -4790 8395
rect -4770 8375 -4750 8395
rect -4730 8375 -4710 8395
rect -4690 8375 -4670 8395
rect -4650 8375 -4630 8395
rect -4610 8375 -4590 8395
rect -4570 8375 -4550 8395
rect -4530 8375 -4510 8395
rect -4490 8375 -4470 8395
rect -4450 8375 -4430 8395
rect -4410 8375 -4390 8395
rect -4370 8375 -4350 8395
rect -4330 8375 -4310 8395
rect -4290 8375 -4270 8395
rect -4250 8375 -4230 8395
rect -4210 8375 -4190 8395
rect -4170 8375 -4150 8395
rect -4130 8375 -4110 8395
rect -4090 8375 -4070 8395
rect -4050 8375 -4030 8395
rect -4010 8375 -3990 8395
rect -3970 8375 -3950 8395
rect -3930 8375 -3910 8395
rect -3890 8375 -3870 8395
rect -3850 8375 -3830 8395
rect -3810 8375 -3790 8395
rect -3770 8375 -3750 8395
rect -3730 8375 -3710 8395
rect -3690 8375 -3670 8395
rect -3650 8375 -3630 8395
rect -3610 8375 -3590 8395
rect -3570 8375 -3550 8395
rect -3530 8375 -3510 8395
rect -3490 8375 -3470 8395
rect -3450 8375 -3430 8395
rect -3410 8375 -3390 8395
rect -3370 8375 -3350 8395
rect -3330 8375 -3310 8395
rect -3290 8375 -3270 8395
rect -3250 8375 -3230 8395
rect -3210 8375 -3190 8395
rect -5650 8293 -5630 8313
rect -5610 8293 -5590 8313
rect -5570 8293 -5550 8313
rect -5530 8293 -5510 8313
rect -5490 8293 -5470 8313
rect -5450 8293 -5430 8313
rect -5410 8293 -5390 8313
rect -5370 8293 -5350 8313
rect -5330 8293 -5310 8313
rect -5290 8293 -5270 8313
rect -5250 8293 -5230 8313
rect -5210 8293 -5190 8313
rect -5170 8293 -5150 8313
rect -5130 8293 -5110 8313
rect -5090 8293 -5070 8313
rect -5050 8293 -5030 8313
rect -5010 8293 -4990 8313
rect -4970 8293 -4950 8313
rect -4930 8293 -4910 8313
rect -4890 8293 -4870 8313
rect -4850 8293 -4830 8313
rect -4810 8293 -4790 8313
rect -4770 8293 -4750 8313
rect -4730 8293 -4710 8313
rect -4690 8293 -4670 8313
rect -4650 8293 -4630 8313
rect -4610 8293 -4590 8313
rect -4570 8293 -4550 8313
rect -4530 8293 -4510 8313
rect -4490 8293 -4470 8313
rect -4450 8293 -4430 8313
rect -4410 8293 -4390 8313
rect -4370 8293 -4350 8313
rect -4330 8293 -4310 8313
rect -4290 8293 -4270 8313
rect -4250 8293 -4230 8313
rect -4210 8293 -4190 8313
rect -4170 8293 -4150 8313
rect -4130 8293 -4110 8313
rect -4090 8293 -4070 8313
rect -4050 8293 -4030 8313
rect -4010 8293 -3990 8313
rect -3970 8293 -3950 8313
rect -3930 8293 -3910 8313
rect -3890 8293 -3870 8313
rect -3850 8293 -3830 8313
rect -3810 8293 -3790 8313
rect -3770 8293 -3750 8313
rect -3730 8293 -3710 8313
rect -3690 8293 -3670 8313
rect -3650 8293 -3630 8313
rect -3610 8293 -3590 8313
rect -3570 8293 -3550 8313
rect -3530 8293 -3510 8313
rect -3490 8293 -3470 8313
rect -3450 8293 -3430 8313
rect -3410 8293 -3390 8313
rect -3370 8293 -3350 8313
rect -3330 8293 -3310 8313
rect -3290 8293 -3270 8313
rect -3250 8293 -3230 8313
rect -3210 8293 -3190 8313
rect -5650 8211 -5630 8231
rect -5610 8211 -5590 8231
rect -5570 8211 -5550 8231
rect -5530 8211 -5510 8231
rect -5490 8211 -5470 8231
rect -5450 8211 -5430 8231
rect -5410 8211 -5390 8231
rect -5370 8211 -5350 8231
rect -5330 8211 -5310 8231
rect -5290 8211 -5270 8231
rect -5250 8211 -5230 8231
rect -5210 8211 -5190 8231
rect -5170 8211 -5150 8231
rect -5130 8211 -5110 8231
rect -5090 8211 -5070 8231
rect -5050 8211 -5030 8231
rect -5010 8211 -4990 8231
rect -4970 8211 -4950 8231
rect -4930 8211 -4910 8231
rect -4890 8211 -4870 8231
rect -4850 8211 -4830 8231
rect -4810 8211 -4790 8231
rect -4770 8211 -4750 8231
rect -4730 8211 -4710 8231
rect -4690 8211 -4670 8231
rect -4650 8211 -4630 8231
rect -4610 8211 -4590 8231
rect -4570 8211 -4550 8231
rect -4530 8211 -4510 8231
rect -4490 8211 -4470 8231
rect -4450 8211 -4430 8231
rect -4410 8211 -4390 8231
rect -4370 8211 -4350 8231
rect -4330 8211 -4310 8231
rect -4290 8211 -4270 8231
rect -4250 8211 -4230 8231
rect -4210 8211 -4190 8231
rect -4170 8211 -4150 8231
rect -4130 8211 -4110 8231
rect -4090 8211 -4070 8231
rect -4050 8211 -4030 8231
rect -4010 8211 -3990 8231
rect -3970 8211 -3950 8231
rect -3930 8211 -3910 8231
rect -3890 8211 -3870 8231
rect -3850 8211 -3830 8231
rect -3810 8211 -3790 8231
rect -3770 8211 -3750 8231
rect -3730 8211 -3710 8231
rect -3690 8211 -3670 8231
rect -3650 8211 -3630 8231
rect -3610 8211 -3590 8231
rect -3570 8211 -3550 8231
rect -3530 8211 -3510 8231
rect -3490 8211 -3470 8231
rect -3450 8211 -3430 8231
rect -3410 8211 -3390 8231
rect -3370 8211 -3350 8231
rect -3330 8211 -3310 8231
rect -3290 8211 -3270 8231
rect -3250 8211 -3230 8231
rect -3210 8211 -3190 8231
rect -5650 8129 -5630 8149
rect -5610 8129 -5590 8149
rect -5570 8129 -5550 8149
rect -5530 8129 -5510 8149
rect -5490 8129 -5470 8149
rect -5450 8129 -5430 8149
rect -5410 8129 -5390 8149
rect -5370 8129 -5350 8149
rect -5330 8129 -5310 8149
rect -5290 8129 -5270 8149
rect -5250 8129 -5230 8149
rect -5210 8129 -5190 8149
rect -5170 8129 -5150 8149
rect -5130 8129 -5110 8149
rect -5090 8129 -5070 8149
rect -5050 8129 -5030 8149
rect -5010 8129 -4990 8149
rect -4970 8129 -4950 8149
rect -4930 8129 -4910 8149
rect -4890 8129 -4870 8149
rect -4850 8129 -4830 8149
rect -4810 8129 -4790 8149
rect -4770 8129 -4750 8149
rect -4730 8129 -4710 8149
rect -4690 8129 -4670 8149
rect -4650 8129 -4630 8149
rect -4610 8129 -4590 8149
rect -4570 8129 -4550 8149
rect -4530 8129 -4510 8149
rect -4490 8129 -4470 8149
rect -4450 8129 -4430 8149
rect -4410 8129 -4390 8149
rect -4370 8129 -4350 8149
rect -4330 8129 -4310 8149
rect -4290 8129 -4270 8149
rect -4250 8129 -4230 8149
rect -4210 8129 -4190 8149
rect -4170 8129 -4150 8149
rect -4130 8129 -4110 8149
rect -4090 8129 -4070 8149
rect -4050 8129 -4030 8149
rect -4010 8129 -3990 8149
rect -3970 8129 -3950 8149
rect -3930 8129 -3910 8149
rect -3890 8129 -3870 8149
rect -3850 8129 -3830 8149
rect -3810 8129 -3790 8149
rect -3770 8129 -3750 8149
rect -3730 8129 -3710 8149
rect -3690 8129 -3670 8149
rect -3650 8129 -3630 8149
rect -3610 8129 -3590 8149
rect -3570 8129 -3550 8149
rect -3530 8129 -3510 8149
rect -3490 8129 -3470 8149
rect -3450 8129 -3430 8149
rect -3410 8129 -3390 8149
rect -3370 8129 -3350 8149
rect -3330 8129 -3310 8149
rect -3290 8129 -3270 8149
rect -3250 8129 -3230 8149
rect -3210 8129 -3190 8149
rect -5650 8047 -5630 8067
rect -5610 8047 -5590 8067
rect -5570 8047 -5550 8067
rect -5530 8047 -5510 8067
rect -5490 8047 -5470 8067
rect -5450 8047 -5430 8067
rect -5410 8047 -5390 8067
rect -5370 8047 -5350 8067
rect -5330 8047 -5310 8067
rect -5290 8047 -5270 8067
rect -5250 8047 -5230 8067
rect -5210 8047 -5190 8067
rect -5170 8047 -5150 8067
rect -5130 8047 -5110 8067
rect -5090 8047 -5070 8067
rect -5050 8047 -5030 8067
rect -5010 8047 -4990 8067
rect -4970 8047 -4950 8067
rect -4930 8047 -4910 8067
rect -4890 8047 -4870 8067
rect -4850 8047 -4830 8067
rect -4810 8047 -4790 8067
rect -4770 8047 -4750 8067
rect -4730 8047 -4710 8067
rect -4690 8047 -4670 8067
rect -4650 8047 -4630 8067
rect -4610 8047 -4590 8067
rect -4570 8047 -4550 8067
rect -4530 8047 -4510 8067
rect -4490 8047 -4470 8067
rect -4450 8047 -4430 8067
rect -4410 8047 -4390 8067
rect -4370 8047 -4350 8067
rect -4330 8047 -4310 8067
rect -4290 8047 -4270 8067
rect -4250 8047 -4230 8067
rect -4210 8047 -4190 8067
rect -4170 8047 -4150 8067
rect -4130 8047 -4110 8067
rect -4090 8047 -4070 8067
rect -4050 8047 -4030 8067
rect -4010 8047 -3990 8067
rect -3970 8047 -3950 8067
rect -3930 8047 -3910 8067
rect -3890 8047 -3870 8067
rect -3850 8047 -3830 8067
rect -3810 8047 -3790 8067
rect -3770 8047 -3750 8067
rect -3730 8047 -3710 8067
rect -3690 8047 -3670 8067
rect -3650 8047 -3630 8067
rect -3610 8047 -3590 8067
rect -3570 8047 -3550 8067
rect -3530 8047 -3510 8067
rect -3490 8047 -3470 8067
rect -3450 8047 -3430 8067
rect -3410 8047 -3390 8067
rect -3370 8047 -3350 8067
rect -3330 8047 -3310 8067
rect -3290 8047 -3270 8067
rect -3250 8047 -3230 8067
rect -3210 8047 -3190 8067
rect -5650 7965 -5630 7985
rect -5610 7965 -5590 7985
rect -5570 7965 -5550 7985
rect -5530 7965 -5510 7985
rect -5490 7965 -5470 7985
rect -5450 7965 -5430 7985
rect -5410 7965 -5390 7985
rect -5370 7965 -5350 7985
rect -5330 7965 -5310 7985
rect -5290 7965 -5270 7985
rect -5250 7965 -5230 7985
rect -5210 7965 -5190 7985
rect -5170 7965 -5150 7985
rect -5130 7965 -5110 7985
rect -5090 7965 -5070 7985
rect -5050 7965 -5030 7985
rect -5010 7965 -4990 7985
rect -4970 7965 -4950 7985
rect -4930 7965 -4910 7985
rect -4890 7965 -4870 7985
rect -4850 7965 -4830 7985
rect -4810 7965 -4790 7985
rect -4770 7965 -4750 7985
rect -4730 7965 -4710 7985
rect -4690 7965 -4670 7985
rect -4650 7965 -4630 7985
rect -4610 7965 -4590 7985
rect -4570 7965 -4550 7985
rect -4530 7965 -4510 7985
rect -4490 7965 -4470 7985
rect -4450 7965 -4430 7985
rect -4410 7965 -4390 7985
rect -4370 7965 -4350 7985
rect -4330 7965 -4310 7985
rect -4290 7965 -4270 7985
rect -4250 7965 -4230 7985
rect -4210 7965 -4190 7985
rect -4170 7965 -4150 7985
rect -4130 7965 -4110 7985
rect -4090 7965 -4070 7985
rect -4050 7965 -4030 7985
rect -4010 7965 -3990 7985
rect -3970 7965 -3950 7985
rect -3930 7965 -3910 7985
rect -3890 7965 -3870 7985
rect -3850 7965 -3830 7985
rect -3810 7965 -3790 7985
rect -3770 7965 -3750 7985
rect -3730 7965 -3710 7985
rect -3690 7965 -3670 7985
rect -3650 7965 -3630 7985
rect -3610 7965 -3590 7985
rect -3570 7965 -3550 7985
rect -3530 7965 -3510 7985
rect -3490 7965 -3470 7985
rect -3450 7965 -3430 7985
rect -3410 7965 -3390 7985
rect -3370 7965 -3350 7985
rect -3330 7965 -3310 7985
rect -3290 7965 -3270 7985
rect -3250 7965 -3230 7985
rect -3210 7965 -3190 7985
rect -5650 7883 -5630 7903
rect -5610 7883 -5590 7903
rect -5570 7883 -5550 7903
rect -5530 7883 -5510 7903
rect -5490 7883 -5470 7903
rect -5450 7883 -5430 7903
rect -5410 7883 -5390 7903
rect -5370 7883 -5350 7903
rect -5330 7883 -5310 7903
rect -5290 7883 -5270 7903
rect -5250 7883 -5230 7903
rect -5210 7883 -5190 7903
rect -5170 7883 -5150 7903
rect -5130 7883 -5110 7903
rect -5090 7883 -5070 7903
rect -5050 7883 -5030 7903
rect -5010 7883 -4990 7903
rect -4970 7883 -4950 7903
rect -4930 7883 -4910 7903
rect -4890 7883 -4870 7903
rect -4850 7883 -4830 7903
rect -4810 7883 -4790 7903
rect -4770 7883 -4750 7903
rect -4730 7883 -4710 7903
rect -4690 7883 -4670 7903
rect -4650 7883 -4630 7903
rect -4610 7883 -4590 7903
rect -4570 7883 -4550 7903
rect -4530 7883 -4510 7903
rect -4490 7883 -4470 7903
rect -4450 7883 -4430 7903
rect -4410 7883 -4390 7903
rect -4370 7883 -4350 7903
rect -4330 7883 -4310 7903
rect -4290 7883 -4270 7903
rect -4250 7883 -4230 7903
rect -4210 7883 -4190 7903
rect -4170 7883 -4150 7903
rect -4130 7883 -4110 7903
rect -4090 7883 -4070 7903
rect -4050 7883 -4030 7903
rect -4010 7883 -3990 7903
rect -3970 7883 -3950 7903
rect -3930 7883 -3910 7903
rect -3890 7883 -3870 7903
rect -3850 7883 -3830 7903
rect -3810 7883 -3790 7903
rect -3770 7883 -3750 7903
rect -3730 7883 -3710 7903
rect -3690 7883 -3670 7903
rect -3650 7883 -3630 7903
rect -3610 7883 -3590 7903
rect -3570 7883 -3550 7903
rect -3530 7883 -3510 7903
rect -3490 7883 -3470 7903
rect -3450 7883 -3430 7903
rect -3410 7883 -3390 7903
rect -3370 7883 -3350 7903
rect -3330 7883 -3310 7903
rect -3290 7883 -3270 7903
rect -3250 7883 -3230 7903
rect -3210 7883 -3190 7903
rect -5650 7801 -5630 7821
rect -5610 7801 -5590 7821
rect -5570 7801 -5550 7821
rect -5530 7801 -5510 7821
rect -5490 7801 -5470 7821
rect -5450 7801 -5430 7821
rect -5410 7801 -5390 7821
rect -5370 7801 -5350 7821
rect -5330 7801 -5310 7821
rect -5290 7801 -5270 7821
rect -5250 7801 -5230 7821
rect -5210 7801 -5190 7821
rect -5170 7801 -5150 7821
rect -5130 7801 -5110 7821
rect -5090 7801 -5070 7821
rect -5050 7801 -5030 7821
rect -5010 7801 -4990 7821
rect -4970 7801 -4950 7821
rect -4930 7801 -4910 7821
rect -4890 7801 -4870 7821
rect -4850 7801 -4830 7821
rect -4810 7801 -4790 7821
rect -4770 7801 -4750 7821
rect -4730 7801 -4710 7821
rect -4690 7801 -4670 7821
rect -4650 7801 -4630 7821
rect -4610 7801 -4590 7821
rect -4570 7801 -4550 7821
rect -4530 7801 -4510 7821
rect -4490 7801 -4470 7821
rect -4450 7801 -4430 7821
rect -4410 7801 -4390 7821
rect -4370 7801 -4350 7821
rect -4330 7801 -4310 7821
rect -4290 7801 -4270 7821
rect -4250 7801 -4230 7821
rect -4210 7801 -4190 7821
rect -4170 7801 -4150 7821
rect -4130 7801 -4110 7821
rect -4090 7801 -4070 7821
rect -4050 7801 -4030 7821
rect -4010 7801 -3990 7821
rect -3970 7801 -3950 7821
rect -3930 7801 -3910 7821
rect -3890 7801 -3870 7821
rect -3850 7801 -3830 7821
rect -3810 7801 -3790 7821
rect -3770 7801 -3750 7821
rect -3730 7801 -3710 7821
rect -3690 7801 -3670 7821
rect -3650 7801 -3630 7821
rect -3610 7801 -3590 7821
rect -3570 7801 -3550 7821
rect -3530 7801 -3510 7821
rect -3490 7801 -3470 7821
rect -3450 7801 -3430 7821
rect -3410 7801 -3390 7821
rect -3370 7801 -3350 7821
rect -3330 7801 -3310 7821
rect -3290 7801 -3270 7821
rect -3250 7801 -3230 7821
rect -3210 7801 -3190 7821
rect -5650 7719 -5630 7739
rect -5610 7719 -5590 7739
rect -5570 7719 -5550 7739
rect -5530 7719 -5510 7739
rect -5490 7719 -5470 7739
rect -5450 7719 -5430 7739
rect -5410 7719 -5390 7739
rect -5370 7719 -5350 7739
rect -5330 7719 -5310 7739
rect -5290 7719 -5270 7739
rect -5250 7719 -5230 7739
rect -5210 7719 -5190 7739
rect -5170 7719 -5150 7739
rect -5130 7719 -5110 7739
rect -5090 7719 -5070 7739
rect -5050 7719 -5030 7739
rect -5010 7719 -4990 7739
rect -4970 7719 -4950 7739
rect -4930 7719 -4910 7739
rect -4890 7719 -4870 7739
rect -4850 7719 -4830 7739
rect -4810 7719 -4790 7739
rect -4770 7719 -4750 7739
rect -4730 7719 -4710 7739
rect -4690 7719 -4670 7739
rect -4650 7719 -4630 7739
rect -4610 7719 -4590 7739
rect -4570 7719 -4550 7739
rect -4530 7719 -4510 7739
rect -4490 7719 -4470 7739
rect -4450 7719 -4430 7739
rect -4410 7719 -4390 7739
rect -4370 7719 -4350 7739
rect -4330 7719 -4310 7739
rect -4290 7719 -4270 7739
rect -4250 7719 -4230 7739
rect -4210 7719 -4190 7739
rect -4170 7719 -4150 7739
rect -4130 7719 -4110 7739
rect -4090 7719 -4070 7739
rect -4050 7719 -4030 7739
rect -4010 7719 -3990 7739
rect -3970 7719 -3950 7739
rect -3930 7719 -3910 7739
rect -3890 7719 -3870 7739
rect -3850 7719 -3830 7739
rect -3810 7719 -3790 7739
rect -3770 7719 -3750 7739
rect -3730 7719 -3710 7739
rect -3690 7719 -3670 7739
rect -3650 7719 -3630 7739
rect -3610 7719 -3590 7739
rect -3570 7719 -3550 7739
rect -3530 7719 -3510 7739
rect -3490 7719 -3470 7739
rect -3450 7719 -3430 7739
rect -3410 7719 -3390 7739
rect -3370 7719 -3350 7739
rect -3330 7719 -3310 7739
rect -3290 7719 -3270 7739
rect -3250 7719 -3230 7739
rect -3210 7719 -3190 7739
rect -5650 7637 -5630 7657
rect -5610 7637 -5590 7657
rect -5570 7637 -5550 7657
rect -5530 7637 -5510 7657
rect -5490 7637 -5470 7657
rect -5450 7637 -5430 7657
rect -5410 7637 -5390 7657
rect -5370 7637 -5350 7657
rect -5330 7637 -5310 7657
rect -5290 7637 -5270 7657
rect -5250 7637 -5230 7657
rect -5210 7637 -5190 7657
rect -5170 7637 -5150 7657
rect -5130 7637 -5110 7657
rect -5090 7637 -5070 7657
rect -5050 7637 -5030 7657
rect -5010 7637 -4990 7657
rect -4970 7637 -4950 7657
rect -4930 7637 -4910 7657
rect -4890 7637 -4870 7657
rect -4850 7637 -4830 7657
rect -4810 7637 -4790 7657
rect -4770 7637 -4750 7657
rect -4730 7637 -4710 7657
rect -4690 7637 -4670 7657
rect -4650 7637 -4630 7657
rect -4610 7637 -4590 7657
rect -4570 7637 -4550 7657
rect -4530 7637 -4510 7657
rect -4490 7637 -4470 7657
rect -4450 7637 -4430 7657
rect -4410 7637 -4390 7657
rect -4370 7637 -4350 7657
rect -4330 7637 -4310 7657
rect -4290 7637 -4270 7657
rect -4250 7637 -4230 7657
rect -4210 7637 -4190 7657
rect -4170 7637 -4150 7657
rect -4130 7637 -4110 7657
rect -4090 7637 -4070 7657
rect -4050 7637 -4030 7657
rect -4010 7637 -3990 7657
rect -3970 7637 -3950 7657
rect -3930 7637 -3910 7657
rect -3890 7637 -3870 7657
rect -3850 7637 -3830 7657
rect -3810 7637 -3790 7657
rect -3770 7637 -3750 7657
rect -3730 7637 -3710 7657
rect -3690 7637 -3670 7657
rect -3650 7637 -3630 7657
rect -3610 7637 -3590 7657
rect -3570 7637 -3550 7657
rect -3530 7637 -3510 7657
rect -3490 7637 -3470 7657
rect -3450 7637 -3430 7657
rect -3410 7637 -3390 7657
rect -3370 7637 -3350 7657
rect -3330 7637 -3310 7657
rect -3290 7637 -3270 7657
rect -3250 7637 -3230 7657
rect -3210 7637 -3190 7657
rect -5650 7555 -5630 7575
rect -5610 7555 -5590 7575
rect -5570 7555 -5550 7575
rect -5530 7555 -5510 7575
rect -5490 7555 -5470 7575
rect -5450 7555 -5430 7575
rect -5410 7555 -5390 7575
rect -5370 7555 -5350 7575
rect -5330 7555 -5310 7575
rect -5290 7555 -5270 7575
rect -5250 7555 -5230 7575
rect -5210 7555 -5190 7575
rect -5170 7555 -5150 7575
rect -5130 7555 -5110 7575
rect -5090 7555 -5070 7575
rect -5050 7555 -5030 7575
rect -5010 7555 -4990 7575
rect -4970 7555 -4950 7575
rect -4930 7555 -4910 7575
rect -4890 7555 -4870 7575
rect -4850 7555 -4830 7575
rect -4810 7555 -4790 7575
rect -4770 7555 -4750 7575
rect -4730 7555 -4710 7575
rect -4690 7555 -4670 7575
rect -4650 7555 -4630 7575
rect -4610 7555 -4590 7575
rect -4570 7555 -4550 7575
rect -4530 7555 -4510 7575
rect -4490 7555 -4470 7575
rect -4450 7555 -4430 7575
rect -4410 7555 -4390 7575
rect -4370 7555 -4350 7575
rect -4330 7555 -4310 7575
rect -4290 7555 -4270 7575
rect -4250 7555 -4230 7575
rect -4210 7555 -4190 7575
rect -4170 7555 -4150 7575
rect -4130 7555 -4110 7575
rect -4090 7555 -4070 7575
rect -4050 7555 -4030 7575
rect -4010 7555 -3990 7575
rect -3970 7555 -3950 7575
rect -3930 7555 -3910 7575
rect -3890 7555 -3870 7575
rect -3850 7555 -3830 7575
rect -3810 7555 -3790 7575
rect -3770 7555 -3750 7575
rect -3730 7555 -3710 7575
rect -3690 7555 -3670 7575
rect -3650 7555 -3630 7575
rect -3610 7555 -3590 7575
rect -3570 7555 -3550 7575
rect -3530 7555 -3510 7575
rect -3490 7555 -3470 7575
rect -3450 7555 -3430 7575
rect -3410 7555 -3390 7575
rect -3370 7555 -3350 7575
rect -3330 7555 -3310 7575
rect -3290 7555 -3270 7575
rect -3250 7555 -3230 7575
rect -3210 7555 -3190 7575
rect -5650 7473 -5630 7493
rect -5610 7473 -5590 7493
rect -5570 7473 -5550 7493
rect -5530 7473 -5510 7493
rect -5490 7473 -5470 7493
rect -5450 7473 -5430 7493
rect -5410 7473 -5390 7493
rect -5370 7473 -5350 7493
rect -5330 7473 -5310 7493
rect -5290 7473 -5270 7493
rect -5250 7473 -5230 7493
rect -5210 7473 -5190 7493
rect -5170 7473 -5150 7493
rect -5130 7473 -5110 7493
rect -5090 7473 -5070 7493
rect -5050 7473 -5030 7493
rect -5010 7473 -4990 7493
rect -4970 7473 -4950 7493
rect -4930 7473 -4910 7493
rect -4890 7473 -4870 7493
rect -4850 7473 -4830 7493
rect -4810 7473 -4790 7493
rect -4770 7473 -4750 7493
rect -4730 7473 -4710 7493
rect -4690 7473 -4670 7493
rect -4650 7473 -4630 7493
rect -4610 7473 -4590 7493
rect -4570 7473 -4550 7493
rect -4530 7473 -4510 7493
rect -4490 7473 -4470 7493
rect -4450 7473 -4430 7493
rect -4410 7473 -4390 7493
rect -4370 7473 -4350 7493
rect -4330 7473 -4310 7493
rect -4290 7473 -4270 7493
rect -4250 7473 -4230 7493
rect -4210 7473 -4190 7493
rect -4170 7473 -4150 7493
rect -4130 7473 -4110 7493
rect -4090 7473 -4070 7493
rect -4050 7473 -4030 7493
rect -4010 7473 -3990 7493
rect -3970 7473 -3950 7493
rect -3930 7473 -3910 7493
rect -3890 7473 -3870 7493
rect -3850 7473 -3830 7493
rect -3810 7473 -3790 7493
rect -3770 7473 -3750 7493
rect -3730 7473 -3710 7493
rect -3690 7473 -3670 7493
rect -3650 7473 -3630 7493
rect -3610 7473 -3590 7493
rect -3570 7473 -3550 7493
rect -3530 7473 -3510 7493
rect -3490 7473 -3470 7493
rect -3450 7473 -3430 7493
rect -3410 7473 -3390 7493
rect -3370 7473 -3350 7493
rect -3330 7473 -3310 7493
rect -3290 7473 -3270 7493
rect -3250 7473 -3230 7493
rect -3210 7473 -3190 7493
rect -5650 7391 -5630 7411
rect -5610 7391 -5590 7411
rect -5570 7391 -5550 7411
rect -5530 7391 -5510 7411
rect -5490 7391 -5470 7411
rect -5450 7391 -5430 7411
rect -5410 7391 -5390 7411
rect -5370 7391 -5350 7411
rect -5330 7391 -5310 7411
rect -5290 7391 -5270 7411
rect -5250 7391 -5230 7411
rect -5210 7391 -5190 7411
rect -5170 7391 -5150 7411
rect -5130 7391 -5110 7411
rect -5090 7391 -5070 7411
rect -5050 7391 -5030 7411
rect -5010 7391 -4990 7411
rect -4970 7391 -4950 7411
rect -4930 7391 -4910 7411
rect -4890 7391 -4870 7411
rect -4850 7391 -4830 7411
rect -4810 7391 -4790 7411
rect -4770 7391 -4750 7411
rect -4730 7391 -4710 7411
rect -4690 7391 -4670 7411
rect -4650 7391 -4630 7411
rect -4610 7391 -4590 7411
rect -4570 7391 -4550 7411
rect -4530 7391 -4510 7411
rect -4490 7391 -4470 7411
rect -4450 7391 -4430 7411
rect -4410 7391 -4390 7411
rect -4370 7391 -4350 7411
rect -4330 7391 -4310 7411
rect -4290 7391 -4270 7411
rect -4250 7391 -4230 7411
rect -4210 7391 -4190 7411
rect -4170 7391 -4150 7411
rect -4130 7391 -4110 7411
rect -4090 7391 -4070 7411
rect -4050 7391 -4030 7411
rect -4010 7391 -3990 7411
rect -3970 7391 -3950 7411
rect -3930 7391 -3910 7411
rect -3890 7391 -3870 7411
rect -3850 7391 -3830 7411
rect -3810 7391 -3790 7411
rect -3770 7391 -3750 7411
rect -3730 7391 -3710 7411
rect -3690 7391 -3670 7411
rect -3650 7391 -3630 7411
rect -3610 7391 -3590 7411
rect -3570 7391 -3550 7411
rect -3530 7391 -3510 7411
rect -3490 7391 -3470 7411
rect -3450 7391 -3430 7411
rect -3410 7391 -3390 7411
rect -3370 7391 -3350 7411
rect -3330 7391 -3310 7411
rect -3290 7391 -3270 7411
rect -3250 7391 -3230 7411
rect -3210 7391 -3190 7411
rect -5650 7309 -5630 7329
rect -5610 7309 -5590 7329
rect -5570 7309 -5550 7329
rect -5530 7309 -5510 7329
rect -5490 7309 -5470 7329
rect -5450 7309 -5430 7329
rect -5410 7309 -5390 7329
rect -5370 7309 -5350 7329
rect -5330 7309 -5310 7329
rect -5290 7309 -5270 7329
rect -5250 7309 -5230 7329
rect -5210 7309 -5190 7329
rect -5170 7309 -5150 7329
rect -5130 7309 -5110 7329
rect -5090 7309 -5070 7329
rect -5050 7309 -5030 7329
rect -5010 7309 -4990 7329
rect -4970 7309 -4950 7329
rect -4930 7309 -4910 7329
rect -4890 7309 -4870 7329
rect -4850 7309 -4830 7329
rect -4810 7309 -4790 7329
rect -4770 7309 -4750 7329
rect -4730 7309 -4710 7329
rect -4690 7309 -4670 7329
rect -4650 7309 -4630 7329
rect -4610 7309 -4590 7329
rect -4570 7309 -4550 7329
rect -4530 7309 -4510 7329
rect -4490 7309 -4470 7329
rect -4450 7309 -4430 7329
rect -4410 7309 -4390 7329
rect -4370 7309 -4350 7329
rect -4330 7309 -4310 7329
rect -4290 7309 -4270 7329
rect -4250 7309 -4230 7329
rect -4210 7309 -4190 7329
rect -4170 7309 -4150 7329
rect -4130 7309 -4110 7329
rect -4090 7309 -4070 7329
rect -4050 7309 -4030 7329
rect -4010 7309 -3990 7329
rect -3970 7309 -3950 7329
rect -3930 7309 -3910 7329
rect -3890 7309 -3870 7329
rect -3850 7309 -3830 7329
rect -3810 7309 -3790 7329
rect -3770 7309 -3750 7329
rect -3730 7309 -3710 7329
rect -3690 7309 -3670 7329
rect -3650 7309 -3630 7329
rect -3610 7309 -3590 7329
rect -3570 7309 -3550 7329
rect -3530 7309 -3510 7329
rect -3490 7309 -3470 7329
rect -3450 7309 -3430 7329
rect -3410 7309 -3390 7329
rect -3370 7309 -3350 7329
rect -3330 7309 -3310 7329
rect -3290 7309 -3270 7329
rect -3250 7309 -3230 7329
rect -3210 7309 -3190 7329
rect -5650 7227 -5630 7247
rect -5610 7227 -5590 7247
rect -5570 7227 -5550 7247
rect -5530 7227 -5510 7247
rect -5490 7227 -5470 7247
rect -5450 7227 -5430 7247
rect -5410 7227 -5390 7247
rect -5370 7227 -5350 7247
rect -5330 7227 -5310 7247
rect -5290 7227 -5270 7247
rect -5250 7227 -5230 7247
rect -5210 7227 -5190 7247
rect -5170 7227 -5150 7247
rect -5130 7227 -5110 7247
rect -5090 7227 -5070 7247
rect -5050 7227 -5030 7247
rect -5010 7227 -4990 7247
rect -4970 7227 -4950 7247
rect -4930 7227 -4910 7247
rect -4890 7227 -4870 7247
rect -4850 7227 -4830 7247
rect -4810 7227 -4790 7247
rect -4770 7227 -4750 7247
rect -4730 7227 -4710 7247
rect -4690 7227 -4670 7247
rect -4650 7227 -4630 7247
rect -4610 7227 -4590 7247
rect -4570 7227 -4550 7247
rect -4530 7227 -4510 7247
rect -4490 7227 -4470 7247
rect -4450 7227 -4430 7247
rect -4410 7227 -4390 7247
rect -4370 7227 -4350 7247
rect -4330 7227 -4310 7247
rect -4290 7227 -4270 7247
rect -4250 7227 -4230 7247
rect -4210 7227 -4190 7247
rect -4170 7227 -4150 7247
rect -4130 7227 -4110 7247
rect -4090 7227 -4070 7247
rect -4050 7227 -4030 7247
rect -4010 7227 -3990 7247
rect -3970 7227 -3950 7247
rect -3930 7227 -3910 7247
rect -3890 7227 -3870 7247
rect -3850 7227 -3830 7247
rect -3810 7227 -3790 7247
rect -3770 7227 -3750 7247
rect -3730 7227 -3710 7247
rect -3690 7227 -3670 7247
rect -3650 7227 -3630 7247
rect -3610 7227 -3590 7247
rect -3570 7227 -3550 7247
rect -3530 7227 -3510 7247
rect -3490 7227 -3470 7247
rect -3450 7227 -3430 7247
rect -3410 7227 -3390 7247
rect -3370 7227 -3350 7247
rect -3330 7227 -3310 7247
rect -3290 7227 -3270 7247
rect -3250 7227 -3230 7247
rect -3210 7227 -3190 7247
rect -5650 7145 -5630 7165
rect -5610 7145 -5590 7165
rect -5570 7145 -5550 7165
rect -5530 7145 -5510 7165
rect -5490 7145 -5470 7165
rect -5450 7145 -5430 7165
rect -5410 7145 -5390 7165
rect -5370 7145 -5350 7165
rect -5330 7145 -5310 7165
rect -5290 7145 -5270 7165
rect -5250 7145 -5230 7165
rect -5210 7145 -5190 7165
rect -5170 7145 -5150 7165
rect -5130 7145 -5110 7165
rect -5090 7145 -5070 7165
rect -5050 7145 -5030 7165
rect -5010 7145 -4990 7165
rect -4970 7145 -4950 7165
rect -4930 7145 -4910 7165
rect -4890 7145 -4870 7165
rect -4850 7145 -4830 7165
rect -4810 7145 -4790 7165
rect -4770 7145 -4750 7165
rect -4730 7145 -4710 7165
rect -4690 7145 -4670 7165
rect -4650 7145 -4630 7165
rect -4610 7145 -4590 7165
rect -4570 7145 -4550 7165
rect -4530 7145 -4510 7165
rect -4490 7145 -4470 7165
rect -4450 7145 -4430 7165
rect -4410 7145 -4390 7165
rect -4370 7145 -4350 7165
rect -4330 7145 -4310 7165
rect -4290 7145 -4270 7165
rect -4250 7145 -4230 7165
rect -4210 7145 -4190 7165
rect -4170 7145 -4150 7165
rect -4130 7145 -4110 7165
rect -4090 7145 -4070 7165
rect -4050 7145 -4030 7165
rect -4010 7145 -3990 7165
rect -3970 7145 -3950 7165
rect -3930 7145 -3910 7165
rect -3890 7145 -3870 7165
rect -3850 7145 -3830 7165
rect -3810 7145 -3790 7165
rect -3770 7145 -3750 7165
rect -3730 7145 -3710 7165
rect -3690 7145 -3670 7165
rect -3650 7145 -3630 7165
rect -3610 7145 -3590 7165
rect -3570 7145 -3550 7165
rect -3530 7145 -3510 7165
rect -3490 7145 -3470 7165
rect -3450 7145 -3430 7165
rect -3410 7145 -3390 7165
rect -3370 7145 -3350 7165
rect -3330 7145 -3310 7165
rect -3290 7145 -3270 7165
rect -3250 7145 -3230 7165
rect -3210 7145 -3190 7165
rect -5650 7063 -5630 7083
rect -5610 7063 -5590 7083
rect -5570 7063 -5550 7083
rect -5530 7063 -5510 7083
rect -5490 7063 -5470 7083
rect -5450 7063 -5430 7083
rect -5410 7063 -5390 7083
rect -5370 7063 -5350 7083
rect -5330 7063 -5310 7083
rect -5290 7063 -5270 7083
rect -5250 7063 -5230 7083
rect -5210 7063 -5190 7083
rect -5170 7063 -5150 7083
rect -5130 7063 -5110 7083
rect -5090 7063 -5070 7083
rect -5050 7063 -5030 7083
rect -5010 7063 -4990 7083
rect -4970 7063 -4950 7083
rect -4930 7063 -4910 7083
rect -4890 7063 -4870 7083
rect -4850 7063 -4830 7083
rect -4810 7063 -4790 7083
rect -4770 7063 -4750 7083
rect -4730 7063 -4710 7083
rect -4690 7063 -4670 7083
rect -4650 7063 -4630 7083
rect -4610 7063 -4590 7083
rect -4570 7063 -4550 7083
rect -4530 7063 -4510 7083
rect -4490 7063 -4470 7083
rect -4450 7063 -4430 7083
rect -4410 7063 -4390 7083
rect -4370 7063 -4350 7083
rect -4330 7063 -4310 7083
rect -4290 7063 -4270 7083
rect -4250 7063 -4230 7083
rect -4210 7063 -4190 7083
rect -4170 7063 -4150 7083
rect -4130 7063 -4110 7083
rect -4090 7063 -4070 7083
rect -4050 7063 -4030 7083
rect -4010 7063 -3990 7083
rect -3970 7063 -3950 7083
rect -3930 7063 -3910 7083
rect -3890 7063 -3870 7083
rect -3850 7063 -3830 7083
rect -3810 7063 -3790 7083
rect -3770 7063 -3750 7083
rect -3730 7063 -3710 7083
rect -3690 7063 -3670 7083
rect -3650 7063 -3630 7083
rect -3610 7063 -3590 7083
rect -3570 7063 -3550 7083
rect -3530 7063 -3510 7083
rect -3490 7063 -3470 7083
rect -3450 7063 -3430 7083
rect -3410 7063 -3390 7083
rect -3370 7063 -3350 7083
rect -3330 7063 -3310 7083
rect -3290 7063 -3270 7083
rect -3250 7063 -3230 7083
rect -3210 7063 -3190 7083
rect -5650 6981 -5630 7001
rect -5610 6981 -5590 7001
rect -5570 6981 -5550 7001
rect -5530 6981 -5510 7001
rect -5490 6981 -5470 7001
rect -5450 6981 -5430 7001
rect -5410 6981 -5390 7001
rect -5370 6981 -5350 7001
rect -5330 6981 -5310 7001
rect -5290 6981 -5270 7001
rect -5250 6981 -5230 7001
rect -5210 6981 -5190 7001
rect -5170 6981 -5150 7001
rect -5130 6981 -5110 7001
rect -5090 6981 -5070 7001
rect -5050 6981 -5030 7001
rect -5010 6981 -4990 7001
rect -4970 6981 -4950 7001
rect -4930 6981 -4910 7001
rect -4890 6981 -4870 7001
rect -4850 6981 -4830 7001
rect -4810 6981 -4790 7001
rect -4770 6981 -4750 7001
rect -4730 6981 -4710 7001
rect -4690 6981 -4670 7001
rect -4650 6981 -4630 7001
rect -4610 6981 -4590 7001
rect -4570 6981 -4550 7001
rect -4530 6981 -4510 7001
rect -4490 6981 -4470 7001
rect -4450 6981 -4430 7001
rect -4410 6981 -4390 7001
rect -4370 6981 -4350 7001
rect -4330 6981 -4310 7001
rect -4290 6981 -4270 7001
rect -4250 6981 -4230 7001
rect -4210 6981 -4190 7001
rect -4170 6981 -4150 7001
rect -4130 6981 -4110 7001
rect -4090 6981 -4070 7001
rect -4050 6981 -4030 7001
rect -4010 6981 -3990 7001
rect -3970 6981 -3950 7001
rect -3930 6981 -3910 7001
rect -3890 6981 -3870 7001
rect -3850 6981 -3830 7001
rect -3810 6981 -3790 7001
rect -3770 6981 -3750 7001
rect -3730 6981 -3710 7001
rect -3690 6981 -3670 7001
rect -3650 6981 -3630 7001
rect -3610 6981 -3590 7001
rect -3570 6981 -3550 7001
rect -3530 6981 -3510 7001
rect -3490 6981 -3470 7001
rect -3450 6981 -3430 7001
rect -3410 6981 -3390 7001
rect -3370 6981 -3350 7001
rect -3330 6981 -3310 7001
rect -3290 6981 -3270 7001
rect -3250 6981 -3230 7001
rect -3210 6981 -3190 7001
rect -5650 6899 -5630 6919
rect -5610 6899 -5590 6919
rect -5570 6899 -5550 6919
rect -5530 6899 -5510 6919
rect -5490 6899 -5470 6919
rect -5450 6899 -5430 6919
rect -5410 6899 -5390 6919
rect -5370 6899 -5350 6919
rect -5330 6899 -5310 6919
rect -5290 6899 -5270 6919
rect -5250 6899 -5230 6919
rect -5210 6899 -5190 6919
rect -5170 6899 -5150 6919
rect -5130 6899 -5110 6919
rect -5090 6899 -5070 6919
rect -5050 6899 -5030 6919
rect -5010 6899 -4990 6919
rect -4970 6899 -4950 6919
rect -4930 6899 -4910 6919
rect -4890 6899 -4870 6919
rect -4850 6899 -4830 6919
rect -4810 6899 -4790 6919
rect -4770 6899 -4750 6919
rect -4730 6899 -4710 6919
rect -4690 6899 -4670 6919
rect -4650 6899 -4630 6919
rect -4610 6899 -4590 6919
rect -4570 6899 -4550 6919
rect -4530 6899 -4510 6919
rect -4490 6899 -4470 6919
rect -4450 6899 -4430 6919
rect -4410 6899 -4390 6919
rect -4370 6899 -4350 6919
rect -4330 6899 -4310 6919
rect -4290 6899 -4270 6919
rect -4250 6899 -4230 6919
rect -4210 6899 -4190 6919
rect -4170 6899 -4150 6919
rect -4130 6899 -4110 6919
rect -4090 6899 -4070 6919
rect -4050 6899 -4030 6919
rect -4010 6899 -3990 6919
rect -3970 6899 -3950 6919
rect -3930 6899 -3910 6919
rect -3890 6899 -3870 6919
rect -3850 6899 -3830 6919
rect -3810 6899 -3790 6919
rect -3770 6899 -3750 6919
rect -3730 6899 -3710 6919
rect -3690 6899 -3670 6919
rect -3650 6899 -3630 6919
rect -3610 6899 -3590 6919
rect -3570 6899 -3550 6919
rect -3530 6899 -3510 6919
rect -3490 6899 -3470 6919
rect -3450 6899 -3430 6919
rect -3410 6899 -3390 6919
rect -3370 6899 -3350 6919
rect -3330 6899 -3310 6919
rect -3290 6899 -3270 6919
rect -3250 6899 -3230 6919
rect -3210 6899 -3190 6919
rect -5650 6817 -5630 6837
rect -5610 6817 -5590 6837
rect -5570 6817 -5550 6837
rect -5530 6817 -5510 6837
rect -5490 6817 -5470 6837
rect -5450 6817 -5430 6837
rect -5410 6817 -5390 6837
rect -5370 6817 -5350 6837
rect -5330 6817 -5310 6837
rect -5290 6817 -5270 6837
rect -5250 6817 -5230 6837
rect -5210 6817 -5190 6837
rect -5170 6817 -5150 6837
rect -5130 6817 -5110 6837
rect -5090 6817 -5070 6837
rect -5050 6817 -5030 6837
rect -5010 6817 -4990 6837
rect -4970 6817 -4950 6837
rect -4930 6817 -4910 6837
rect -4890 6817 -4870 6837
rect -4850 6817 -4830 6837
rect -4810 6817 -4790 6837
rect -4770 6817 -4750 6837
rect -4730 6817 -4710 6837
rect -4690 6817 -4670 6837
rect -4650 6817 -4630 6837
rect -4610 6817 -4590 6837
rect -4570 6817 -4550 6837
rect -4530 6817 -4510 6837
rect -4490 6817 -4470 6837
rect -4450 6817 -4430 6837
rect -4410 6817 -4390 6837
rect -4370 6817 -4350 6837
rect -4330 6817 -4310 6837
rect -4290 6817 -4270 6837
rect -4250 6817 -4230 6837
rect -4210 6817 -4190 6837
rect -4170 6817 -4150 6837
rect -4130 6817 -4110 6837
rect -4090 6817 -4070 6837
rect -4050 6817 -4030 6837
rect -4010 6817 -3990 6837
rect -3970 6817 -3950 6837
rect -3930 6817 -3910 6837
rect -3890 6817 -3870 6837
rect -3850 6817 -3830 6837
rect -3810 6817 -3790 6837
rect -3770 6817 -3750 6837
rect -3730 6817 -3710 6837
rect -3690 6817 -3670 6837
rect -3650 6817 -3630 6837
rect -3610 6817 -3590 6837
rect -3570 6817 -3550 6837
rect -3530 6817 -3510 6837
rect -3490 6817 -3470 6837
rect -3450 6817 -3430 6837
rect -3410 6817 -3390 6837
rect -3370 6817 -3350 6837
rect -3330 6817 -3310 6837
rect -3290 6817 -3270 6837
rect -3250 6817 -3230 6837
rect -3210 6817 -3190 6837
rect -5650 6735 -5630 6755
rect -5610 6735 -5590 6755
rect -5570 6735 -5550 6755
rect -5530 6735 -5510 6755
rect -5490 6735 -5470 6755
rect -5450 6735 -5430 6755
rect -5410 6735 -5390 6755
rect -5370 6735 -5350 6755
rect -5330 6735 -5310 6755
rect -5290 6735 -5270 6755
rect -5250 6735 -5230 6755
rect -5210 6735 -5190 6755
rect -5170 6735 -5150 6755
rect -5130 6735 -5110 6755
rect -5090 6735 -5070 6755
rect -5050 6735 -5030 6755
rect -5010 6735 -4990 6755
rect -4970 6735 -4950 6755
rect -4930 6735 -4910 6755
rect -4890 6735 -4870 6755
rect -4850 6735 -4830 6755
rect -4810 6735 -4790 6755
rect -4770 6735 -4750 6755
rect -4730 6735 -4710 6755
rect -4690 6735 -4670 6755
rect -4650 6735 -4630 6755
rect -4610 6735 -4590 6755
rect -4570 6735 -4550 6755
rect -4530 6735 -4510 6755
rect -4490 6735 -4470 6755
rect -4450 6735 -4430 6755
rect -4410 6735 -4390 6755
rect -4370 6735 -4350 6755
rect -4330 6735 -4310 6755
rect -4290 6735 -4270 6755
rect -4250 6735 -4230 6755
rect -4210 6735 -4190 6755
rect -4170 6735 -4150 6755
rect -4130 6735 -4110 6755
rect -4090 6735 -4070 6755
rect -4050 6735 -4030 6755
rect -4010 6735 -3990 6755
rect -3970 6735 -3950 6755
rect -3930 6735 -3910 6755
rect -3890 6735 -3870 6755
rect -3850 6735 -3830 6755
rect -3810 6735 -3790 6755
rect -3770 6735 -3750 6755
rect -3730 6735 -3710 6755
rect -3690 6735 -3670 6755
rect -3650 6735 -3630 6755
rect -3610 6735 -3590 6755
rect -3570 6735 -3550 6755
rect -3530 6735 -3510 6755
rect -3490 6735 -3470 6755
rect -3450 6735 -3430 6755
rect -3410 6735 -3390 6755
rect -3370 6735 -3350 6755
rect -3330 6735 -3310 6755
rect -3290 6735 -3270 6755
rect -3250 6735 -3230 6755
rect -3210 6735 -3190 6755
rect -5650 6653 -5630 6673
rect -5610 6653 -5590 6673
rect -5570 6653 -5550 6673
rect -5530 6653 -5510 6673
rect -5490 6653 -5470 6673
rect -5450 6653 -5430 6673
rect -5410 6653 -5390 6673
rect -5370 6653 -5350 6673
rect -5330 6653 -5310 6673
rect -5290 6653 -5270 6673
rect -5250 6653 -5230 6673
rect -5210 6653 -5190 6673
rect -5170 6653 -5150 6673
rect -5130 6653 -5110 6673
rect -5090 6653 -5070 6673
rect -5050 6653 -5030 6673
rect -5010 6653 -4990 6673
rect -4970 6653 -4950 6673
rect -4930 6653 -4910 6673
rect -4890 6653 -4870 6673
rect -4850 6653 -4830 6673
rect -4810 6653 -4790 6673
rect -4770 6653 -4750 6673
rect -4730 6653 -4710 6673
rect -4690 6653 -4670 6673
rect -4650 6653 -4630 6673
rect -4610 6653 -4590 6673
rect -4570 6653 -4550 6673
rect -4530 6653 -4510 6673
rect -4490 6653 -4470 6673
rect -4450 6653 -4430 6673
rect -4410 6653 -4390 6673
rect -4370 6653 -4350 6673
rect -4330 6653 -4310 6673
rect -4290 6653 -4270 6673
rect -4250 6653 -4230 6673
rect -4210 6653 -4190 6673
rect -4170 6653 -4150 6673
rect -4130 6653 -4110 6673
rect -4090 6653 -4070 6673
rect -4050 6653 -4030 6673
rect -4010 6653 -3990 6673
rect -3970 6653 -3950 6673
rect -3930 6653 -3910 6673
rect -3890 6653 -3870 6673
rect -3850 6653 -3830 6673
rect -3810 6653 -3790 6673
rect -3770 6653 -3750 6673
rect -3730 6653 -3710 6673
rect -3690 6653 -3670 6673
rect -3650 6653 -3630 6673
rect -3610 6653 -3590 6673
rect -3570 6653 -3550 6673
rect -3530 6653 -3510 6673
rect -3490 6653 -3470 6673
rect -3450 6653 -3430 6673
rect -3410 6653 -3390 6673
rect -3370 6653 -3350 6673
rect -3330 6653 -3310 6673
rect -3290 6653 -3270 6673
rect -3250 6653 -3230 6673
rect -3210 6653 -3190 6673
rect -5650 6571 -5630 6591
rect -5610 6571 -5590 6591
rect -5570 6571 -5550 6591
rect -5530 6571 -5510 6591
rect -5490 6571 -5470 6591
rect -5450 6571 -5430 6591
rect -5410 6571 -5390 6591
rect -5370 6571 -5350 6591
rect -5330 6571 -5310 6591
rect -5290 6571 -5270 6591
rect -5250 6571 -5230 6591
rect -5210 6571 -5190 6591
rect -5170 6571 -5150 6591
rect -5130 6571 -5110 6591
rect -5090 6571 -5070 6591
rect -5050 6571 -5030 6591
rect -5010 6571 -4990 6591
rect -4970 6571 -4950 6591
rect -4930 6571 -4910 6591
rect -4890 6571 -4870 6591
rect -4850 6571 -4830 6591
rect -4810 6571 -4790 6591
rect -4770 6571 -4750 6591
rect -4730 6571 -4710 6591
rect -4690 6571 -4670 6591
rect -4650 6571 -4630 6591
rect -4610 6571 -4590 6591
rect -4570 6571 -4550 6591
rect -4530 6571 -4510 6591
rect -4490 6571 -4470 6591
rect -4450 6571 -4430 6591
rect -4410 6571 -4390 6591
rect -4370 6571 -4350 6591
rect -4330 6571 -4310 6591
rect -4290 6571 -4270 6591
rect -4250 6571 -4230 6591
rect -4210 6571 -4190 6591
rect -4170 6571 -4150 6591
rect -4130 6571 -4110 6591
rect -4090 6571 -4070 6591
rect -4050 6571 -4030 6591
rect -4010 6571 -3990 6591
rect -3970 6571 -3950 6591
rect -3930 6571 -3910 6591
rect -3890 6571 -3870 6591
rect -3850 6571 -3830 6591
rect -3810 6571 -3790 6591
rect -3770 6571 -3750 6591
rect -3730 6571 -3710 6591
rect -3690 6571 -3670 6591
rect -3650 6571 -3630 6591
rect -3610 6571 -3590 6591
rect -3570 6571 -3550 6591
rect -3530 6571 -3510 6591
rect -3490 6571 -3470 6591
rect -3450 6571 -3430 6591
rect -3410 6571 -3390 6591
rect -3370 6571 -3350 6591
rect -3330 6571 -3310 6591
rect -3290 6571 -3270 6591
rect -3250 6571 -3230 6591
rect -3210 6571 -3190 6591
rect -5650 6489 -5630 6509
rect -5610 6489 -5590 6509
rect -5570 6489 -5550 6509
rect -5530 6489 -5510 6509
rect -5490 6489 -5470 6509
rect -5450 6489 -5430 6509
rect -5410 6489 -5390 6509
rect -5370 6489 -5350 6509
rect -5330 6489 -5310 6509
rect -5290 6489 -5270 6509
rect -5250 6489 -5230 6509
rect -5210 6489 -5190 6509
rect -5170 6489 -5150 6509
rect -5130 6489 -5110 6509
rect -5090 6489 -5070 6509
rect -5050 6489 -5030 6509
rect -5010 6489 -4990 6509
rect -4970 6489 -4950 6509
rect -4930 6489 -4910 6509
rect -4890 6489 -4870 6509
rect -4850 6489 -4830 6509
rect -4810 6489 -4790 6509
rect -4770 6489 -4750 6509
rect -4730 6489 -4710 6509
rect -4690 6489 -4670 6509
rect -4650 6489 -4630 6509
rect -4610 6489 -4590 6509
rect -4570 6489 -4550 6509
rect -4530 6489 -4510 6509
rect -4490 6489 -4470 6509
rect -4450 6489 -4430 6509
rect -4410 6489 -4390 6509
rect -4370 6489 -4350 6509
rect -4330 6489 -4310 6509
rect -4290 6489 -4270 6509
rect -4250 6489 -4230 6509
rect -4210 6489 -4190 6509
rect -4170 6489 -4150 6509
rect -4130 6489 -4110 6509
rect -4090 6489 -4070 6509
rect -4050 6489 -4030 6509
rect -4010 6489 -3990 6509
rect -3970 6489 -3950 6509
rect -3930 6489 -3910 6509
rect -3890 6489 -3870 6509
rect -3850 6489 -3830 6509
rect -3810 6489 -3790 6509
rect -3770 6489 -3750 6509
rect -3730 6489 -3710 6509
rect -3690 6489 -3670 6509
rect -3650 6489 -3630 6509
rect -3610 6489 -3590 6509
rect -3570 6489 -3550 6509
rect -3530 6489 -3510 6509
rect -3490 6489 -3470 6509
rect -3450 6489 -3430 6509
rect -3410 6489 -3390 6509
rect -3370 6489 -3350 6509
rect -3330 6489 -3310 6509
rect -3290 6489 -3270 6509
rect -3250 6489 -3230 6509
rect -3210 6489 -3190 6509
rect -5650 6407 -5630 6427
rect -5610 6407 -5590 6427
rect -5570 6407 -5550 6427
rect -5530 6407 -5510 6427
rect -5490 6407 -5470 6427
rect -5450 6407 -5430 6427
rect -5410 6407 -5390 6427
rect -5370 6407 -5350 6427
rect -5330 6407 -5310 6427
rect -5290 6407 -5270 6427
rect -5250 6407 -5230 6427
rect -5210 6407 -5190 6427
rect -5170 6407 -5150 6427
rect -5130 6407 -5110 6427
rect -5090 6407 -5070 6427
rect -5050 6407 -5030 6427
rect -5010 6407 -4990 6427
rect -4970 6407 -4950 6427
rect -4930 6407 -4910 6427
rect -4890 6407 -4870 6427
rect -4850 6407 -4830 6427
rect -4810 6407 -4790 6427
rect -4770 6407 -4750 6427
rect -4730 6407 -4710 6427
rect -4690 6407 -4670 6427
rect -4650 6407 -4630 6427
rect -4610 6407 -4590 6427
rect -4570 6407 -4550 6427
rect -4530 6407 -4510 6427
rect -4490 6407 -4470 6427
rect -4450 6407 -4430 6427
rect -4410 6407 -4390 6427
rect -4370 6407 -4350 6427
rect -4330 6407 -4310 6427
rect -4290 6407 -4270 6427
rect -4250 6407 -4230 6427
rect -4210 6407 -4190 6427
rect -4170 6407 -4150 6427
rect -4130 6407 -4110 6427
rect -4090 6407 -4070 6427
rect -4050 6407 -4030 6427
rect -4010 6407 -3990 6427
rect -3970 6407 -3950 6427
rect -3930 6407 -3910 6427
rect -3890 6407 -3870 6427
rect -3850 6407 -3830 6427
rect -3810 6407 -3790 6427
rect -3770 6407 -3750 6427
rect -3730 6407 -3710 6427
rect -3690 6407 -3670 6427
rect -3650 6407 -3630 6427
rect -3610 6407 -3590 6427
rect -3570 6407 -3550 6427
rect -3530 6407 -3510 6427
rect -3490 6407 -3470 6427
rect -3450 6407 -3430 6427
rect -3410 6407 -3390 6427
rect -3370 6407 -3350 6427
rect -3330 6407 -3310 6427
rect -3290 6407 -3270 6427
rect -3250 6407 -3230 6427
rect -3210 6407 -3190 6427
rect -5650 6325 -5630 6345
rect -5610 6325 -5590 6345
rect -5570 6325 -5550 6345
rect -5530 6325 -5510 6345
rect -5490 6325 -5470 6345
rect -5450 6325 -5430 6345
rect -5410 6325 -5390 6345
rect -5370 6325 -5350 6345
rect -5330 6325 -5310 6345
rect -5290 6325 -5270 6345
rect -5250 6325 -5230 6345
rect -5210 6325 -5190 6345
rect -5170 6325 -5150 6345
rect -5130 6325 -5110 6345
rect -5090 6325 -5070 6345
rect -5050 6325 -5030 6345
rect -5010 6325 -4990 6345
rect -4970 6325 -4950 6345
rect -4930 6325 -4910 6345
rect -4890 6325 -4870 6345
rect -4850 6325 -4830 6345
rect -4810 6325 -4790 6345
rect -4770 6325 -4750 6345
rect -4730 6325 -4710 6345
rect -4690 6325 -4670 6345
rect -4650 6325 -4630 6345
rect -4610 6325 -4590 6345
rect -4570 6325 -4550 6345
rect -4530 6325 -4510 6345
rect -4490 6325 -4470 6345
rect -4450 6325 -4430 6345
rect -4410 6325 -4390 6345
rect -4370 6325 -4350 6345
rect -4330 6325 -4310 6345
rect -4290 6325 -4270 6345
rect -4250 6325 -4230 6345
rect -4210 6325 -4190 6345
rect -4170 6325 -4150 6345
rect -4130 6325 -4110 6345
rect -4090 6325 -4070 6345
rect -4050 6325 -4030 6345
rect -4010 6325 -3990 6345
rect -3970 6325 -3950 6345
rect -3930 6325 -3910 6345
rect -3890 6325 -3870 6345
rect -3850 6325 -3830 6345
rect -3810 6325 -3790 6345
rect -3770 6325 -3750 6345
rect -3730 6325 -3710 6345
rect -3690 6325 -3670 6345
rect -3650 6325 -3630 6345
rect -3610 6325 -3590 6345
rect -3570 6325 -3550 6345
rect -3530 6325 -3510 6345
rect -3490 6325 -3470 6345
rect -3450 6325 -3430 6345
rect -3410 6325 -3390 6345
rect -3370 6325 -3350 6345
rect -3330 6325 -3310 6345
rect -3290 6325 -3270 6345
rect -3250 6325 -3230 6345
rect -3210 6325 -3190 6345
rect -1950 8457 -1930 8477
rect -1910 8457 -1890 8477
rect -1870 8457 -1850 8477
rect -1830 8457 -1810 8477
rect -1790 8457 -1770 8477
rect -1750 8457 -1730 8477
rect -1710 8457 -1690 8477
rect -1670 8457 -1650 8477
rect -1630 8457 -1610 8477
rect -1590 8457 -1570 8477
rect -1550 8457 -1530 8477
rect -1510 8457 -1490 8477
rect -1470 8457 -1450 8477
rect -1430 8457 -1410 8477
rect -1390 8457 -1370 8477
rect -1350 8457 -1330 8477
rect -1310 8457 -1290 8477
rect -1270 8457 -1250 8477
rect -1230 8457 -1210 8477
rect -1190 8457 -1170 8477
rect -1150 8457 -1130 8477
rect -1110 8457 -1090 8477
rect -1070 8457 -1050 8477
rect -1030 8457 -1010 8477
rect -990 8457 -970 8477
rect -950 8457 -930 8477
rect -910 8457 -890 8477
rect -870 8457 -850 8477
rect -830 8457 -810 8477
rect -790 8457 -770 8477
rect -750 8457 -730 8477
rect -710 8457 -690 8477
rect -670 8457 -650 8477
rect -630 8457 -610 8477
rect -590 8457 -570 8477
rect -550 8457 -530 8477
rect -510 8457 -490 8477
rect -470 8457 -450 8477
rect -430 8457 -410 8477
rect -390 8457 -370 8477
rect -350 8457 -330 8477
rect -310 8457 -290 8477
rect -270 8457 -250 8477
rect -230 8457 -210 8477
rect -190 8457 -170 8477
rect -150 8457 -130 8477
rect -110 8457 -90 8477
rect -70 8457 -50 8477
rect -30 8457 -10 8477
rect 10 8457 30 8477
rect 50 8457 70 8477
rect 90 8457 110 8477
rect 130 8457 150 8477
rect 170 8457 190 8477
rect 210 8457 230 8477
rect 250 8457 270 8477
rect 290 8457 310 8477
rect 330 8457 350 8477
rect 370 8457 390 8477
rect 410 8457 430 8477
rect 450 8457 470 8477
rect 490 8457 510 8477
rect -1950 8375 -1930 8395
rect -1910 8375 -1890 8395
rect -1870 8375 -1850 8395
rect -1830 8375 -1810 8395
rect -1790 8375 -1770 8395
rect -1750 8375 -1730 8395
rect -1710 8375 -1690 8395
rect -1670 8375 -1650 8395
rect -1630 8375 -1610 8395
rect -1590 8375 -1570 8395
rect -1550 8375 -1530 8395
rect -1510 8375 -1490 8395
rect -1470 8375 -1450 8395
rect -1430 8375 -1410 8395
rect -1390 8375 -1370 8395
rect -1350 8375 -1330 8395
rect -1310 8375 -1290 8395
rect -1270 8375 -1250 8395
rect -1230 8375 -1210 8395
rect -1190 8375 -1170 8395
rect -1150 8375 -1130 8395
rect -1110 8375 -1090 8395
rect -1070 8375 -1050 8395
rect -1030 8375 -1010 8395
rect -990 8375 -970 8395
rect -950 8375 -930 8395
rect -910 8375 -890 8395
rect -870 8375 -850 8395
rect -830 8375 -810 8395
rect -790 8375 -770 8395
rect -750 8375 -730 8395
rect -710 8375 -690 8395
rect -670 8375 -650 8395
rect -630 8375 -610 8395
rect -590 8375 -570 8395
rect -550 8375 -530 8395
rect -510 8375 -490 8395
rect -470 8375 -450 8395
rect -430 8375 -410 8395
rect -390 8375 -370 8395
rect -350 8375 -330 8395
rect -310 8375 -290 8395
rect -270 8375 -250 8395
rect -230 8375 -210 8395
rect -190 8375 -170 8395
rect -150 8375 -130 8395
rect -110 8375 -90 8395
rect -70 8375 -50 8395
rect -30 8375 -10 8395
rect 10 8375 30 8395
rect 50 8375 70 8395
rect 90 8375 110 8395
rect 130 8375 150 8395
rect 170 8375 190 8395
rect 210 8375 230 8395
rect 250 8375 270 8395
rect 290 8375 310 8395
rect 330 8375 350 8395
rect 370 8375 390 8395
rect 410 8375 430 8395
rect 450 8375 470 8395
rect 490 8375 510 8395
rect -1950 8293 -1930 8313
rect -1910 8293 -1890 8313
rect -1870 8293 -1850 8313
rect -1830 8293 -1810 8313
rect -1790 8293 -1770 8313
rect -1750 8293 -1730 8313
rect -1710 8293 -1690 8313
rect -1670 8293 -1650 8313
rect -1630 8293 -1610 8313
rect -1590 8293 -1570 8313
rect -1550 8293 -1530 8313
rect -1510 8293 -1490 8313
rect -1470 8293 -1450 8313
rect -1430 8293 -1410 8313
rect -1390 8293 -1370 8313
rect -1350 8293 -1330 8313
rect -1310 8293 -1290 8313
rect -1270 8293 -1250 8313
rect -1230 8293 -1210 8313
rect -1190 8293 -1170 8313
rect -1150 8293 -1130 8313
rect -1110 8293 -1090 8313
rect -1070 8293 -1050 8313
rect -1030 8293 -1010 8313
rect -990 8293 -970 8313
rect -950 8293 -930 8313
rect -910 8293 -890 8313
rect -870 8293 -850 8313
rect -830 8293 -810 8313
rect -790 8293 -770 8313
rect -750 8293 -730 8313
rect -710 8293 -690 8313
rect -670 8293 -650 8313
rect -630 8293 -610 8313
rect -590 8293 -570 8313
rect -550 8293 -530 8313
rect -510 8293 -490 8313
rect -470 8293 -450 8313
rect -430 8293 -410 8313
rect -390 8293 -370 8313
rect -350 8293 -330 8313
rect -310 8293 -290 8313
rect -270 8293 -250 8313
rect -230 8293 -210 8313
rect -190 8293 -170 8313
rect -150 8293 -130 8313
rect -110 8293 -90 8313
rect -70 8293 -50 8313
rect -30 8293 -10 8313
rect 10 8293 30 8313
rect 50 8293 70 8313
rect 90 8293 110 8313
rect 130 8293 150 8313
rect 170 8293 190 8313
rect 210 8293 230 8313
rect 250 8293 270 8313
rect 290 8293 310 8313
rect 330 8293 350 8313
rect 370 8293 390 8313
rect 410 8293 430 8313
rect 450 8293 470 8313
rect 490 8293 510 8313
rect -1950 8211 -1930 8231
rect -1910 8211 -1890 8231
rect -1870 8211 -1850 8231
rect -1830 8211 -1810 8231
rect -1790 8211 -1770 8231
rect -1750 8211 -1730 8231
rect -1710 8211 -1690 8231
rect -1670 8211 -1650 8231
rect -1630 8211 -1610 8231
rect -1590 8211 -1570 8231
rect -1550 8211 -1530 8231
rect -1510 8211 -1490 8231
rect -1470 8211 -1450 8231
rect -1430 8211 -1410 8231
rect -1390 8211 -1370 8231
rect -1350 8211 -1330 8231
rect -1310 8211 -1290 8231
rect -1270 8211 -1250 8231
rect -1230 8211 -1210 8231
rect -1190 8211 -1170 8231
rect -1150 8211 -1130 8231
rect -1110 8211 -1090 8231
rect -1070 8211 -1050 8231
rect -1030 8211 -1010 8231
rect -990 8211 -970 8231
rect -950 8211 -930 8231
rect -910 8211 -890 8231
rect -870 8211 -850 8231
rect -830 8211 -810 8231
rect -790 8211 -770 8231
rect -750 8211 -730 8231
rect -710 8211 -690 8231
rect -670 8211 -650 8231
rect -630 8211 -610 8231
rect -590 8211 -570 8231
rect -550 8211 -530 8231
rect -510 8211 -490 8231
rect -470 8211 -450 8231
rect -430 8211 -410 8231
rect -390 8211 -370 8231
rect -350 8211 -330 8231
rect -310 8211 -290 8231
rect -270 8211 -250 8231
rect -230 8211 -210 8231
rect -190 8211 -170 8231
rect -150 8211 -130 8231
rect -110 8211 -90 8231
rect -70 8211 -50 8231
rect -30 8211 -10 8231
rect 10 8211 30 8231
rect 50 8211 70 8231
rect 90 8211 110 8231
rect 130 8211 150 8231
rect 170 8211 190 8231
rect 210 8211 230 8231
rect 250 8211 270 8231
rect 290 8211 310 8231
rect 330 8211 350 8231
rect 370 8211 390 8231
rect 410 8211 430 8231
rect 450 8211 470 8231
rect 490 8211 510 8231
rect -1950 8129 -1930 8149
rect -1910 8129 -1890 8149
rect -1870 8129 -1850 8149
rect -1830 8129 -1810 8149
rect -1790 8129 -1770 8149
rect -1750 8129 -1730 8149
rect -1710 8129 -1690 8149
rect -1670 8129 -1650 8149
rect -1630 8129 -1610 8149
rect -1590 8129 -1570 8149
rect -1550 8129 -1530 8149
rect -1510 8129 -1490 8149
rect -1470 8129 -1450 8149
rect -1430 8129 -1410 8149
rect -1390 8129 -1370 8149
rect -1350 8129 -1330 8149
rect -1310 8129 -1290 8149
rect -1270 8129 -1250 8149
rect -1230 8129 -1210 8149
rect -1190 8129 -1170 8149
rect -1150 8129 -1130 8149
rect -1110 8129 -1090 8149
rect -1070 8129 -1050 8149
rect -1030 8129 -1010 8149
rect -990 8129 -970 8149
rect -950 8129 -930 8149
rect -910 8129 -890 8149
rect -870 8129 -850 8149
rect -830 8129 -810 8149
rect -790 8129 -770 8149
rect -750 8129 -730 8149
rect -710 8129 -690 8149
rect -670 8129 -650 8149
rect -630 8129 -610 8149
rect -590 8129 -570 8149
rect -550 8129 -530 8149
rect -510 8129 -490 8149
rect -470 8129 -450 8149
rect -430 8129 -410 8149
rect -390 8129 -370 8149
rect -350 8129 -330 8149
rect -310 8129 -290 8149
rect -270 8129 -250 8149
rect -230 8129 -210 8149
rect -190 8129 -170 8149
rect -150 8129 -130 8149
rect -110 8129 -90 8149
rect -70 8129 -50 8149
rect -30 8129 -10 8149
rect 10 8129 30 8149
rect 50 8129 70 8149
rect 90 8129 110 8149
rect 130 8129 150 8149
rect 170 8129 190 8149
rect 210 8129 230 8149
rect 250 8129 270 8149
rect 290 8129 310 8149
rect 330 8129 350 8149
rect 370 8129 390 8149
rect 410 8129 430 8149
rect 450 8129 470 8149
rect 490 8129 510 8149
rect -1950 8047 -1930 8067
rect -1910 8047 -1890 8067
rect -1870 8047 -1850 8067
rect -1830 8047 -1810 8067
rect -1790 8047 -1770 8067
rect -1750 8047 -1730 8067
rect -1710 8047 -1690 8067
rect -1670 8047 -1650 8067
rect -1630 8047 -1610 8067
rect -1590 8047 -1570 8067
rect -1550 8047 -1530 8067
rect -1510 8047 -1490 8067
rect -1470 8047 -1450 8067
rect -1430 8047 -1410 8067
rect -1390 8047 -1370 8067
rect -1350 8047 -1330 8067
rect -1310 8047 -1290 8067
rect -1270 8047 -1250 8067
rect -1230 8047 -1210 8067
rect -1190 8047 -1170 8067
rect -1150 8047 -1130 8067
rect -1110 8047 -1090 8067
rect -1070 8047 -1050 8067
rect -1030 8047 -1010 8067
rect -990 8047 -970 8067
rect -950 8047 -930 8067
rect -910 8047 -890 8067
rect -870 8047 -850 8067
rect -830 8047 -810 8067
rect -790 8047 -770 8067
rect -750 8047 -730 8067
rect -710 8047 -690 8067
rect -670 8047 -650 8067
rect -630 8047 -610 8067
rect -590 8047 -570 8067
rect -550 8047 -530 8067
rect -510 8047 -490 8067
rect -470 8047 -450 8067
rect -430 8047 -410 8067
rect -390 8047 -370 8067
rect -350 8047 -330 8067
rect -310 8047 -290 8067
rect -270 8047 -250 8067
rect -230 8047 -210 8067
rect -190 8047 -170 8067
rect -150 8047 -130 8067
rect -110 8047 -90 8067
rect -70 8047 -50 8067
rect -30 8047 -10 8067
rect 10 8047 30 8067
rect 50 8047 70 8067
rect 90 8047 110 8067
rect 130 8047 150 8067
rect 170 8047 190 8067
rect 210 8047 230 8067
rect 250 8047 270 8067
rect 290 8047 310 8067
rect 330 8047 350 8067
rect 370 8047 390 8067
rect 410 8047 430 8067
rect 450 8047 470 8067
rect 490 8047 510 8067
rect -1950 7965 -1930 7985
rect -1910 7965 -1890 7985
rect -1870 7965 -1850 7985
rect -1830 7965 -1810 7985
rect -1790 7965 -1770 7985
rect -1750 7965 -1730 7985
rect -1710 7965 -1690 7985
rect -1670 7965 -1650 7985
rect -1630 7965 -1610 7985
rect -1590 7965 -1570 7985
rect -1550 7965 -1530 7985
rect -1510 7965 -1490 7985
rect -1470 7965 -1450 7985
rect -1430 7965 -1410 7985
rect -1390 7965 -1370 7985
rect -1350 7965 -1330 7985
rect -1310 7965 -1290 7985
rect -1270 7965 -1250 7985
rect -1230 7965 -1210 7985
rect -1190 7965 -1170 7985
rect -1150 7965 -1130 7985
rect -1110 7965 -1090 7985
rect -1070 7965 -1050 7985
rect -1030 7965 -1010 7985
rect -990 7965 -970 7985
rect -950 7965 -930 7985
rect -910 7965 -890 7985
rect -870 7965 -850 7985
rect -830 7965 -810 7985
rect -790 7965 -770 7985
rect -750 7965 -730 7985
rect -710 7965 -690 7985
rect -670 7965 -650 7985
rect -630 7965 -610 7985
rect -590 7965 -570 7985
rect -550 7965 -530 7985
rect -510 7965 -490 7985
rect -470 7965 -450 7985
rect -430 7965 -410 7985
rect -390 7965 -370 7985
rect -350 7965 -330 7985
rect -310 7965 -290 7985
rect -270 7965 -250 7985
rect -230 7965 -210 7985
rect -190 7965 -170 7985
rect -150 7965 -130 7985
rect -110 7965 -90 7985
rect -70 7965 -50 7985
rect -30 7965 -10 7985
rect 10 7965 30 7985
rect 50 7965 70 7985
rect 90 7965 110 7985
rect 130 7965 150 7985
rect 170 7965 190 7985
rect 210 7965 230 7985
rect 250 7965 270 7985
rect 290 7965 310 7985
rect 330 7965 350 7985
rect 370 7965 390 7985
rect 410 7965 430 7985
rect 450 7965 470 7985
rect 490 7965 510 7985
rect -1950 7883 -1930 7903
rect -1910 7883 -1890 7903
rect -1870 7883 -1850 7903
rect -1830 7883 -1810 7903
rect -1790 7883 -1770 7903
rect -1750 7883 -1730 7903
rect -1710 7883 -1690 7903
rect -1670 7883 -1650 7903
rect -1630 7883 -1610 7903
rect -1590 7883 -1570 7903
rect -1550 7883 -1530 7903
rect -1510 7883 -1490 7903
rect -1470 7883 -1450 7903
rect -1430 7883 -1410 7903
rect -1390 7883 -1370 7903
rect -1350 7883 -1330 7903
rect -1310 7883 -1290 7903
rect -1270 7883 -1250 7903
rect -1230 7883 -1210 7903
rect -1190 7883 -1170 7903
rect -1150 7883 -1130 7903
rect -1110 7883 -1090 7903
rect -1070 7883 -1050 7903
rect -1030 7883 -1010 7903
rect -990 7883 -970 7903
rect -950 7883 -930 7903
rect -910 7883 -890 7903
rect -870 7883 -850 7903
rect -830 7883 -810 7903
rect -790 7883 -770 7903
rect -750 7883 -730 7903
rect -710 7883 -690 7903
rect -670 7883 -650 7903
rect -630 7883 -610 7903
rect -590 7883 -570 7903
rect -550 7883 -530 7903
rect -510 7883 -490 7903
rect -470 7883 -450 7903
rect -430 7883 -410 7903
rect -390 7883 -370 7903
rect -350 7883 -330 7903
rect -310 7883 -290 7903
rect -270 7883 -250 7903
rect -230 7883 -210 7903
rect -190 7883 -170 7903
rect -150 7883 -130 7903
rect -110 7883 -90 7903
rect -70 7883 -50 7903
rect -30 7883 -10 7903
rect 10 7883 30 7903
rect 50 7883 70 7903
rect 90 7883 110 7903
rect 130 7883 150 7903
rect 170 7883 190 7903
rect 210 7883 230 7903
rect 250 7883 270 7903
rect 290 7883 310 7903
rect 330 7883 350 7903
rect 370 7883 390 7903
rect 410 7883 430 7903
rect 450 7883 470 7903
rect 490 7883 510 7903
rect -1950 7801 -1930 7821
rect -1910 7801 -1890 7821
rect -1870 7801 -1850 7821
rect -1830 7801 -1810 7821
rect -1790 7801 -1770 7821
rect -1750 7801 -1730 7821
rect -1710 7801 -1690 7821
rect -1670 7801 -1650 7821
rect -1630 7801 -1610 7821
rect -1590 7801 -1570 7821
rect -1550 7801 -1530 7821
rect -1510 7801 -1490 7821
rect -1470 7801 -1450 7821
rect -1430 7801 -1410 7821
rect -1390 7801 -1370 7821
rect -1350 7801 -1330 7821
rect -1310 7801 -1290 7821
rect -1270 7801 -1250 7821
rect -1230 7801 -1210 7821
rect -1190 7801 -1170 7821
rect -1150 7801 -1130 7821
rect -1110 7801 -1090 7821
rect -1070 7801 -1050 7821
rect -1030 7801 -1010 7821
rect -990 7801 -970 7821
rect -950 7801 -930 7821
rect -910 7801 -890 7821
rect -870 7801 -850 7821
rect -830 7801 -810 7821
rect -790 7801 -770 7821
rect -750 7801 -730 7821
rect -710 7801 -690 7821
rect -670 7801 -650 7821
rect -630 7801 -610 7821
rect -590 7801 -570 7821
rect -550 7801 -530 7821
rect -510 7801 -490 7821
rect -470 7801 -450 7821
rect -430 7801 -410 7821
rect -390 7801 -370 7821
rect -350 7801 -330 7821
rect -310 7801 -290 7821
rect -270 7801 -250 7821
rect -230 7801 -210 7821
rect -190 7801 -170 7821
rect -150 7801 -130 7821
rect -110 7801 -90 7821
rect -70 7801 -50 7821
rect -30 7801 -10 7821
rect 10 7801 30 7821
rect 50 7801 70 7821
rect 90 7801 110 7821
rect 130 7801 150 7821
rect 170 7801 190 7821
rect 210 7801 230 7821
rect 250 7801 270 7821
rect 290 7801 310 7821
rect 330 7801 350 7821
rect 370 7801 390 7821
rect 410 7801 430 7821
rect 450 7801 470 7821
rect 490 7801 510 7821
rect -1950 7719 -1930 7739
rect -1910 7719 -1890 7739
rect -1870 7719 -1850 7739
rect -1830 7719 -1810 7739
rect -1790 7719 -1770 7739
rect -1750 7719 -1730 7739
rect -1710 7719 -1690 7739
rect -1670 7719 -1650 7739
rect -1630 7719 -1610 7739
rect -1590 7719 -1570 7739
rect -1550 7719 -1530 7739
rect -1510 7719 -1490 7739
rect -1470 7719 -1450 7739
rect -1430 7719 -1410 7739
rect -1390 7719 -1370 7739
rect -1350 7719 -1330 7739
rect -1310 7719 -1290 7739
rect -1270 7719 -1250 7739
rect -1230 7719 -1210 7739
rect -1190 7719 -1170 7739
rect -1150 7719 -1130 7739
rect -1110 7719 -1090 7739
rect -1070 7719 -1050 7739
rect -1030 7719 -1010 7739
rect -990 7719 -970 7739
rect -950 7719 -930 7739
rect -910 7719 -890 7739
rect -870 7719 -850 7739
rect -830 7719 -810 7739
rect -790 7719 -770 7739
rect -750 7719 -730 7739
rect -710 7719 -690 7739
rect -670 7719 -650 7739
rect -630 7719 -610 7739
rect -590 7719 -570 7739
rect -550 7719 -530 7739
rect -510 7719 -490 7739
rect -470 7719 -450 7739
rect -430 7719 -410 7739
rect -390 7719 -370 7739
rect -350 7719 -330 7739
rect -310 7719 -290 7739
rect -270 7719 -250 7739
rect -230 7719 -210 7739
rect -190 7719 -170 7739
rect -150 7719 -130 7739
rect -110 7719 -90 7739
rect -70 7719 -50 7739
rect -30 7719 -10 7739
rect 10 7719 30 7739
rect 50 7719 70 7739
rect 90 7719 110 7739
rect 130 7719 150 7739
rect 170 7719 190 7739
rect 210 7719 230 7739
rect 250 7719 270 7739
rect 290 7719 310 7739
rect 330 7719 350 7739
rect 370 7719 390 7739
rect 410 7719 430 7739
rect 450 7719 470 7739
rect 490 7719 510 7739
rect -1950 7637 -1930 7657
rect -1910 7637 -1890 7657
rect -1870 7637 -1850 7657
rect -1830 7637 -1810 7657
rect -1790 7637 -1770 7657
rect -1750 7637 -1730 7657
rect -1710 7637 -1690 7657
rect -1670 7637 -1650 7657
rect -1630 7637 -1610 7657
rect -1590 7637 -1570 7657
rect -1550 7637 -1530 7657
rect -1510 7637 -1490 7657
rect -1470 7637 -1450 7657
rect -1430 7637 -1410 7657
rect -1390 7637 -1370 7657
rect -1350 7637 -1330 7657
rect -1310 7637 -1290 7657
rect -1270 7637 -1250 7657
rect -1230 7637 -1210 7657
rect -1190 7637 -1170 7657
rect -1150 7637 -1130 7657
rect -1110 7637 -1090 7657
rect -1070 7637 -1050 7657
rect -1030 7637 -1010 7657
rect -990 7637 -970 7657
rect -950 7637 -930 7657
rect -910 7637 -890 7657
rect -870 7637 -850 7657
rect -830 7637 -810 7657
rect -790 7637 -770 7657
rect -750 7637 -730 7657
rect -710 7637 -690 7657
rect -670 7637 -650 7657
rect -630 7637 -610 7657
rect -590 7637 -570 7657
rect -550 7637 -530 7657
rect -510 7637 -490 7657
rect -470 7637 -450 7657
rect -430 7637 -410 7657
rect -390 7637 -370 7657
rect -350 7637 -330 7657
rect -310 7637 -290 7657
rect -270 7637 -250 7657
rect -230 7637 -210 7657
rect -190 7637 -170 7657
rect -150 7637 -130 7657
rect -110 7637 -90 7657
rect -70 7637 -50 7657
rect -30 7637 -10 7657
rect 10 7637 30 7657
rect 50 7637 70 7657
rect 90 7637 110 7657
rect 130 7637 150 7657
rect 170 7637 190 7657
rect 210 7637 230 7657
rect 250 7637 270 7657
rect 290 7637 310 7657
rect 330 7637 350 7657
rect 370 7637 390 7657
rect 410 7637 430 7657
rect 450 7637 470 7657
rect 490 7637 510 7657
rect -1950 7555 -1930 7575
rect -1910 7555 -1890 7575
rect -1870 7555 -1850 7575
rect -1830 7555 -1810 7575
rect -1790 7555 -1770 7575
rect -1750 7555 -1730 7575
rect -1710 7555 -1690 7575
rect -1670 7555 -1650 7575
rect -1630 7555 -1610 7575
rect -1590 7555 -1570 7575
rect -1550 7555 -1530 7575
rect -1510 7555 -1490 7575
rect -1470 7555 -1450 7575
rect -1430 7555 -1410 7575
rect -1390 7555 -1370 7575
rect -1350 7555 -1330 7575
rect -1310 7555 -1290 7575
rect -1270 7555 -1250 7575
rect -1230 7555 -1210 7575
rect -1190 7555 -1170 7575
rect -1150 7555 -1130 7575
rect -1110 7555 -1090 7575
rect -1070 7555 -1050 7575
rect -1030 7555 -1010 7575
rect -990 7555 -970 7575
rect -950 7555 -930 7575
rect -910 7555 -890 7575
rect -870 7555 -850 7575
rect -830 7555 -810 7575
rect -790 7555 -770 7575
rect -750 7555 -730 7575
rect -710 7555 -690 7575
rect -670 7555 -650 7575
rect -630 7555 -610 7575
rect -590 7555 -570 7575
rect -550 7555 -530 7575
rect -510 7555 -490 7575
rect -470 7555 -450 7575
rect -430 7555 -410 7575
rect -390 7555 -370 7575
rect -350 7555 -330 7575
rect -310 7555 -290 7575
rect -270 7555 -250 7575
rect -230 7555 -210 7575
rect -190 7555 -170 7575
rect -150 7555 -130 7575
rect -110 7555 -90 7575
rect -70 7555 -50 7575
rect -30 7555 -10 7575
rect 10 7555 30 7575
rect 50 7555 70 7575
rect 90 7555 110 7575
rect 130 7555 150 7575
rect 170 7555 190 7575
rect 210 7555 230 7575
rect 250 7555 270 7575
rect 290 7555 310 7575
rect 330 7555 350 7575
rect 370 7555 390 7575
rect 410 7555 430 7575
rect 450 7555 470 7575
rect 490 7555 510 7575
rect -1950 7473 -1930 7493
rect -1910 7473 -1890 7493
rect -1870 7473 -1850 7493
rect -1830 7473 -1810 7493
rect -1790 7473 -1770 7493
rect -1750 7473 -1730 7493
rect -1710 7473 -1690 7493
rect -1670 7473 -1650 7493
rect -1630 7473 -1610 7493
rect -1590 7473 -1570 7493
rect -1550 7473 -1530 7493
rect -1510 7473 -1490 7493
rect -1470 7473 -1450 7493
rect -1430 7473 -1410 7493
rect -1390 7473 -1370 7493
rect -1350 7473 -1330 7493
rect -1310 7473 -1290 7493
rect -1270 7473 -1250 7493
rect -1230 7473 -1210 7493
rect -1190 7473 -1170 7493
rect -1150 7473 -1130 7493
rect -1110 7473 -1090 7493
rect -1070 7473 -1050 7493
rect -1030 7473 -1010 7493
rect -990 7473 -970 7493
rect -950 7473 -930 7493
rect -910 7473 -890 7493
rect -870 7473 -850 7493
rect -830 7473 -810 7493
rect -790 7473 -770 7493
rect -750 7473 -730 7493
rect -710 7473 -690 7493
rect -670 7473 -650 7493
rect -630 7473 -610 7493
rect -590 7473 -570 7493
rect -550 7473 -530 7493
rect -510 7473 -490 7493
rect -470 7473 -450 7493
rect -430 7473 -410 7493
rect -390 7473 -370 7493
rect -350 7473 -330 7493
rect -310 7473 -290 7493
rect -270 7473 -250 7493
rect -230 7473 -210 7493
rect -190 7473 -170 7493
rect -150 7473 -130 7493
rect -110 7473 -90 7493
rect -70 7473 -50 7493
rect -30 7473 -10 7493
rect 10 7473 30 7493
rect 50 7473 70 7493
rect 90 7473 110 7493
rect 130 7473 150 7493
rect 170 7473 190 7493
rect 210 7473 230 7493
rect 250 7473 270 7493
rect 290 7473 310 7493
rect 330 7473 350 7493
rect 370 7473 390 7493
rect 410 7473 430 7493
rect 450 7473 470 7493
rect 490 7473 510 7493
rect -1950 7391 -1930 7411
rect -1910 7391 -1890 7411
rect -1870 7391 -1850 7411
rect -1830 7391 -1810 7411
rect -1790 7391 -1770 7411
rect -1750 7391 -1730 7411
rect -1710 7391 -1690 7411
rect -1670 7391 -1650 7411
rect -1630 7391 -1610 7411
rect -1590 7391 -1570 7411
rect -1550 7391 -1530 7411
rect -1510 7391 -1490 7411
rect -1470 7391 -1450 7411
rect -1430 7391 -1410 7411
rect -1390 7391 -1370 7411
rect -1350 7391 -1330 7411
rect -1310 7391 -1290 7411
rect -1270 7391 -1250 7411
rect -1230 7391 -1210 7411
rect -1190 7391 -1170 7411
rect -1150 7391 -1130 7411
rect -1110 7391 -1090 7411
rect -1070 7391 -1050 7411
rect -1030 7391 -1010 7411
rect -990 7391 -970 7411
rect -950 7391 -930 7411
rect -910 7391 -890 7411
rect -870 7391 -850 7411
rect -830 7391 -810 7411
rect -790 7391 -770 7411
rect -750 7391 -730 7411
rect -710 7391 -690 7411
rect -670 7391 -650 7411
rect -630 7391 -610 7411
rect -590 7391 -570 7411
rect -550 7391 -530 7411
rect -510 7391 -490 7411
rect -470 7391 -450 7411
rect -430 7391 -410 7411
rect -390 7391 -370 7411
rect -350 7391 -330 7411
rect -310 7391 -290 7411
rect -270 7391 -250 7411
rect -230 7391 -210 7411
rect -190 7391 -170 7411
rect -150 7391 -130 7411
rect -110 7391 -90 7411
rect -70 7391 -50 7411
rect -30 7391 -10 7411
rect 10 7391 30 7411
rect 50 7391 70 7411
rect 90 7391 110 7411
rect 130 7391 150 7411
rect 170 7391 190 7411
rect 210 7391 230 7411
rect 250 7391 270 7411
rect 290 7391 310 7411
rect 330 7391 350 7411
rect 370 7391 390 7411
rect 410 7391 430 7411
rect 450 7391 470 7411
rect 490 7391 510 7411
rect -1950 7309 -1930 7329
rect -1910 7309 -1890 7329
rect -1870 7309 -1850 7329
rect -1830 7309 -1810 7329
rect -1790 7309 -1770 7329
rect -1750 7309 -1730 7329
rect -1710 7309 -1690 7329
rect -1670 7309 -1650 7329
rect -1630 7309 -1610 7329
rect -1590 7309 -1570 7329
rect -1550 7309 -1530 7329
rect -1510 7309 -1490 7329
rect -1470 7309 -1450 7329
rect -1430 7309 -1410 7329
rect -1390 7309 -1370 7329
rect -1350 7309 -1330 7329
rect -1310 7309 -1290 7329
rect -1270 7309 -1250 7329
rect -1230 7309 -1210 7329
rect -1190 7309 -1170 7329
rect -1150 7309 -1130 7329
rect -1110 7309 -1090 7329
rect -1070 7309 -1050 7329
rect -1030 7309 -1010 7329
rect -990 7309 -970 7329
rect -950 7309 -930 7329
rect -910 7309 -890 7329
rect -870 7309 -850 7329
rect -830 7309 -810 7329
rect -790 7309 -770 7329
rect -750 7309 -730 7329
rect -710 7309 -690 7329
rect -670 7309 -650 7329
rect -630 7309 -610 7329
rect -590 7309 -570 7329
rect -550 7309 -530 7329
rect -510 7309 -490 7329
rect -470 7309 -450 7329
rect -430 7309 -410 7329
rect -390 7309 -370 7329
rect -350 7309 -330 7329
rect -310 7309 -290 7329
rect -270 7309 -250 7329
rect -230 7309 -210 7329
rect -190 7309 -170 7329
rect -150 7309 -130 7329
rect -110 7309 -90 7329
rect -70 7309 -50 7329
rect -30 7309 -10 7329
rect 10 7309 30 7329
rect 50 7309 70 7329
rect 90 7309 110 7329
rect 130 7309 150 7329
rect 170 7309 190 7329
rect 210 7309 230 7329
rect 250 7309 270 7329
rect 290 7309 310 7329
rect 330 7309 350 7329
rect 370 7309 390 7329
rect 410 7309 430 7329
rect 450 7309 470 7329
rect 490 7309 510 7329
rect -1950 7227 -1930 7247
rect -1910 7227 -1890 7247
rect -1870 7227 -1850 7247
rect -1830 7227 -1810 7247
rect -1790 7227 -1770 7247
rect -1750 7227 -1730 7247
rect -1710 7227 -1690 7247
rect -1670 7227 -1650 7247
rect -1630 7227 -1610 7247
rect -1590 7227 -1570 7247
rect -1550 7227 -1530 7247
rect -1510 7227 -1490 7247
rect -1470 7227 -1450 7247
rect -1430 7227 -1410 7247
rect -1390 7227 -1370 7247
rect -1350 7227 -1330 7247
rect -1310 7227 -1290 7247
rect -1270 7227 -1250 7247
rect -1230 7227 -1210 7247
rect -1190 7227 -1170 7247
rect -1150 7227 -1130 7247
rect -1110 7227 -1090 7247
rect -1070 7227 -1050 7247
rect -1030 7227 -1010 7247
rect -990 7227 -970 7247
rect -950 7227 -930 7247
rect -910 7227 -890 7247
rect -870 7227 -850 7247
rect -830 7227 -810 7247
rect -790 7227 -770 7247
rect -750 7227 -730 7247
rect -710 7227 -690 7247
rect -670 7227 -650 7247
rect -630 7227 -610 7247
rect -590 7227 -570 7247
rect -550 7227 -530 7247
rect -510 7227 -490 7247
rect -470 7227 -450 7247
rect -430 7227 -410 7247
rect -390 7227 -370 7247
rect -350 7227 -330 7247
rect -310 7227 -290 7247
rect -270 7227 -250 7247
rect -230 7227 -210 7247
rect -190 7227 -170 7247
rect -150 7227 -130 7247
rect -110 7227 -90 7247
rect -70 7227 -50 7247
rect -30 7227 -10 7247
rect 10 7227 30 7247
rect 50 7227 70 7247
rect 90 7227 110 7247
rect 130 7227 150 7247
rect 170 7227 190 7247
rect 210 7227 230 7247
rect 250 7227 270 7247
rect 290 7227 310 7247
rect 330 7227 350 7247
rect 370 7227 390 7247
rect 410 7227 430 7247
rect 450 7227 470 7247
rect 490 7227 510 7247
rect -1950 7145 -1930 7165
rect -1910 7145 -1890 7165
rect -1870 7145 -1850 7165
rect -1830 7145 -1810 7165
rect -1790 7145 -1770 7165
rect -1750 7145 -1730 7165
rect -1710 7145 -1690 7165
rect -1670 7145 -1650 7165
rect -1630 7145 -1610 7165
rect -1590 7145 -1570 7165
rect -1550 7145 -1530 7165
rect -1510 7145 -1490 7165
rect -1470 7145 -1450 7165
rect -1430 7145 -1410 7165
rect -1390 7145 -1370 7165
rect -1350 7145 -1330 7165
rect -1310 7145 -1290 7165
rect -1270 7145 -1250 7165
rect -1230 7145 -1210 7165
rect -1190 7145 -1170 7165
rect -1150 7145 -1130 7165
rect -1110 7145 -1090 7165
rect -1070 7145 -1050 7165
rect -1030 7145 -1010 7165
rect -990 7145 -970 7165
rect -950 7145 -930 7165
rect -910 7145 -890 7165
rect -870 7145 -850 7165
rect -830 7145 -810 7165
rect -790 7145 -770 7165
rect -750 7145 -730 7165
rect -710 7145 -690 7165
rect -670 7145 -650 7165
rect -630 7145 -610 7165
rect -590 7145 -570 7165
rect -550 7145 -530 7165
rect -510 7145 -490 7165
rect -470 7145 -450 7165
rect -430 7145 -410 7165
rect -390 7145 -370 7165
rect -350 7145 -330 7165
rect -310 7145 -290 7165
rect -270 7145 -250 7165
rect -230 7145 -210 7165
rect -190 7145 -170 7165
rect -150 7145 -130 7165
rect -110 7145 -90 7165
rect -70 7145 -50 7165
rect -30 7145 -10 7165
rect 10 7145 30 7165
rect 50 7145 70 7165
rect 90 7145 110 7165
rect 130 7145 150 7165
rect 170 7145 190 7165
rect 210 7145 230 7165
rect 250 7145 270 7165
rect 290 7145 310 7165
rect 330 7145 350 7165
rect 370 7145 390 7165
rect 410 7145 430 7165
rect 450 7145 470 7165
rect 490 7145 510 7165
rect -1950 7063 -1930 7083
rect -1910 7063 -1890 7083
rect -1870 7063 -1850 7083
rect -1830 7063 -1810 7083
rect -1790 7063 -1770 7083
rect -1750 7063 -1730 7083
rect -1710 7063 -1690 7083
rect -1670 7063 -1650 7083
rect -1630 7063 -1610 7083
rect -1590 7063 -1570 7083
rect -1550 7063 -1530 7083
rect -1510 7063 -1490 7083
rect -1470 7063 -1450 7083
rect -1430 7063 -1410 7083
rect -1390 7063 -1370 7083
rect -1350 7063 -1330 7083
rect -1310 7063 -1290 7083
rect -1270 7063 -1250 7083
rect -1230 7063 -1210 7083
rect -1190 7063 -1170 7083
rect -1150 7063 -1130 7083
rect -1110 7063 -1090 7083
rect -1070 7063 -1050 7083
rect -1030 7063 -1010 7083
rect -990 7063 -970 7083
rect -950 7063 -930 7083
rect -910 7063 -890 7083
rect -870 7063 -850 7083
rect -830 7063 -810 7083
rect -790 7063 -770 7083
rect -750 7063 -730 7083
rect -710 7063 -690 7083
rect -670 7063 -650 7083
rect -630 7063 -610 7083
rect -590 7063 -570 7083
rect -550 7063 -530 7083
rect -510 7063 -490 7083
rect -470 7063 -450 7083
rect -430 7063 -410 7083
rect -390 7063 -370 7083
rect -350 7063 -330 7083
rect -310 7063 -290 7083
rect -270 7063 -250 7083
rect -230 7063 -210 7083
rect -190 7063 -170 7083
rect -150 7063 -130 7083
rect -110 7063 -90 7083
rect -70 7063 -50 7083
rect -30 7063 -10 7083
rect 10 7063 30 7083
rect 50 7063 70 7083
rect 90 7063 110 7083
rect 130 7063 150 7083
rect 170 7063 190 7083
rect 210 7063 230 7083
rect 250 7063 270 7083
rect 290 7063 310 7083
rect 330 7063 350 7083
rect 370 7063 390 7083
rect 410 7063 430 7083
rect 450 7063 470 7083
rect 490 7063 510 7083
rect -1950 6981 -1930 7001
rect -1910 6981 -1890 7001
rect -1870 6981 -1850 7001
rect -1830 6981 -1810 7001
rect -1790 6981 -1770 7001
rect -1750 6981 -1730 7001
rect -1710 6981 -1690 7001
rect -1670 6981 -1650 7001
rect -1630 6981 -1610 7001
rect -1590 6981 -1570 7001
rect -1550 6981 -1530 7001
rect -1510 6981 -1490 7001
rect -1470 6981 -1450 7001
rect -1430 6981 -1410 7001
rect -1390 6981 -1370 7001
rect -1350 6981 -1330 7001
rect -1310 6981 -1290 7001
rect -1270 6981 -1250 7001
rect -1230 6981 -1210 7001
rect -1190 6981 -1170 7001
rect -1150 6981 -1130 7001
rect -1110 6981 -1090 7001
rect -1070 6981 -1050 7001
rect -1030 6981 -1010 7001
rect -990 6981 -970 7001
rect -950 6981 -930 7001
rect -910 6981 -890 7001
rect -870 6981 -850 7001
rect -830 6981 -810 7001
rect -790 6981 -770 7001
rect -750 6981 -730 7001
rect -710 6981 -690 7001
rect -670 6981 -650 7001
rect -630 6981 -610 7001
rect -590 6981 -570 7001
rect -550 6981 -530 7001
rect -510 6981 -490 7001
rect -470 6981 -450 7001
rect -430 6981 -410 7001
rect -390 6981 -370 7001
rect -350 6981 -330 7001
rect -310 6981 -290 7001
rect -270 6981 -250 7001
rect -230 6981 -210 7001
rect -190 6981 -170 7001
rect -150 6981 -130 7001
rect -110 6981 -90 7001
rect -70 6981 -50 7001
rect -30 6981 -10 7001
rect 10 6981 30 7001
rect 50 6981 70 7001
rect 90 6981 110 7001
rect 130 6981 150 7001
rect 170 6981 190 7001
rect 210 6981 230 7001
rect 250 6981 270 7001
rect 290 6981 310 7001
rect 330 6981 350 7001
rect 370 6981 390 7001
rect 410 6981 430 7001
rect 450 6981 470 7001
rect 490 6981 510 7001
rect -1950 6899 -1930 6919
rect -1910 6899 -1890 6919
rect -1870 6899 -1850 6919
rect -1830 6899 -1810 6919
rect -1790 6899 -1770 6919
rect -1750 6899 -1730 6919
rect -1710 6899 -1690 6919
rect -1670 6899 -1650 6919
rect -1630 6899 -1610 6919
rect -1590 6899 -1570 6919
rect -1550 6899 -1530 6919
rect -1510 6899 -1490 6919
rect -1470 6899 -1450 6919
rect -1430 6899 -1410 6919
rect -1390 6899 -1370 6919
rect -1350 6899 -1330 6919
rect -1310 6899 -1290 6919
rect -1270 6899 -1250 6919
rect -1230 6899 -1210 6919
rect -1190 6899 -1170 6919
rect -1150 6899 -1130 6919
rect -1110 6899 -1090 6919
rect -1070 6899 -1050 6919
rect -1030 6899 -1010 6919
rect -990 6899 -970 6919
rect -950 6899 -930 6919
rect -910 6899 -890 6919
rect -870 6899 -850 6919
rect -830 6899 -810 6919
rect -790 6899 -770 6919
rect -750 6899 -730 6919
rect -710 6899 -690 6919
rect -670 6899 -650 6919
rect -630 6899 -610 6919
rect -590 6899 -570 6919
rect -550 6899 -530 6919
rect -510 6899 -490 6919
rect -470 6899 -450 6919
rect -430 6899 -410 6919
rect -390 6899 -370 6919
rect -350 6899 -330 6919
rect -310 6899 -290 6919
rect -270 6899 -250 6919
rect -230 6899 -210 6919
rect -190 6899 -170 6919
rect -150 6899 -130 6919
rect -110 6899 -90 6919
rect -70 6899 -50 6919
rect -30 6899 -10 6919
rect 10 6899 30 6919
rect 50 6899 70 6919
rect 90 6899 110 6919
rect 130 6899 150 6919
rect 170 6899 190 6919
rect 210 6899 230 6919
rect 250 6899 270 6919
rect 290 6899 310 6919
rect 330 6899 350 6919
rect 370 6899 390 6919
rect 410 6899 430 6919
rect 450 6899 470 6919
rect 490 6899 510 6919
rect -1950 6817 -1930 6837
rect -1910 6817 -1890 6837
rect -1870 6817 -1850 6837
rect -1830 6817 -1810 6837
rect -1790 6817 -1770 6837
rect -1750 6817 -1730 6837
rect -1710 6817 -1690 6837
rect -1670 6817 -1650 6837
rect -1630 6817 -1610 6837
rect -1590 6817 -1570 6837
rect -1550 6817 -1530 6837
rect -1510 6817 -1490 6837
rect -1470 6817 -1450 6837
rect -1430 6817 -1410 6837
rect -1390 6817 -1370 6837
rect -1350 6817 -1330 6837
rect -1310 6817 -1290 6837
rect -1270 6817 -1250 6837
rect -1230 6817 -1210 6837
rect -1190 6817 -1170 6837
rect -1150 6817 -1130 6837
rect -1110 6817 -1090 6837
rect -1070 6817 -1050 6837
rect -1030 6817 -1010 6837
rect -990 6817 -970 6837
rect -950 6817 -930 6837
rect -910 6817 -890 6837
rect -870 6817 -850 6837
rect -830 6817 -810 6837
rect -790 6817 -770 6837
rect -750 6817 -730 6837
rect -710 6817 -690 6837
rect -670 6817 -650 6837
rect -630 6817 -610 6837
rect -590 6817 -570 6837
rect -550 6817 -530 6837
rect -510 6817 -490 6837
rect -470 6817 -450 6837
rect -430 6817 -410 6837
rect -390 6817 -370 6837
rect -350 6817 -330 6837
rect -310 6817 -290 6837
rect -270 6817 -250 6837
rect -230 6817 -210 6837
rect -190 6817 -170 6837
rect -150 6817 -130 6837
rect -110 6817 -90 6837
rect -70 6817 -50 6837
rect -30 6817 -10 6837
rect 10 6817 30 6837
rect 50 6817 70 6837
rect 90 6817 110 6837
rect 130 6817 150 6837
rect 170 6817 190 6837
rect 210 6817 230 6837
rect 250 6817 270 6837
rect 290 6817 310 6837
rect 330 6817 350 6837
rect 370 6817 390 6837
rect 410 6817 430 6837
rect 450 6817 470 6837
rect 490 6817 510 6837
rect -1950 6735 -1930 6755
rect -1910 6735 -1890 6755
rect -1870 6735 -1850 6755
rect -1830 6735 -1810 6755
rect -1790 6735 -1770 6755
rect -1750 6735 -1730 6755
rect -1710 6735 -1690 6755
rect -1670 6735 -1650 6755
rect -1630 6735 -1610 6755
rect -1590 6735 -1570 6755
rect -1550 6735 -1530 6755
rect -1510 6735 -1490 6755
rect -1470 6735 -1450 6755
rect -1430 6735 -1410 6755
rect -1390 6735 -1370 6755
rect -1350 6735 -1330 6755
rect -1310 6735 -1290 6755
rect -1270 6735 -1250 6755
rect -1230 6735 -1210 6755
rect -1190 6735 -1170 6755
rect -1150 6735 -1130 6755
rect -1110 6735 -1090 6755
rect -1070 6735 -1050 6755
rect -1030 6735 -1010 6755
rect -990 6735 -970 6755
rect -950 6735 -930 6755
rect -910 6735 -890 6755
rect -870 6735 -850 6755
rect -830 6735 -810 6755
rect -790 6735 -770 6755
rect -750 6735 -730 6755
rect -710 6735 -690 6755
rect -670 6735 -650 6755
rect -630 6735 -610 6755
rect -590 6735 -570 6755
rect -550 6735 -530 6755
rect -510 6735 -490 6755
rect -470 6735 -450 6755
rect -430 6735 -410 6755
rect -390 6735 -370 6755
rect -350 6735 -330 6755
rect -310 6735 -290 6755
rect -270 6735 -250 6755
rect -230 6735 -210 6755
rect -190 6735 -170 6755
rect -150 6735 -130 6755
rect -110 6735 -90 6755
rect -70 6735 -50 6755
rect -30 6735 -10 6755
rect 10 6735 30 6755
rect 50 6735 70 6755
rect 90 6735 110 6755
rect 130 6735 150 6755
rect 170 6735 190 6755
rect 210 6735 230 6755
rect 250 6735 270 6755
rect 290 6735 310 6755
rect 330 6735 350 6755
rect 370 6735 390 6755
rect 410 6735 430 6755
rect 450 6735 470 6755
rect 490 6735 510 6755
rect -1950 6653 -1930 6673
rect -1910 6653 -1890 6673
rect -1870 6653 -1850 6673
rect -1830 6653 -1810 6673
rect -1790 6653 -1770 6673
rect -1750 6653 -1730 6673
rect -1710 6653 -1690 6673
rect -1670 6653 -1650 6673
rect -1630 6653 -1610 6673
rect -1590 6653 -1570 6673
rect -1550 6653 -1530 6673
rect -1510 6653 -1490 6673
rect -1470 6653 -1450 6673
rect -1430 6653 -1410 6673
rect -1390 6653 -1370 6673
rect -1350 6653 -1330 6673
rect -1310 6653 -1290 6673
rect -1270 6653 -1250 6673
rect -1230 6653 -1210 6673
rect -1190 6653 -1170 6673
rect -1150 6653 -1130 6673
rect -1110 6653 -1090 6673
rect -1070 6653 -1050 6673
rect -1030 6653 -1010 6673
rect -990 6653 -970 6673
rect -950 6653 -930 6673
rect -910 6653 -890 6673
rect -870 6653 -850 6673
rect -830 6653 -810 6673
rect -790 6653 -770 6673
rect -750 6653 -730 6673
rect -710 6653 -690 6673
rect -670 6653 -650 6673
rect -630 6653 -610 6673
rect -590 6653 -570 6673
rect -550 6653 -530 6673
rect -510 6653 -490 6673
rect -470 6653 -450 6673
rect -430 6653 -410 6673
rect -390 6653 -370 6673
rect -350 6653 -330 6673
rect -310 6653 -290 6673
rect -270 6653 -250 6673
rect -230 6653 -210 6673
rect -190 6653 -170 6673
rect -150 6653 -130 6673
rect -110 6653 -90 6673
rect -70 6653 -50 6673
rect -30 6653 -10 6673
rect 10 6653 30 6673
rect 50 6653 70 6673
rect 90 6653 110 6673
rect 130 6653 150 6673
rect 170 6653 190 6673
rect 210 6653 230 6673
rect 250 6653 270 6673
rect 290 6653 310 6673
rect 330 6653 350 6673
rect 370 6653 390 6673
rect 410 6653 430 6673
rect 450 6653 470 6673
rect 490 6653 510 6673
rect -1950 6571 -1930 6591
rect -1910 6571 -1890 6591
rect -1870 6571 -1850 6591
rect -1830 6571 -1810 6591
rect -1790 6571 -1770 6591
rect -1750 6571 -1730 6591
rect -1710 6571 -1690 6591
rect -1670 6571 -1650 6591
rect -1630 6571 -1610 6591
rect -1590 6571 -1570 6591
rect -1550 6571 -1530 6591
rect -1510 6571 -1490 6591
rect -1470 6571 -1450 6591
rect -1430 6571 -1410 6591
rect -1390 6571 -1370 6591
rect -1350 6571 -1330 6591
rect -1310 6571 -1290 6591
rect -1270 6571 -1250 6591
rect -1230 6571 -1210 6591
rect -1190 6571 -1170 6591
rect -1150 6571 -1130 6591
rect -1110 6571 -1090 6591
rect -1070 6571 -1050 6591
rect -1030 6571 -1010 6591
rect -990 6571 -970 6591
rect -950 6571 -930 6591
rect -910 6571 -890 6591
rect -870 6571 -850 6591
rect -830 6571 -810 6591
rect -790 6571 -770 6591
rect -750 6571 -730 6591
rect -710 6571 -690 6591
rect -670 6571 -650 6591
rect -630 6571 -610 6591
rect -590 6571 -570 6591
rect -550 6571 -530 6591
rect -510 6571 -490 6591
rect -470 6571 -450 6591
rect -430 6571 -410 6591
rect -390 6571 -370 6591
rect -350 6571 -330 6591
rect -310 6571 -290 6591
rect -270 6571 -250 6591
rect -230 6571 -210 6591
rect -190 6571 -170 6591
rect -150 6571 -130 6591
rect -110 6571 -90 6591
rect -70 6571 -50 6591
rect -30 6571 -10 6591
rect 10 6571 30 6591
rect 50 6571 70 6591
rect 90 6571 110 6591
rect 130 6571 150 6591
rect 170 6571 190 6591
rect 210 6571 230 6591
rect 250 6571 270 6591
rect 290 6571 310 6591
rect 330 6571 350 6591
rect 370 6571 390 6591
rect 410 6571 430 6591
rect 450 6571 470 6591
rect 490 6571 510 6591
rect -1950 6489 -1930 6509
rect -1910 6489 -1890 6509
rect -1870 6489 -1850 6509
rect -1830 6489 -1810 6509
rect -1790 6489 -1770 6509
rect -1750 6489 -1730 6509
rect -1710 6489 -1690 6509
rect -1670 6489 -1650 6509
rect -1630 6489 -1610 6509
rect -1590 6489 -1570 6509
rect -1550 6489 -1530 6509
rect -1510 6489 -1490 6509
rect -1470 6489 -1450 6509
rect -1430 6489 -1410 6509
rect -1390 6489 -1370 6509
rect -1350 6489 -1330 6509
rect -1310 6489 -1290 6509
rect -1270 6489 -1250 6509
rect -1230 6489 -1210 6509
rect -1190 6489 -1170 6509
rect -1150 6489 -1130 6509
rect -1110 6489 -1090 6509
rect -1070 6489 -1050 6509
rect -1030 6489 -1010 6509
rect -990 6489 -970 6509
rect -950 6489 -930 6509
rect -910 6489 -890 6509
rect -870 6489 -850 6509
rect -830 6489 -810 6509
rect -790 6489 -770 6509
rect -750 6489 -730 6509
rect -710 6489 -690 6509
rect -670 6489 -650 6509
rect -630 6489 -610 6509
rect -590 6489 -570 6509
rect -550 6489 -530 6509
rect -510 6489 -490 6509
rect -470 6489 -450 6509
rect -430 6489 -410 6509
rect -390 6489 -370 6509
rect -350 6489 -330 6509
rect -310 6489 -290 6509
rect -270 6489 -250 6509
rect -230 6489 -210 6509
rect -190 6489 -170 6509
rect -150 6489 -130 6509
rect -110 6489 -90 6509
rect -70 6489 -50 6509
rect -30 6489 -10 6509
rect 10 6489 30 6509
rect 50 6489 70 6509
rect 90 6489 110 6509
rect 130 6489 150 6509
rect 170 6489 190 6509
rect 210 6489 230 6509
rect 250 6489 270 6509
rect 290 6489 310 6509
rect 330 6489 350 6509
rect 370 6489 390 6509
rect 410 6489 430 6509
rect 450 6489 470 6509
rect 490 6489 510 6509
rect -1950 6407 -1930 6427
rect -1910 6407 -1890 6427
rect -1870 6407 -1850 6427
rect -1830 6407 -1810 6427
rect -1790 6407 -1770 6427
rect -1750 6407 -1730 6427
rect -1710 6407 -1690 6427
rect -1670 6407 -1650 6427
rect -1630 6407 -1610 6427
rect -1590 6407 -1570 6427
rect -1550 6407 -1530 6427
rect -1510 6407 -1490 6427
rect -1470 6407 -1450 6427
rect -1430 6407 -1410 6427
rect -1390 6407 -1370 6427
rect -1350 6407 -1330 6427
rect -1310 6407 -1290 6427
rect -1270 6407 -1250 6427
rect -1230 6407 -1210 6427
rect -1190 6407 -1170 6427
rect -1150 6407 -1130 6427
rect -1110 6407 -1090 6427
rect -1070 6407 -1050 6427
rect -1030 6407 -1010 6427
rect -990 6407 -970 6427
rect -950 6407 -930 6427
rect -910 6407 -890 6427
rect -870 6407 -850 6427
rect -830 6407 -810 6427
rect -790 6407 -770 6427
rect -750 6407 -730 6427
rect -710 6407 -690 6427
rect -670 6407 -650 6427
rect -630 6407 -610 6427
rect -590 6407 -570 6427
rect -550 6407 -530 6427
rect -510 6407 -490 6427
rect -470 6407 -450 6427
rect -430 6407 -410 6427
rect -390 6407 -370 6427
rect -350 6407 -330 6427
rect -310 6407 -290 6427
rect -270 6407 -250 6427
rect -230 6407 -210 6427
rect -190 6407 -170 6427
rect -150 6407 -130 6427
rect -110 6407 -90 6427
rect -70 6407 -50 6427
rect -30 6407 -10 6427
rect 10 6407 30 6427
rect 50 6407 70 6427
rect 90 6407 110 6427
rect 130 6407 150 6427
rect 170 6407 190 6427
rect 210 6407 230 6427
rect 250 6407 270 6427
rect 290 6407 310 6427
rect 330 6407 350 6427
rect 370 6407 390 6427
rect 410 6407 430 6427
rect 450 6407 470 6427
rect 490 6407 510 6427
rect -1950 6325 -1930 6345
rect -1910 6325 -1890 6345
rect -1870 6325 -1850 6345
rect -1830 6325 -1810 6345
rect -1790 6325 -1770 6345
rect -1750 6325 -1730 6345
rect -1710 6325 -1690 6345
rect -1670 6325 -1650 6345
rect -1630 6325 -1610 6345
rect -1590 6325 -1570 6345
rect -1550 6325 -1530 6345
rect -1510 6325 -1490 6345
rect -1470 6325 -1450 6345
rect -1430 6325 -1410 6345
rect -1390 6325 -1370 6345
rect -1350 6325 -1330 6345
rect -1310 6325 -1290 6345
rect -1270 6325 -1250 6345
rect -1230 6325 -1210 6345
rect -1190 6325 -1170 6345
rect -1150 6325 -1130 6345
rect -1110 6325 -1090 6345
rect -1070 6325 -1050 6345
rect -1030 6325 -1010 6345
rect -990 6325 -970 6345
rect -950 6325 -930 6345
rect -910 6325 -890 6345
rect -870 6325 -850 6345
rect -830 6325 -810 6345
rect -790 6325 -770 6345
rect -750 6325 -730 6345
rect -710 6325 -690 6345
rect -670 6325 -650 6345
rect -630 6325 -610 6345
rect -590 6325 -570 6345
rect -550 6325 -530 6345
rect -510 6325 -490 6345
rect -470 6325 -450 6345
rect -430 6325 -410 6345
rect -390 6325 -370 6345
rect -350 6325 -330 6345
rect -310 6325 -290 6345
rect -270 6325 -250 6345
rect -230 6325 -210 6345
rect -190 6325 -170 6345
rect -150 6325 -130 6345
rect -110 6325 -90 6345
rect -70 6325 -50 6345
rect -30 6325 -10 6345
rect 10 6325 30 6345
rect 50 6325 70 6345
rect 90 6325 110 6345
rect 130 6325 150 6345
rect 170 6325 190 6345
rect 210 6325 230 6345
rect 250 6325 270 6345
rect 290 6325 310 6345
rect 330 6325 350 6345
rect 370 6325 390 6345
rect 410 6325 430 6345
rect 450 6325 470 6345
rect 490 6325 510 6345
rect -5580 6025 -5550 6045
rect -5530 6025 -5510 6045
rect -5490 6025 -5470 6045
rect -5450 6025 -5430 6045
rect -5410 6025 -5390 6045
rect -5370 6025 -5350 6045
rect -5330 6025 -5310 6045
rect -5290 6025 -5270 6045
rect -5250 6025 -5230 6045
rect -5210 6025 -5190 6045
rect -5170 6025 -5150 6045
rect -5130 6025 -5110 6045
rect -5090 6025 -5070 6045
rect -5050 6025 -5030 6045
rect -5010 6025 -4990 6045
rect -4970 6025 -4950 6045
rect -4930 6025 -4910 6045
rect -4890 6025 -4870 6045
rect -4850 6025 -4830 6045
rect -4810 6025 -4790 6045
rect -4770 6025 -4750 6045
rect -4730 6025 -4710 6045
rect -4690 6025 -4670 6045
rect -4650 6025 -4630 6045
rect -4610 6025 -4590 6045
rect -4570 6025 -4550 6045
rect -4530 6025 -4510 6045
rect -4490 6025 -4470 6045
rect -4450 6025 -4430 6045
rect -4410 6025 -4390 6045
rect -4370 6025 -4350 6045
rect -4330 6025 -4310 6045
rect -4290 6025 -4270 6045
rect -4250 6025 -4230 6045
rect -4210 6025 -4190 6045
rect -4170 6025 -4150 6045
rect -4130 6025 -4110 6045
rect -4090 6025 -4070 6045
rect -4050 6025 -4030 6045
rect -4010 6025 -3990 6045
rect -3970 6025 -3950 6045
rect -3930 6025 -3910 6045
rect -3890 6025 -3870 6045
rect -3850 6025 -3830 6045
rect -3810 6025 -3790 6045
rect -3770 6025 -3750 6045
rect -3730 6025 -3710 6045
rect -3690 6025 -3670 6045
rect -3650 6025 -3630 6045
rect -3610 6025 -3590 6045
rect -3570 6025 -3550 6045
rect -3530 6025 -3510 6045
rect -3490 6025 -3470 6045
rect -3450 6025 -3430 6045
rect -3410 6025 -3390 6045
rect -3370 6025 -3350 6045
rect -3330 6025 -3310 6045
rect -3290 6025 -3270 6045
rect -3250 6025 -3230 6045
rect -3210 6025 -3190 6045
rect -3170 6025 -3150 6045
rect -3130 6025 -3110 6045
rect -2030 6025 -2010 6045
rect -1990 6025 -1970 6045
rect -1950 6025 -1930 6045
rect -1910 6025 -1890 6045
rect -1870 6025 -1850 6045
rect -1830 6025 -1810 6045
rect -1790 6025 -1770 6045
rect -1750 6025 -1730 6045
rect -1710 6025 -1690 6045
rect -1670 6025 -1650 6045
rect -1630 6025 -1610 6045
rect -1590 6025 -1570 6045
rect -1550 6025 -1530 6045
rect -1510 6025 -1490 6045
rect -1470 6025 -1450 6045
rect -1430 6025 -1410 6045
rect -1390 6025 -1370 6045
rect -1350 6025 -1330 6045
rect -1310 6025 -1290 6045
rect -1270 6025 -1250 6045
rect -1230 6025 -1210 6045
rect -1190 6025 -1170 6045
rect -1150 6025 -1130 6045
rect -1110 6025 -1090 6045
rect -1070 6025 -1050 6045
rect -1030 6025 -1010 6045
rect -990 6025 -970 6045
rect -950 6025 -930 6045
rect -910 6025 -890 6045
rect -870 6025 -850 6045
rect -830 6025 -810 6045
rect -790 6025 -770 6045
rect -750 6025 -730 6045
rect -710 6025 -690 6045
rect -670 6025 -650 6045
rect -630 6025 -610 6045
rect -590 6025 -570 6045
rect -550 6025 -530 6045
rect -510 6025 -490 6045
rect -470 6025 -450 6045
rect -430 6025 -410 6045
rect -390 6025 -370 6045
rect -350 6025 -330 6045
rect -310 6025 -290 6045
rect -270 6025 -250 6045
rect -230 6025 -210 6045
rect -190 6025 -170 6045
rect -150 6025 -130 6045
rect -110 6025 -90 6045
rect -70 6025 -50 6045
rect -30 6025 -10 6045
rect 10 6025 30 6045
rect 50 6025 70 6045
rect 90 6025 110 6045
rect 130 6025 150 6045
rect 170 6025 190 6045
rect 210 6025 230 6045
rect 250 6025 270 6045
rect 290 6025 310 6045
rect 330 6025 350 6045
rect 370 6025 390 6045
rect 410 6025 440 6045
rect -5580 5930 -5550 5950
rect -5530 5930 -5510 5950
rect -5490 5930 -5470 5950
rect -5450 5930 -5430 5950
rect -5410 5930 -5390 5950
rect -5370 5930 -5350 5950
rect -5330 5930 -5310 5950
rect -5290 5930 -5270 5950
rect -5250 5930 -5230 5950
rect -5210 5930 -5190 5950
rect -5170 5930 -5150 5950
rect -5130 5930 -5110 5950
rect -5090 5930 -5070 5950
rect -5050 5930 -5030 5950
rect -5010 5930 -4990 5950
rect -4970 5930 -4950 5950
rect -4930 5930 -4910 5950
rect -4890 5930 -4870 5950
rect -4850 5930 -4830 5950
rect -4810 5930 -4790 5950
rect -4770 5930 -4750 5950
rect -4730 5930 -4710 5950
rect -4690 5930 -4670 5950
rect -4650 5930 -4630 5950
rect -4610 5930 -4590 5950
rect -4570 5930 -4550 5950
rect -4530 5930 -4510 5950
rect -4490 5930 -4470 5950
rect -4450 5930 -4430 5950
rect -4410 5930 -4390 5950
rect -4370 5930 -4350 5950
rect -4330 5930 -4310 5950
rect -4290 5930 -4270 5950
rect -4250 5930 -4230 5950
rect -4210 5930 -4190 5950
rect -4170 5930 -4150 5950
rect -4130 5930 -4110 5950
rect -4090 5930 -4070 5950
rect -4050 5930 -4030 5950
rect -4010 5930 -3990 5950
rect -3970 5930 -3950 5950
rect -3930 5930 -3910 5950
rect -3890 5930 -3870 5950
rect -3850 5930 -3830 5950
rect -3810 5930 -3790 5950
rect -3770 5930 -3750 5950
rect -3730 5930 -3710 5950
rect -3690 5930 -3670 5950
rect -3650 5930 -3630 5950
rect -3610 5930 -3590 5950
rect -3570 5930 -3550 5950
rect -3530 5930 -3510 5950
rect -3490 5930 -3470 5950
rect -3450 5930 -3430 5950
rect -3410 5930 -3390 5950
rect -3370 5930 -3350 5950
rect -3330 5930 -3310 5950
rect -3290 5930 -3270 5950
rect -3250 5930 -3230 5950
rect -3210 5930 -3190 5950
rect -3170 5930 -3150 5950
rect -3130 5930 -3110 5950
rect -2030 5930 -2010 5950
rect -1990 5930 -1970 5950
rect -1950 5930 -1930 5950
rect -1910 5930 -1890 5950
rect -1870 5930 -1850 5950
rect -1830 5930 -1810 5950
rect -1790 5930 -1770 5950
rect -1750 5930 -1730 5950
rect -1710 5930 -1690 5950
rect -1670 5930 -1650 5950
rect -1630 5930 -1610 5950
rect -1590 5930 -1570 5950
rect -1550 5930 -1530 5950
rect -1510 5930 -1490 5950
rect -1470 5930 -1450 5950
rect -1430 5930 -1410 5950
rect -1390 5930 -1370 5950
rect -1350 5930 -1330 5950
rect -1310 5930 -1290 5950
rect -1270 5930 -1250 5950
rect -1230 5930 -1210 5950
rect -1190 5930 -1170 5950
rect -1150 5930 -1130 5950
rect -1110 5930 -1090 5950
rect -1070 5930 -1050 5950
rect -1030 5930 -1010 5950
rect -990 5930 -970 5950
rect -950 5930 -930 5950
rect -910 5930 -890 5950
rect -870 5930 -850 5950
rect -830 5930 -810 5950
rect -790 5930 -770 5950
rect -750 5930 -730 5950
rect -710 5930 -690 5950
rect -670 5930 -650 5950
rect -630 5930 -610 5950
rect -590 5930 -570 5950
rect -550 5930 -530 5950
rect -510 5930 -490 5950
rect -470 5930 -450 5950
rect -430 5930 -410 5950
rect -390 5930 -370 5950
rect -350 5930 -330 5950
rect -310 5930 -290 5950
rect -270 5930 -250 5950
rect -230 5930 -210 5950
rect -190 5930 -170 5950
rect -150 5930 -130 5950
rect -110 5930 -90 5950
rect -70 5930 -50 5950
rect -30 5930 -10 5950
rect 10 5930 30 5950
rect 50 5930 70 5950
rect 90 5930 110 5950
rect 130 5930 150 5950
rect 170 5930 190 5950
rect 210 5930 230 5950
rect 250 5930 270 5950
rect 290 5930 310 5950
rect 330 5930 350 5950
rect 370 5930 390 5950
rect 410 5930 440 5950
rect -5580 5835 -5550 5855
rect -5530 5835 -5510 5855
rect -5490 5835 -5470 5855
rect -5450 5835 -5430 5855
rect -5410 5835 -5390 5855
rect -5370 5835 -5350 5855
rect -5330 5835 -5310 5855
rect -5290 5835 -5270 5855
rect -5250 5835 -5230 5855
rect -5210 5835 -5190 5855
rect -5170 5835 -5150 5855
rect -5130 5835 -5110 5855
rect -5090 5835 -5070 5855
rect -5050 5835 -5030 5855
rect -5010 5835 -4990 5855
rect -4970 5835 -4950 5855
rect -4930 5835 -4910 5855
rect -4890 5835 -4870 5855
rect -4850 5835 -4830 5855
rect -4810 5835 -4790 5855
rect -4770 5835 -4750 5855
rect -4730 5835 -4710 5855
rect -4690 5835 -4670 5855
rect -4650 5835 -4630 5855
rect -4610 5835 -4590 5855
rect -4570 5835 -4550 5855
rect -4530 5835 -4510 5855
rect -4490 5835 -4470 5855
rect -4450 5835 -4430 5855
rect -4410 5835 -4390 5855
rect -4370 5835 -4350 5855
rect -4330 5835 -4310 5855
rect -4290 5835 -4270 5855
rect -4250 5835 -4230 5855
rect -4210 5835 -4190 5855
rect -4170 5835 -4150 5855
rect -4130 5835 -4110 5855
rect -4090 5835 -4070 5855
rect -4050 5835 -4030 5855
rect -4010 5835 -3990 5855
rect -3970 5835 -3950 5855
rect -3930 5835 -3910 5855
rect -3890 5835 -3870 5855
rect -3850 5835 -3830 5855
rect -3810 5835 -3790 5855
rect -3770 5835 -3750 5855
rect -3730 5835 -3710 5855
rect -3690 5835 -3670 5855
rect -3650 5835 -3630 5855
rect -3610 5835 -3590 5855
rect -3570 5835 -3550 5855
rect -3530 5835 -3510 5855
rect -3490 5835 -3470 5855
rect -3450 5835 -3430 5855
rect -3410 5835 -3390 5855
rect -3370 5835 -3350 5855
rect -3330 5835 -3310 5855
rect -3290 5835 -3270 5855
rect -3250 5835 -3230 5855
rect -3210 5835 -3190 5855
rect -3170 5835 -3150 5855
rect -3130 5835 -3110 5855
rect -2030 5835 -2010 5855
rect -1990 5835 -1970 5855
rect -1950 5835 -1930 5855
rect -1910 5835 -1890 5855
rect -1870 5835 -1850 5855
rect -1830 5835 -1810 5855
rect -1790 5835 -1770 5855
rect -1750 5835 -1730 5855
rect -1710 5835 -1690 5855
rect -1670 5835 -1650 5855
rect -1630 5835 -1610 5855
rect -1590 5835 -1570 5855
rect -1550 5835 -1530 5855
rect -1510 5835 -1490 5855
rect -1470 5835 -1450 5855
rect -1430 5835 -1410 5855
rect -1390 5835 -1370 5855
rect -1350 5835 -1330 5855
rect -1310 5835 -1290 5855
rect -1270 5835 -1250 5855
rect -1230 5835 -1210 5855
rect -1190 5835 -1170 5855
rect -1150 5835 -1130 5855
rect -1110 5835 -1090 5855
rect -1070 5835 -1050 5855
rect -1030 5835 -1010 5855
rect -990 5835 -970 5855
rect -950 5835 -930 5855
rect -910 5835 -890 5855
rect -870 5835 -850 5855
rect -830 5835 -810 5855
rect -790 5835 -770 5855
rect -750 5835 -730 5855
rect -710 5835 -690 5855
rect -670 5835 -650 5855
rect -630 5835 -610 5855
rect -590 5835 -570 5855
rect -550 5835 -530 5855
rect -510 5835 -490 5855
rect -470 5835 -450 5855
rect -430 5835 -410 5855
rect -390 5835 -370 5855
rect -350 5835 -330 5855
rect -310 5835 -290 5855
rect -270 5835 -250 5855
rect -230 5835 -210 5855
rect -190 5835 -170 5855
rect -150 5835 -130 5855
rect -110 5835 -90 5855
rect -70 5835 -50 5855
rect -30 5835 -10 5855
rect 10 5835 30 5855
rect 50 5835 70 5855
rect 90 5835 110 5855
rect 130 5835 150 5855
rect 170 5835 190 5855
rect 210 5835 230 5855
rect 250 5835 270 5855
rect 290 5835 310 5855
rect 330 5835 350 5855
rect 370 5835 390 5855
rect 410 5835 440 5855
rect -5580 5740 -5550 5760
rect -5530 5740 -5510 5760
rect -5490 5740 -5470 5760
rect -5450 5740 -5430 5760
rect -5410 5740 -5390 5760
rect -5370 5740 -5350 5760
rect -5330 5740 -5310 5760
rect -5290 5740 -5270 5760
rect -5250 5740 -5230 5760
rect -5210 5740 -5190 5760
rect -5170 5740 -5150 5760
rect -5130 5740 -5110 5760
rect -5090 5740 -5070 5760
rect -5050 5740 -5030 5760
rect -5010 5740 -4990 5760
rect -4970 5740 -4950 5760
rect -4930 5740 -4910 5760
rect -4890 5740 -4870 5760
rect -4850 5740 -4830 5760
rect -4810 5740 -4790 5760
rect -4770 5740 -4750 5760
rect -4730 5740 -4710 5760
rect -4690 5740 -4670 5760
rect -4650 5740 -4630 5760
rect -4610 5740 -4590 5760
rect -4570 5740 -4550 5760
rect -4530 5740 -4510 5760
rect -4490 5740 -4470 5760
rect -4450 5740 -4430 5760
rect -4410 5740 -4390 5760
rect -4370 5740 -4350 5760
rect -4330 5740 -4310 5760
rect -4290 5740 -4270 5760
rect -4250 5740 -4230 5760
rect -4210 5740 -4190 5760
rect -4170 5740 -4150 5760
rect -4130 5740 -4110 5760
rect -4090 5740 -4070 5760
rect -4050 5740 -4030 5760
rect -4010 5740 -3990 5760
rect -3970 5740 -3950 5760
rect -3930 5740 -3910 5760
rect -3890 5740 -3870 5760
rect -3850 5740 -3830 5760
rect -3810 5740 -3790 5760
rect -3770 5740 -3750 5760
rect -3730 5740 -3710 5760
rect -3690 5740 -3670 5760
rect -3650 5740 -3630 5760
rect -3610 5740 -3590 5760
rect -3570 5740 -3550 5760
rect -3530 5740 -3510 5760
rect -3490 5740 -3470 5760
rect -3450 5740 -3430 5760
rect -3410 5740 -3390 5760
rect -3370 5740 -3350 5760
rect -3330 5740 -3310 5760
rect -3290 5740 -3270 5760
rect -3250 5740 -3230 5760
rect -3210 5740 -3190 5760
rect -3170 5740 -3150 5760
rect -3130 5740 -3110 5760
rect -2030 5740 -2010 5760
rect -1990 5740 -1970 5760
rect -1950 5740 -1930 5760
rect -1910 5740 -1890 5760
rect -1870 5740 -1850 5760
rect -1830 5740 -1810 5760
rect -1790 5740 -1770 5760
rect -1750 5740 -1730 5760
rect -1710 5740 -1690 5760
rect -1670 5740 -1650 5760
rect -1630 5740 -1610 5760
rect -1590 5740 -1570 5760
rect -1550 5740 -1530 5760
rect -1510 5740 -1490 5760
rect -1470 5740 -1450 5760
rect -1430 5740 -1410 5760
rect -1390 5740 -1370 5760
rect -1350 5740 -1330 5760
rect -1310 5740 -1290 5760
rect -1270 5740 -1250 5760
rect -1230 5740 -1210 5760
rect -1190 5740 -1170 5760
rect -1150 5740 -1130 5760
rect -1110 5740 -1090 5760
rect -1070 5740 -1050 5760
rect -1030 5740 -1010 5760
rect -990 5740 -970 5760
rect -950 5740 -930 5760
rect -910 5740 -890 5760
rect -870 5740 -850 5760
rect -830 5740 -810 5760
rect -790 5740 -770 5760
rect -750 5740 -730 5760
rect -710 5740 -690 5760
rect -670 5740 -650 5760
rect -630 5740 -610 5760
rect -590 5740 -570 5760
rect -550 5740 -530 5760
rect -510 5740 -490 5760
rect -470 5740 -450 5760
rect -430 5740 -410 5760
rect -390 5740 -370 5760
rect -350 5740 -330 5760
rect -310 5740 -290 5760
rect -270 5740 -250 5760
rect -230 5740 -210 5760
rect -190 5740 -170 5760
rect -150 5740 -130 5760
rect -110 5740 -90 5760
rect -70 5740 -50 5760
rect -30 5740 -10 5760
rect 10 5740 30 5760
rect 50 5740 70 5760
rect 90 5740 110 5760
rect 130 5740 150 5760
rect 170 5740 190 5760
rect 210 5740 230 5760
rect 250 5740 270 5760
rect 290 5740 310 5760
rect 330 5740 350 5760
rect 370 5740 390 5760
rect 410 5740 440 5760
rect -5580 5645 -5550 5665
rect -5530 5645 -5510 5665
rect -5490 5645 -5470 5665
rect -5450 5645 -5430 5665
rect -5410 5645 -5390 5665
rect -5370 5645 -5350 5665
rect -5330 5645 -5310 5665
rect -5290 5645 -5270 5665
rect -5250 5645 -5230 5665
rect -5210 5645 -5190 5665
rect -5170 5645 -5150 5665
rect -5130 5645 -5110 5665
rect -5090 5645 -5070 5665
rect -5050 5645 -5030 5665
rect -5010 5645 -4990 5665
rect -4970 5645 -4950 5665
rect -4930 5645 -4910 5665
rect -4890 5645 -4870 5665
rect -4850 5645 -4830 5665
rect -4810 5645 -4790 5665
rect -4770 5645 -4750 5665
rect -4730 5645 -4710 5665
rect -4690 5645 -4670 5665
rect -4650 5645 -4630 5665
rect -4610 5645 -4590 5665
rect -4570 5645 -4550 5665
rect -4530 5645 -4510 5665
rect -4490 5645 -4470 5665
rect -4450 5645 -4430 5665
rect -4410 5645 -4390 5665
rect -4370 5645 -4350 5665
rect -4330 5645 -4310 5665
rect -4290 5645 -4270 5665
rect -4250 5645 -4230 5665
rect -4210 5645 -4190 5665
rect -4170 5645 -4150 5665
rect -4130 5645 -4110 5665
rect -4090 5645 -4070 5665
rect -4050 5645 -4030 5665
rect -4010 5645 -3990 5665
rect -3970 5645 -3950 5665
rect -3930 5645 -3910 5665
rect -3890 5645 -3870 5665
rect -3850 5645 -3830 5665
rect -3810 5645 -3790 5665
rect -3770 5645 -3750 5665
rect -3730 5645 -3710 5665
rect -3690 5645 -3670 5665
rect -3650 5645 -3630 5665
rect -3610 5645 -3590 5665
rect -3570 5645 -3550 5665
rect -3530 5645 -3510 5665
rect -3490 5645 -3470 5665
rect -3450 5645 -3430 5665
rect -3410 5645 -3390 5665
rect -3370 5645 -3350 5665
rect -3330 5645 -3310 5665
rect -3290 5645 -3270 5665
rect -3250 5645 -3230 5665
rect -3210 5645 -3190 5665
rect -3170 5645 -3150 5665
rect -3130 5645 -3110 5665
rect -2030 5645 -2010 5665
rect -1990 5645 -1970 5665
rect -1950 5645 -1930 5665
rect -1910 5645 -1890 5665
rect -1870 5645 -1850 5665
rect -1830 5645 -1810 5665
rect -1790 5645 -1770 5665
rect -1750 5645 -1730 5665
rect -1710 5645 -1690 5665
rect -1670 5645 -1650 5665
rect -1630 5645 -1610 5665
rect -1590 5645 -1570 5665
rect -1550 5645 -1530 5665
rect -1510 5645 -1490 5665
rect -1470 5645 -1450 5665
rect -1430 5645 -1410 5665
rect -1390 5645 -1370 5665
rect -1350 5645 -1330 5665
rect -1310 5645 -1290 5665
rect -1270 5645 -1250 5665
rect -1230 5645 -1210 5665
rect -1190 5645 -1170 5665
rect -1150 5645 -1130 5665
rect -1110 5645 -1090 5665
rect -1070 5645 -1050 5665
rect -1030 5645 -1010 5665
rect -990 5645 -970 5665
rect -950 5645 -930 5665
rect -910 5645 -890 5665
rect -870 5645 -850 5665
rect -830 5645 -810 5665
rect -790 5645 -770 5665
rect -750 5645 -730 5665
rect -710 5645 -690 5665
rect -670 5645 -650 5665
rect -630 5645 -610 5665
rect -590 5645 -570 5665
rect -550 5645 -530 5665
rect -510 5645 -490 5665
rect -470 5645 -450 5665
rect -430 5645 -410 5665
rect -390 5645 -370 5665
rect -350 5645 -330 5665
rect -310 5645 -290 5665
rect -270 5645 -250 5665
rect -230 5645 -210 5665
rect -190 5645 -170 5665
rect -150 5645 -130 5665
rect -110 5645 -90 5665
rect -70 5645 -50 5665
rect -30 5645 -10 5665
rect 10 5645 30 5665
rect 50 5645 70 5665
rect 90 5645 110 5665
rect 130 5645 150 5665
rect 170 5645 190 5665
rect 210 5645 230 5665
rect 250 5645 270 5665
rect 290 5645 310 5665
rect 330 5645 350 5665
rect 370 5645 390 5665
rect 410 5645 440 5665
rect -5580 5550 -5550 5570
rect -5530 5550 -5510 5570
rect -5490 5550 -5470 5570
rect -5450 5550 -5430 5570
rect -5410 5550 -5390 5570
rect -5370 5550 -5350 5570
rect -5330 5550 -5310 5570
rect -5290 5550 -5270 5570
rect -5250 5550 -5230 5570
rect -5210 5550 -5190 5570
rect -5170 5550 -5150 5570
rect -5130 5550 -5110 5570
rect -5090 5550 -5070 5570
rect -5050 5550 -5030 5570
rect -5010 5550 -4990 5570
rect -4970 5550 -4950 5570
rect -4930 5550 -4910 5570
rect -4890 5550 -4870 5570
rect -4850 5550 -4830 5570
rect -4810 5550 -4790 5570
rect -4770 5550 -4750 5570
rect -4730 5550 -4710 5570
rect -4690 5550 -4670 5570
rect -4650 5550 -4630 5570
rect -4610 5550 -4590 5570
rect -4570 5550 -4550 5570
rect -4530 5550 -4510 5570
rect -4490 5550 -4470 5570
rect -4450 5550 -4430 5570
rect -4410 5550 -4390 5570
rect -4370 5550 -4350 5570
rect -4330 5550 -4310 5570
rect -4290 5550 -4270 5570
rect -4250 5550 -4230 5570
rect -4210 5550 -4190 5570
rect -4170 5550 -4150 5570
rect -4130 5550 -4110 5570
rect -4090 5550 -4070 5570
rect -4050 5550 -4030 5570
rect -4010 5550 -3990 5570
rect -3970 5550 -3950 5570
rect -3930 5550 -3910 5570
rect -3890 5550 -3870 5570
rect -3850 5550 -3830 5570
rect -3810 5550 -3790 5570
rect -3770 5550 -3750 5570
rect -3730 5550 -3710 5570
rect -3690 5550 -3670 5570
rect -3650 5550 -3630 5570
rect -3610 5550 -3590 5570
rect -3570 5550 -3550 5570
rect -3530 5550 -3510 5570
rect -3490 5550 -3470 5570
rect -3450 5550 -3430 5570
rect -3410 5550 -3390 5570
rect -3370 5550 -3350 5570
rect -3330 5550 -3310 5570
rect -3290 5550 -3270 5570
rect -3250 5550 -3230 5570
rect -3210 5550 -3190 5570
rect -3170 5550 -3150 5570
rect -3130 5550 -3110 5570
rect -2030 5550 -2010 5570
rect -1990 5550 -1970 5570
rect -1950 5550 -1930 5570
rect -1910 5550 -1890 5570
rect -1870 5550 -1850 5570
rect -1830 5550 -1810 5570
rect -1790 5550 -1770 5570
rect -1750 5550 -1730 5570
rect -1710 5550 -1690 5570
rect -1670 5550 -1650 5570
rect -1630 5550 -1610 5570
rect -1590 5550 -1570 5570
rect -1550 5550 -1530 5570
rect -1510 5550 -1490 5570
rect -1470 5550 -1450 5570
rect -1430 5550 -1410 5570
rect -1390 5550 -1370 5570
rect -1350 5550 -1330 5570
rect -1310 5550 -1290 5570
rect -1270 5550 -1250 5570
rect -1230 5550 -1210 5570
rect -1190 5550 -1170 5570
rect -1150 5550 -1130 5570
rect -1110 5550 -1090 5570
rect -1070 5550 -1050 5570
rect -1030 5550 -1010 5570
rect -990 5550 -970 5570
rect -950 5550 -930 5570
rect -910 5550 -890 5570
rect -870 5550 -850 5570
rect -830 5550 -810 5570
rect -790 5550 -770 5570
rect -750 5550 -730 5570
rect -710 5550 -690 5570
rect -670 5550 -650 5570
rect -630 5550 -610 5570
rect -590 5550 -570 5570
rect -550 5550 -530 5570
rect -510 5550 -490 5570
rect -470 5550 -450 5570
rect -430 5550 -410 5570
rect -390 5550 -370 5570
rect -350 5550 -330 5570
rect -310 5550 -290 5570
rect -270 5550 -250 5570
rect -230 5550 -210 5570
rect -190 5550 -170 5570
rect -150 5550 -130 5570
rect -110 5550 -90 5570
rect -70 5550 -50 5570
rect -30 5550 -10 5570
rect 10 5550 30 5570
rect 50 5550 70 5570
rect 90 5550 110 5570
rect 130 5550 150 5570
rect 170 5550 190 5570
rect 210 5550 230 5570
rect 250 5550 270 5570
rect 290 5550 310 5570
rect 330 5550 350 5570
rect 370 5550 390 5570
rect 410 5550 440 5570
rect -5580 5455 -5550 5475
rect -5530 5455 -5510 5475
rect -5490 5455 -5470 5475
rect -5450 5455 -5430 5475
rect -5410 5455 -5390 5475
rect -5370 5455 -5350 5475
rect -5330 5455 -5310 5475
rect -5290 5455 -5270 5475
rect -5250 5455 -5230 5475
rect -5210 5455 -5190 5475
rect -5170 5455 -5150 5475
rect -5130 5455 -5110 5475
rect -5090 5455 -5070 5475
rect -5050 5455 -5030 5475
rect -5010 5455 -4990 5475
rect -4970 5455 -4950 5475
rect -4930 5455 -4910 5475
rect -4890 5455 -4870 5475
rect -4850 5455 -4830 5475
rect -4810 5455 -4790 5475
rect -4770 5455 -4750 5475
rect -4730 5455 -4710 5475
rect -4690 5455 -4670 5475
rect -4650 5455 -4630 5475
rect -4610 5455 -4590 5475
rect -4570 5455 -4550 5475
rect -4530 5455 -4510 5475
rect -4490 5455 -4470 5475
rect -4450 5455 -4430 5475
rect -4410 5455 -4390 5475
rect -4370 5455 -4350 5475
rect -4330 5455 -4310 5475
rect -4290 5455 -4270 5475
rect -4250 5455 -4230 5475
rect -4210 5455 -4190 5475
rect -4170 5455 -4150 5475
rect -4130 5455 -4110 5475
rect -4090 5455 -4070 5475
rect -4050 5455 -4030 5475
rect -4010 5455 -3990 5475
rect -3970 5455 -3950 5475
rect -3930 5455 -3910 5475
rect -3890 5455 -3870 5475
rect -3850 5455 -3830 5475
rect -3810 5455 -3790 5475
rect -3770 5455 -3750 5475
rect -3730 5455 -3710 5475
rect -3690 5455 -3670 5475
rect -3650 5455 -3630 5475
rect -3610 5455 -3590 5475
rect -3570 5455 -3550 5475
rect -3530 5455 -3510 5475
rect -3490 5455 -3470 5475
rect -3450 5455 -3430 5475
rect -3410 5455 -3390 5475
rect -3370 5455 -3350 5475
rect -3330 5455 -3310 5475
rect -3290 5455 -3270 5475
rect -3250 5455 -3230 5475
rect -3210 5455 -3190 5475
rect -3170 5455 -3150 5475
rect -3130 5455 -3110 5475
rect -2030 5455 -2010 5475
rect -1990 5455 -1970 5475
rect -1950 5455 -1930 5475
rect -1910 5455 -1890 5475
rect -1870 5455 -1850 5475
rect -1830 5455 -1810 5475
rect -1790 5455 -1770 5475
rect -1750 5455 -1730 5475
rect -1710 5455 -1690 5475
rect -1670 5455 -1650 5475
rect -1630 5455 -1610 5475
rect -1590 5455 -1570 5475
rect -1550 5455 -1530 5475
rect -1510 5455 -1490 5475
rect -1470 5455 -1450 5475
rect -1430 5455 -1410 5475
rect -1390 5455 -1370 5475
rect -1350 5455 -1330 5475
rect -1310 5455 -1290 5475
rect -1270 5455 -1250 5475
rect -1230 5455 -1210 5475
rect -1190 5455 -1170 5475
rect -1150 5455 -1130 5475
rect -1110 5455 -1090 5475
rect -1070 5455 -1050 5475
rect -1030 5455 -1010 5475
rect -990 5455 -970 5475
rect -950 5455 -930 5475
rect -910 5455 -890 5475
rect -870 5455 -850 5475
rect -830 5455 -810 5475
rect -790 5455 -770 5475
rect -750 5455 -730 5475
rect -710 5455 -690 5475
rect -670 5455 -650 5475
rect -630 5455 -610 5475
rect -590 5455 -570 5475
rect -550 5455 -530 5475
rect -510 5455 -490 5475
rect -470 5455 -450 5475
rect -430 5455 -410 5475
rect -390 5455 -370 5475
rect -350 5455 -330 5475
rect -310 5455 -290 5475
rect -270 5455 -250 5475
rect -230 5455 -210 5475
rect -190 5455 -170 5475
rect -150 5455 -130 5475
rect -110 5455 -90 5475
rect -70 5455 -50 5475
rect -30 5455 -10 5475
rect 10 5455 30 5475
rect 50 5455 70 5475
rect 90 5455 110 5475
rect 130 5455 150 5475
rect 170 5455 190 5475
rect 210 5455 230 5475
rect 250 5455 270 5475
rect 290 5455 310 5475
rect 330 5455 350 5475
rect 370 5455 390 5475
rect 410 5455 440 5475
rect -5580 5360 -5550 5380
rect -5530 5360 -5510 5380
rect -5490 5360 -5470 5380
rect -5450 5360 -5430 5380
rect -5410 5360 -5390 5380
rect -5370 5360 -5350 5380
rect -5330 5360 -5310 5380
rect -5290 5360 -5270 5380
rect -5250 5360 -5230 5380
rect -5210 5360 -5190 5380
rect -5170 5360 -5150 5380
rect -5130 5360 -5110 5380
rect -5090 5360 -5070 5380
rect -5050 5360 -5030 5380
rect -5010 5360 -4990 5380
rect -4970 5360 -4950 5380
rect -4930 5360 -4910 5380
rect -4890 5360 -4870 5380
rect -4850 5360 -4830 5380
rect -4810 5360 -4790 5380
rect -4770 5360 -4750 5380
rect -4730 5360 -4710 5380
rect -4690 5360 -4670 5380
rect -4650 5360 -4630 5380
rect -4610 5360 -4590 5380
rect -4570 5360 -4550 5380
rect -4530 5360 -4510 5380
rect -4490 5360 -4470 5380
rect -4450 5360 -4430 5380
rect -4410 5360 -4390 5380
rect -4370 5360 -4350 5380
rect -4330 5360 -4310 5380
rect -4290 5360 -4270 5380
rect -4250 5360 -4230 5380
rect -4210 5360 -4190 5380
rect -4170 5360 -4150 5380
rect -4130 5360 -4110 5380
rect -4090 5360 -4070 5380
rect -4050 5360 -4030 5380
rect -4010 5360 -3990 5380
rect -3970 5360 -3950 5380
rect -3930 5360 -3910 5380
rect -3890 5360 -3870 5380
rect -3850 5360 -3830 5380
rect -3810 5360 -3790 5380
rect -3770 5360 -3750 5380
rect -3730 5360 -3710 5380
rect -3690 5360 -3670 5380
rect -3650 5360 -3630 5380
rect -3610 5360 -3590 5380
rect -3570 5360 -3550 5380
rect -3530 5360 -3510 5380
rect -3490 5360 -3470 5380
rect -3450 5360 -3430 5380
rect -3410 5360 -3390 5380
rect -3370 5360 -3350 5380
rect -3330 5360 -3310 5380
rect -3290 5360 -3270 5380
rect -3250 5360 -3230 5380
rect -3210 5360 -3190 5380
rect -3170 5360 -3150 5380
rect -3130 5360 -3110 5380
rect -2030 5360 -2010 5380
rect -1990 5360 -1970 5380
rect -1950 5360 -1930 5380
rect -1910 5360 -1890 5380
rect -1870 5360 -1850 5380
rect -1830 5360 -1810 5380
rect -1790 5360 -1770 5380
rect -1750 5360 -1730 5380
rect -1710 5360 -1690 5380
rect -1670 5360 -1650 5380
rect -1630 5360 -1610 5380
rect -1590 5360 -1570 5380
rect -1550 5360 -1530 5380
rect -1510 5360 -1490 5380
rect -1470 5360 -1450 5380
rect -1430 5360 -1410 5380
rect -1390 5360 -1370 5380
rect -1350 5360 -1330 5380
rect -1310 5360 -1290 5380
rect -1270 5360 -1250 5380
rect -1230 5360 -1210 5380
rect -1190 5360 -1170 5380
rect -1150 5360 -1130 5380
rect -1110 5360 -1090 5380
rect -1070 5360 -1050 5380
rect -1030 5360 -1010 5380
rect -990 5360 -970 5380
rect -950 5360 -930 5380
rect -910 5360 -890 5380
rect -870 5360 -850 5380
rect -830 5360 -810 5380
rect -790 5360 -770 5380
rect -750 5360 -730 5380
rect -710 5360 -690 5380
rect -670 5360 -650 5380
rect -630 5360 -610 5380
rect -590 5360 -570 5380
rect -550 5360 -530 5380
rect -510 5360 -490 5380
rect -470 5360 -450 5380
rect -430 5360 -410 5380
rect -390 5360 -370 5380
rect -350 5360 -330 5380
rect -310 5360 -290 5380
rect -270 5360 -250 5380
rect -230 5360 -210 5380
rect -190 5360 -170 5380
rect -150 5360 -130 5380
rect -110 5360 -90 5380
rect -70 5360 -50 5380
rect -30 5360 -10 5380
rect 10 5360 30 5380
rect 50 5360 70 5380
rect 90 5360 110 5380
rect 130 5360 150 5380
rect 170 5360 190 5380
rect 210 5360 230 5380
rect 250 5360 270 5380
rect 290 5360 310 5380
rect 330 5360 350 5380
rect 370 5360 390 5380
rect 410 5360 440 5380
rect -5580 5265 -5550 5285
rect -5530 5265 -5510 5285
rect -5490 5265 -5470 5285
rect -5450 5265 -5430 5285
rect -5410 5265 -5390 5285
rect -5370 5265 -5350 5285
rect -5330 5265 -5310 5285
rect -5290 5265 -5270 5285
rect -5250 5265 -5230 5285
rect -5210 5265 -5190 5285
rect -5170 5265 -5150 5285
rect -5130 5265 -5110 5285
rect -5090 5265 -5070 5285
rect -5050 5265 -5030 5285
rect -5010 5265 -4990 5285
rect -4970 5265 -4950 5285
rect -4930 5265 -4910 5285
rect -4890 5265 -4870 5285
rect -4850 5265 -4830 5285
rect -4810 5265 -4790 5285
rect -4770 5265 -4750 5285
rect -4730 5265 -4710 5285
rect -4690 5265 -4670 5285
rect -4650 5265 -4630 5285
rect -4610 5265 -4590 5285
rect -4570 5265 -4550 5285
rect -4530 5265 -4510 5285
rect -4490 5265 -4470 5285
rect -4450 5265 -4430 5285
rect -4410 5265 -4390 5285
rect -4370 5265 -4350 5285
rect -4330 5265 -4310 5285
rect -4290 5265 -4270 5285
rect -4250 5265 -4230 5285
rect -4210 5265 -4190 5285
rect -4170 5265 -4150 5285
rect -4130 5265 -4110 5285
rect -4090 5265 -4070 5285
rect -4050 5265 -4030 5285
rect -4010 5265 -3990 5285
rect -3970 5265 -3950 5285
rect -3930 5265 -3910 5285
rect -3890 5265 -3870 5285
rect -3850 5265 -3830 5285
rect -3810 5265 -3790 5285
rect -3770 5265 -3750 5285
rect -3730 5265 -3710 5285
rect -3690 5265 -3670 5285
rect -3650 5265 -3630 5285
rect -3610 5265 -3590 5285
rect -3570 5265 -3550 5285
rect -3530 5265 -3510 5285
rect -3490 5265 -3470 5285
rect -3450 5265 -3430 5285
rect -3410 5265 -3390 5285
rect -3370 5265 -3350 5285
rect -3330 5265 -3310 5285
rect -3290 5265 -3270 5285
rect -3250 5265 -3230 5285
rect -3210 5265 -3190 5285
rect -3170 5265 -3150 5285
rect -3130 5265 -3110 5285
rect -2030 5265 -2010 5285
rect -1990 5265 -1970 5285
rect -1950 5265 -1930 5285
rect -1910 5265 -1890 5285
rect -1870 5265 -1850 5285
rect -1830 5265 -1810 5285
rect -1790 5265 -1770 5285
rect -1750 5265 -1730 5285
rect -1710 5265 -1690 5285
rect -1670 5265 -1650 5285
rect -1630 5265 -1610 5285
rect -1590 5265 -1570 5285
rect -1550 5265 -1530 5285
rect -1510 5265 -1490 5285
rect -1470 5265 -1450 5285
rect -1430 5265 -1410 5285
rect -1390 5265 -1370 5285
rect -1350 5265 -1330 5285
rect -1310 5265 -1290 5285
rect -1270 5265 -1250 5285
rect -1230 5265 -1210 5285
rect -1190 5265 -1170 5285
rect -1150 5265 -1130 5285
rect -1110 5265 -1090 5285
rect -1070 5265 -1050 5285
rect -1030 5265 -1010 5285
rect -990 5265 -970 5285
rect -950 5265 -930 5285
rect -910 5265 -890 5285
rect -870 5265 -850 5285
rect -830 5265 -810 5285
rect -790 5265 -770 5285
rect -750 5265 -730 5285
rect -710 5265 -690 5285
rect -670 5265 -650 5285
rect -630 5265 -610 5285
rect -590 5265 -570 5285
rect -550 5265 -530 5285
rect -510 5265 -490 5285
rect -470 5265 -450 5285
rect -430 5265 -410 5285
rect -390 5265 -370 5285
rect -350 5265 -330 5285
rect -310 5265 -290 5285
rect -270 5265 -250 5285
rect -230 5265 -210 5285
rect -190 5265 -170 5285
rect -150 5265 -130 5285
rect -110 5265 -90 5285
rect -70 5265 -50 5285
rect -30 5265 -10 5285
rect 10 5265 30 5285
rect 50 5265 70 5285
rect 90 5265 110 5285
rect 130 5265 150 5285
rect 170 5265 190 5285
rect 210 5265 230 5285
rect 250 5265 270 5285
rect 290 5265 310 5285
rect 330 5265 350 5285
rect 370 5265 390 5285
rect 410 5265 440 5285
rect -5580 5170 -5550 5190
rect -5530 5170 -5510 5190
rect -5490 5170 -5470 5190
rect -5450 5170 -5430 5190
rect -5410 5170 -5390 5190
rect -5370 5170 -5350 5190
rect -5330 5170 -5310 5190
rect -5290 5170 -5270 5190
rect -5250 5170 -5230 5190
rect -5210 5170 -5190 5190
rect -5170 5170 -5150 5190
rect -5130 5170 -5110 5190
rect -5090 5170 -5070 5190
rect -5050 5170 -5030 5190
rect -5010 5170 -4990 5190
rect -4970 5170 -4950 5190
rect -4930 5170 -4910 5190
rect -4890 5170 -4870 5190
rect -4850 5170 -4830 5190
rect -4810 5170 -4790 5190
rect -4770 5170 -4750 5190
rect -4730 5170 -4710 5190
rect -4690 5170 -4670 5190
rect -4650 5170 -4630 5190
rect -4610 5170 -4590 5190
rect -4570 5170 -4550 5190
rect -4530 5170 -4510 5190
rect -4490 5170 -4470 5190
rect -4450 5170 -4430 5190
rect -4410 5170 -4390 5190
rect -4370 5170 -4350 5190
rect -4330 5170 -4310 5190
rect -4290 5170 -4270 5190
rect -4250 5170 -4230 5190
rect -4210 5170 -4190 5190
rect -4170 5170 -4150 5190
rect -4130 5170 -4110 5190
rect -4090 5170 -4070 5190
rect -4050 5170 -4030 5190
rect -4010 5170 -3990 5190
rect -3970 5170 -3950 5190
rect -3930 5170 -3910 5190
rect -3890 5170 -3870 5190
rect -3850 5170 -3830 5190
rect -3810 5170 -3790 5190
rect -3770 5170 -3750 5190
rect -3730 5170 -3710 5190
rect -3690 5170 -3670 5190
rect -3650 5170 -3630 5190
rect -3610 5170 -3590 5190
rect -3570 5170 -3550 5190
rect -3530 5170 -3510 5190
rect -3490 5170 -3470 5190
rect -3450 5170 -3430 5190
rect -3410 5170 -3390 5190
rect -3370 5170 -3350 5190
rect -3330 5170 -3310 5190
rect -3290 5170 -3270 5190
rect -3250 5170 -3230 5190
rect -3210 5170 -3190 5190
rect -3170 5170 -3150 5190
rect -3130 5170 -3110 5190
rect -2030 5170 -2010 5190
rect -1990 5170 -1970 5190
rect -1950 5170 -1930 5190
rect -1910 5170 -1890 5190
rect -1870 5170 -1850 5190
rect -1830 5170 -1810 5190
rect -1790 5170 -1770 5190
rect -1750 5170 -1730 5190
rect -1710 5170 -1690 5190
rect -1670 5170 -1650 5190
rect -1630 5170 -1610 5190
rect -1590 5170 -1570 5190
rect -1550 5170 -1530 5190
rect -1510 5170 -1490 5190
rect -1470 5170 -1450 5190
rect -1430 5170 -1410 5190
rect -1390 5170 -1370 5190
rect -1350 5170 -1330 5190
rect -1310 5170 -1290 5190
rect -1270 5170 -1250 5190
rect -1230 5170 -1210 5190
rect -1190 5170 -1170 5190
rect -1150 5170 -1130 5190
rect -1110 5170 -1090 5190
rect -1070 5170 -1050 5190
rect -1030 5170 -1010 5190
rect -990 5170 -970 5190
rect -950 5170 -930 5190
rect -910 5170 -890 5190
rect -870 5170 -850 5190
rect -830 5170 -810 5190
rect -790 5170 -770 5190
rect -750 5170 -730 5190
rect -710 5170 -690 5190
rect -670 5170 -650 5190
rect -630 5170 -610 5190
rect -590 5170 -570 5190
rect -550 5170 -530 5190
rect -510 5170 -490 5190
rect -470 5170 -450 5190
rect -430 5170 -410 5190
rect -390 5170 -370 5190
rect -350 5170 -330 5190
rect -310 5170 -290 5190
rect -270 5170 -250 5190
rect -230 5170 -210 5190
rect -190 5170 -170 5190
rect -150 5170 -130 5190
rect -110 5170 -90 5190
rect -70 5170 -50 5190
rect -30 5170 -10 5190
rect 10 5170 30 5190
rect 50 5170 70 5190
rect 90 5170 110 5190
rect 130 5170 150 5190
rect 170 5170 190 5190
rect 210 5170 230 5190
rect 250 5170 270 5190
rect 290 5170 310 5190
rect 330 5170 350 5190
rect 370 5170 390 5190
rect 410 5170 440 5190
rect -5580 5075 -5550 5095
rect -5530 5075 -5510 5095
rect -5490 5075 -5470 5095
rect -5450 5075 -5430 5095
rect -5410 5075 -5390 5095
rect -5370 5075 -5350 5095
rect -5330 5075 -5310 5095
rect -5290 5075 -5270 5095
rect -5250 5075 -5230 5095
rect -5210 5075 -5190 5095
rect -5170 5075 -5150 5095
rect -5130 5075 -5110 5095
rect -5090 5075 -5070 5095
rect -5050 5075 -5030 5095
rect -5010 5075 -4990 5095
rect -4970 5075 -4950 5095
rect -4930 5075 -4910 5095
rect -4890 5075 -4870 5095
rect -4850 5075 -4830 5095
rect -4810 5075 -4790 5095
rect -4770 5075 -4750 5095
rect -4730 5075 -4710 5095
rect -4690 5075 -4670 5095
rect -4650 5075 -4630 5095
rect -4610 5075 -4590 5095
rect -4570 5075 -4550 5095
rect -4530 5075 -4510 5095
rect -4490 5075 -4470 5095
rect -4450 5075 -4430 5095
rect -4410 5075 -4390 5095
rect -4370 5075 -4350 5095
rect -4330 5075 -4310 5095
rect -4290 5075 -4270 5095
rect -4250 5075 -4230 5095
rect -4210 5075 -4190 5095
rect -4170 5075 -4150 5095
rect -4130 5075 -4110 5095
rect -4090 5075 -4070 5095
rect -4050 5075 -4030 5095
rect -4010 5075 -3990 5095
rect -3970 5075 -3950 5095
rect -3930 5075 -3910 5095
rect -3890 5075 -3870 5095
rect -3850 5075 -3830 5095
rect -3810 5075 -3790 5095
rect -3770 5075 -3750 5095
rect -3730 5075 -3710 5095
rect -3690 5075 -3670 5095
rect -3650 5075 -3630 5095
rect -3610 5075 -3590 5095
rect -3570 5075 -3550 5095
rect -3530 5075 -3510 5095
rect -3490 5075 -3470 5095
rect -3450 5075 -3430 5095
rect -3410 5075 -3390 5095
rect -3370 5075 -3350 5095
rect -3330 5075 -3310 5095
rect -3290 5075 -3270 5095
rect -3250 5075 -3230 5095
rect -3210 5075 -3190 5095
rect -3170 5075 -3150 5095
rect -3130 5075 -3110 5095
rect -2030 5075 -2010 5095
rect -1990 5075 -1970 5095
rect -1950 5075 -1930 5095
rect -1910 5075 -1890 5095
rect -1870 5075 -1850 5095
rect -1830 5075 -1810 5095
rect -1790 5075 -1770 5095
rect -1750 5075 -1730 5095
rect -1710 5075 -1690 5095
rect -1670 5075 -1650 5095
rect -1630 5075 -1610 5095
rect -1590 5075 -1570 5095
rect -1550 5075 -1530 5095
rect -1510 5075 -1490 5095
rect -1470 5075 -1450 5095
rect -1430 5075 -1410 5095
rect -1390 5075 -1370 5095
rect -1350 5075 -1330 5095
rect -1310 5075 -1290 5095
rect -1270 5075 -1250 5095
rect -1230 5075 -1210 5095
rect -1190 5075 -1170 5095
rect -1150 5075 -1130 5095
rect -1110 5075 -1090 5095
rect -1070 5075 -1050 5095
rect -1030 5075 -1010 5095
rect -990 5075 -970 5095
rect -950 5075 -930 5095
rect -910 5075 -890 5095
rect -870 5075 -850 5095
rect -830 5075 -810 5095
rect -790 5075 -770 5095
rect -750 5075 -730 5095
rect -710 5075 -690 5095
rect -670 5075 -650 5095
rect -630 5075 -610 5095
rect -590 5075 -570 5095
rect -550 5075 -530 5095
rect -510 5075 -490 5095
rect -470 5075 -450 5095
rect -430 5075 -410 5095
rect -390 5075 -370 5095
rect -350 5075 -330 5095
rect -310 5075 -290 5095
rect -270 5075 -250 5095
rect -230 5075 -210 5095
rect -190 5075 -170 5095
rect -150 5075 -130 5095
rect -110 5075 -90 5095
rect -70 5075 -50 5095
rect -30 5075 -10 5095
rect 10 5075 30 5095
rect 50 5075 70 5095
rect 90 5075 110 5095
rect 130 5075 150 5095
rect 170 5075 190 5095
rect 210 5075 230 5095
rect 250 5075 270 5095
rect 290 5075 310 5095
rect 330 5075 350 5095
rect 370 5075 390 5095
rect 410 5075 440 5095
rect -5580 4980 -5550 5000
rect -5530 4980 -5510 5000
rect -5490 4980 -5470 5000
rect -5450 4980 -5430 5000
rect -5410 4980 -5390 5000
rect -5370 4980 -5350 5000
rect -5330 4980 -5310 5000
rect -5290 4980 -5270 5000
rect -5250 4980 -5230 5000
rect -5210 4980 -5190 5000
rect -5170 4980 -5150 5000
rect -5130 4980 -5110 5000
rect -5090 4980 -5070 5000
rect -5050 4980 -5030 5000
rect -5010 4980 -4990 5000
rect -4970 4980 -4950 5000
rect -4930 4980 -4910 5000
rect -4890 4980 -4870 5000
rect -4850 4980 -4830 5000
rect -4810 4980 -4790 5000
rect -4770 4980 -4750 5000
rect -4730 4980 -4710 5000
rect -4690 4980 -4670 5000
rect -4650 4980 -4630 5000
rect -4610 4980 -4590 5000
rect -4570 4980 -4550 5000
rect -4530 4980 -4510 5000
rect -4490 4980 -4470 5000
rect -4450 4980 -4430 5000
rect -4410 4980 -4390 5000
rect -4370 4980 -4350 5000
rect -4330 4980 -4310 5000
rect -4290 4980 -4270 5000
rect -4250 4980 -4230 5000
rect -4210 4980 -4190 5000
rect -4170 4980 -4150 5000
rect -4130 4980 -4110 5000
rect -4090 4980 -4070 5000
rect -4050 4980 -4030 5000
rect -4010 4980 -3990 5000
rect -3970 4980 -3950 5000
rect -3930 4980 -3910 5000
rect -3890 4980 -3870 5000
rect -3850 4980 -3830 5000
rect -3810 4980 -3790 5000
rect -3770 4980 -3750 5000
rect -3730 4980 -3710 5000
rect -3690 4980 -3670 5000
rect -3650 4980 -3630 5000
rect -3610 4980 -3590 5000
rect -3570 4980 -3550 5000
rect -3530 4980 -3510 5000
rect -3490 4980 -3470 5000
rect -3450 4980 -3430 5000
rect -3410 4980 -3390 5000
rect -3370 4980 -3350 5000
rect -3330 4980 -3310 5000
rect -3290 4980 -3270 5000
rect -3250 4980 -3230 5000
rect -3210 4980 -3190 5000
rect -3170 4980 -3150 5000
rect -3130 4980 -3110 5000
rect -2030 4980 -2010 5000
rect -1990 4980 -1970 5000
rect -1950 4980 -1930 5000
rect -1910 4980 -1890 5000
rect -1870 4980 -1850 5000
rect -1830 4980 -1810 5000
rect -1790 4980 -1770 5000
rect -1750 4980 -1730 5000
rect -1710 4980 -1690 5000
rect -1670 4980 -1650 5000
rect -1630 4980 -1610 5000
rect -1590 4980 -1570 5000
rect -1550 4980 -1530 5000
rect -1510 4980 -1490 5000
rect -1470 4980 -1450 5000
rect -1430 4980 -1410 5000
rect -1390 4980 -1370 5000
rect -1350 4980 -1330 5000
rect -1310 4980 -1290 5000
rect -1270 4980 -1250 5000
rect -1230 4980 -1210 5000
rect -1190 4980 -1170 5000
rect -1150 4980 -1130 5000
rect -1110 4980 -1090 5000
rect -1070 4980 -1050 5000
rect -1030 4980 -1010 5000
rect -990 4980 -970 5000
rect -950 4980 -930 5000
rect -910 4980 -890 5000
rect -870 4980 -850 5000
rect -830 4980 -810 5000
rect -790 4980 -770 5000
rect -750 4980 -730 5000
rect -710 4980 -690 5000
rect -670 4980 -650 5000
rect -630 4980 -610 5000
rect -590 4980 -570 5000
rect -550 4980 -530 5000
rect -510 4980 -490 5000
rect -470 4980 -450 5000
rect -430 4980 -410 5000
rect -390 4980 -370 5000
rect -350 4980 -330 5000
rect -310 4980 -290 5000
rect -270 4980 -250 5000
rect -230 4980 -210 5000
rect -190 4980 -170 5000
rect -150 4980 -130 5000
rect -110 4980 -90 5000
rect -70 4980 -50 5000
rect -30 4980 -10 5000
rect 10 4980 30 5000
rect 50 4980 70 5000
rect 90 4980 110 5000
rect 130 4980 150 5000
rect 170 4980 190 5000
rect 210 4980 230 5000
rect 250 4980 270 5000
rect 290 4980 310 5000
rect 330 4980 350 5000
rect 370 4980 390 5000
rect 410 4980 440 5000
rect -5580 4885 -5550 4905
rect -5530 4885 -5510 4905
rect -5490 4885 -5470 4905
rect -5450 4885 -5430 4905
rect -5410 4885 -5390 4905
rect -5370 4885 -5350 4905
rect -5330 4885 -5310 4905
rect -5290 4885 -5270 4905
rect -5250 4885 -5230 4905
rect -5210 4885 -5190 4905
rect -5170 4885 -5150 4905
rect -5130 4885 -5110 4905
rect -5090 4885 -5070 4905
rect -5050 4885 -5030 4905
rect -5010 4885 -4990 4905
rect -4970 4885 -4950 4905
rect -4930 4885 -4910 4905
rect -4890 4885 -4870 4905
rect -4850 4885 -4830 4905
rect -4810 4885 -4790 4905
rect -4770 4885 -4750 4905
rect -4730 4885 -4710 4905
rect -4690 4885 -4670 4905
rect -4650 4885 -4630 4905
rect -4610 4885 -4590 4905
rect -4570 4885 -4550 4905
rect -4530 4885 -4510 4905
rect -4490 4885 -4470 4905
rect -4450 4885 -4430 4905
rect -4410 4885 -4390 4905
rect -4370 4885 -4350 4905
rect -4330 4885 -4310 4905
rect -4290 4885 -4270 4905
rect -4250 4885 -4230 4905
rect -4210 4885 -4190 4905
rect -4170 4885 -4150 4905
rect -4130 4885 -4110 4905
rect -4090 4885 -4070 4905
rect -4050 4885 -4030 4905
rect -4010 4885 -3990 4905
rect -3970 4885 -3950 4905
rect -3930 4885 -3910 4905
rect -3890 4885 -3870 4905
rect -3850 4885 -3830 4905
rect -3810 4885 -3790 4905
rect -3770 4885 -3750 4905
rect -3730 4885 -3710 4905
rect -3690 4885 -3670 4905
rect -3650 4885 -3630 4905
rect -3610 4885 -3590 4905
rect -3570 4885 -3550 4905
rect -3530 4885 -3510 4905
rect -3490 4885 -3470 4905
rect -3450 4885 -3430 4905
rect -3410 4885 -3390 4905
rect -3370 4885 -3350 4905
rect -3330 4885 -3310 4905
rect -3290 4885 -3270 4905
rect -3250 4885 -3230 4905
rect -3210 4885 -3190 4905
rect -3170 4885 -3150 4905
rect -3130 4885 -3110 4905
rect -2030 4885 -2010 4905
rect -1990 4885 -1970 4905
rect -1950 4885 -1930 4905
rect -1910 4885 -1890 4905
rect -1870 4885 -1850 4905
rect -1830 4885 -1810 4905
rect -1790 4885 -1770 4905
rect -1750 4885 -1730 4905
rect -1710 4885 -1690 4905
rect -1670 4885 -1650 4905
rect -1630 4885 -1610 4905
rect -1590 4885 -1570 4905
rect -1550 4885 -1530 4905
rect -1510 4885 -1490 4905
rect -1470 4885 -1450 4905
rect -1430 4885 -1410 4905
rect -1390 4885 -1370 4905
rect -1350 4885 -1330 4905
rect -1310 4885 -1290 4905
rect -1270 4885 -1250 4905
rect -1230 4885 -1210 4905
rect -1190 4885 -1170 4905
rect -1150 4885 -1130 4905
rect -1110 4885 -1090 4905
rect -1070 4885 -1050 4905
rect -1030 4885 -1010 4905
rect -990 4885 -970 4905
rect -950 4885 -930 4905
rect -910 4885 -890 4905
rect -870 4885 -850 4905
rect -830 4885 -810 4905
rect -790 4885 -770 4905
rect -750 4885 -730 4905
rect -710 4885 -690 4905
rect -670 4885 -650 4905
rect -630 4885 -610 4905
rect -590 4885 -570 4905
rect -550 4885 -530 4905
rect -510 4885 -490 4905
rect -470 4885 -450 4905
rect -430 4885 -410 4905
rect -390 4885 -370 4905
rect -350 4885 -330 4905
rect -310 4885 -290 4905
rect -270 4885 -250 4905
rect -230 4885 -210 4905
rect -190 4885 -170 4905
rect -150 4885 -130 4905
rect -110 4885 -90 4905
rect -70 4885 -50 4905
rect -30 4885 -10 4905
rect 10 4885 30 4905
rect 50 4885 70 4905
rect 90 4885 110 4905
rect 130 4885 150 4905
rect 170 4885 190 4905
rect 210 4885 230 4905
rect 250 4885 270 4905
rect 290 4885 310 4905
rect 330 4885 350 4905
rect 370 4885 390 4905
rect 410 4885 440 4905
rect -5580 4790 -5550 4810
rect -5530 4790 -5510 4810
rect -5490 4790 -5470 4810
rect -5450 4790 -5430 4810
rect -5410 4790 -5390 4810
rect -5370 4790 -5350 4810
rect -5330 4790 -5310 4810
rect -5290 4790 -5270 4810
rect -5250 4790 -5230 4810
rect -5210 4790 -5190 4810
rect -5170 4790 -5150 4810
rect -5130 4790 -5110 4810
rect -5090 4790 -5070 4810
rect -5050 4790 -5030 4810
rect -5010 4790 -4990 4810
rect -4970 4790 -4950 4810
rect -4930 4790 -4910 4810
rect -4890 4790 -4870 4810
rect -4850 4790 -4830 4810
rect -4810 4790 -4790 4810
rect -4770 4790 -4750 4810
rect -4730 4790 -4710 4810
rect -4690 4790 -4670 4810
rect -4650 4790 -4630 4810
rect -4610 4790 -4590 4810
rect -4570 4790 -4550 4810
rect -4530 4790 -4510 4810
rect -4490 4790 -4470 4810
rect -4450 4790 -4430 4810
rect -4410 4790 -4390 4810
rect -4370 4790 -4350 4810
rect -4330 4790 -4310 4810
rect -4290 4790 -4270 4810
rect -4250 4790 -4230 4810
rect -4210 4790 -4190 4810
rect -4170 4790 -4150 4810
rect -4130 4790 -4110 4810
rect -4090 4790 -4070 4810
rect -4050 4790 -4030 4810
rect -4010 4790 -3990 4810
rect -3970 4790 -3950 4810
rect -3930 4790 -3910 4810
rect -3890 4790 -3870 4810
rect -3850 4790 -3830 4810
rect -3810 4790 -3790 4810
rect -3770 4790 -3750 4810
rect -3730 4790 -3710 4810
rect -3690 4790 -3670 4810
rect -3650 4790 -3630 4810
rect -3610 4790 -3590 4810
rect -3570 4790 -3550 4810
rect -3530 4790 -3510 4810
rect -3490 4790 -3470 4810
rect -3450 4790 -3430 4810
rect -3410 4790 -3390 4810
rect -3370 4790 -3350 4810
rect -3330 4790 -3310 4810
rect -3290 4790 -3270 4810
rect -3250 4790 -3230 4810
rect -3210 4790 -3190 4810
rect -3170 4790 -3150 4810
rect -3130 4790 -3110 4810
rect -2030 4790 -2010 4810
rect -1990 4790 -1970 4810
rect -1950 4790 -1930 4810
rect -1910 4790 -1890 4810
rect -1870 4790 -1850 4810
rect -1830 4790 -1810 4810
rect -1790 4790 -1770 4810
rect -1750 4790 -1730 4810
rect -1710 4790 -1690 4810
rect -1670 4790 -1650 4810
rect -1630 4790 -1610 4810
rect -1590 4790 -1570 4810
rect -1550 4790 -1530 4810
rect -1510 4790 -1490 4810
rect -1470 4790 -1450 4810
rect -1430 4790 -1410 4810
rect -1390 4790 -1370 4810
rect -1350 4790 -1330 4810
rect -1310 4790 -1290 4810
rect -1270 4790 -1250 4810
rect -1230 4790 -1210 4810
rect -1190 4790 -1170 4810
rect -1150 4790 -1130 4810
rect -1110 4790 -1090 4810
rect -1070 4790 -1050 4810
rect -1030 4790 -1010 4810
rect -990 4790 -970 4810
rect -950 4790 -930 4810
rect -910 4790 -890 4810
rect -870 4790 -850 4810
rect -830 4790 -810 4810
rect -790 4790 -770 4810
rect -750 4790 -730 4810
rect -710 4790 -690 4810
rect -670 4790 -650 4810
rect -630 4790 -610 4810
rect -590 4790 -570 4810
rect -550 4790 -530 4810
rect -510 4790 -490 4810
rect -470 4790 -450 4810
rect -430 4790 -410 4810
rect -390 4790 -370 4810
rect -350 4790 -330 4810
rect -310 4790 -290 4810
rect -270 4790 -250 4810
rect -230 4790 -210 4810
rect -190 4790 -170 4810
rect -150 4790 -130 4810
rect -110 4790 -90 4810
rect -70 4790 -50 4810
rect -30 4790 -10 4810
rect 10 4790 30 4810
rect 50 4790 70 4810
rect 90 4790 110 4810
rect 130 4790 150 4810
rect 170 4790 190 4810
rect 210 4790 230 4810
rect 250 4790 270 4810
rect 290 4790 310 4810
rect 330 4790 350 4810
rect 370 4790 390 4810
rect 410 4790 440 4810
rect -5580 4695 -5550 4715
rect -5530 4695 -5510 4715
rect -5490 4695 -5470 4715
rect -5450 4695 -5430 4715
rect -5410 4695 -5390 4715
rect -5370 4695 -5350 4715
rect -5330 4695 -5310 4715
rect -5290 4695 -5270 4715
rect -5250 4695 -5230 4715
rect -5210 4695 -5190 4715
rect -5170 4695 -5150 4715
rect -5130 4695 -5110 4715
rect -5090 4695 -5070 4715
rect -5050 4695 -5030 4715
rect -5010 4695 -4990 4715
rect -4970 4695 -4950 4715
rect -4930 4695 -4910 4715
rect -4890 4695 -4870 4715
rect -4850 4695 -4830 4715
rect -4810 4695 -4790 4715
rect -4770 4695 -4750 4715
rect -4730 4695 -4710 4715
rect -4690 4695 -4670 4715
rect -4650 4695 -4630 4715
rect -4610 4695 -4590 4715
rect -4570 4695 -4550 4715
rect -4530 4695 -4510 4715
rect -4490 4695 -4470 4715
rect -4450 4695 -4430 4715
rect -4410 4695 -4390 4715
rect -4370 4695 -4350 4715
rect -4330 4695 -4310 4715
rect -4290 4695 -4270 4715
rect -4250 4695 -4230 4715
rect -4210 4695 -4190 4715
rect -4170 4695 -4150 4715
rect -4130 4695 -4110 4715
rect -4090 4695 -4070 4715
rect -4050 4695 -4030 4715
rect -4010 4695 -3990 4715
rect -3970 4695 -3950 4715
rect -3930 4695 -3910 4715
rect -3890 4695 -3870 4715
rect -3850 4695 -3830 4715
rect -3810 4695 -3790 4715
rect -3770 4695 -3750 4715
rect -3730 4695 -3710 4715
rect -3690 4695 -3670 4715
rect -3650 4695 -3630 4715
rect -3610 4695 -3590 4715
rect -3570 4695 -3550 4715
rect -3530 4695 -3510 4715
rect -3490 4695 -3470 4715
rect -3450 4695 -3430 4715
rect -3410 4695 -3390 4715
rect -3370 4695 -3350 4715
rect -3330 4695 -3310 4715
rect -3290 4695 -3270 4715
rect -3250 4695 -3230 4715
rect -3210 4695 -3190 4715
rect -3170 4695 -3150 4715
rect -3130 4695 -3110 4715
rect -2030 4695 -2010 4715
rect -1990 4695 -1970 4715
rect -1950 4695 -1930 4715
rect -1910 4695 -1890 4715
rect -1870 4695 -1850 4715
rect -1830 4695 -1810 4715
rect -1790 4695 -1770 4715
rect -1750 4695 -1730 4715
rect -1710 4695 -1690 4715
rect -1670 4695 -1650 4715
rect -1630 4695 -1610 4715
rect -1590 4695 -1570 4715
rect -1550 4695 -1530 4715
rect -1510 4695 -1490 4715
rect -1470 4695 -1450 4715
rect -1430 4695 -1410 4715
rect -1390 4695 -1370 4715
rect -1350 4695 -1330 4715
rect -1310 4695 -1290 4715
rect -1270 4695 -1250 4715
rect -1230 4695 -1210 4715
rect -1190 4695 -1170 4715
rect -1150 4695 -1130 4715
rect -1110 4695 -1090 4715
rect -1070 4695 -1050 4715
rect -1030 4695 -1010 4715
rect -990 4695 -970 4715
rect -950 4695 -930 4715
rect -910 4695 -890 4715
rect -870 4695 -850 4715
rect -830 4695 -810 4715
rect -790 4695 -770 4715
rect -750 4695 -730 4715
rect -710 4695 -690 4715
rect -670 4695 -650 4715
rect -630 4695 -610 4715
rect -590 4695 -570 4715
rect -550 4695 -530 4715
rect -510 4695 -490 4715
rect -470 4695 -450 4715
rect -430 4695 -410 4715
rect -390 4695 -370 4715
rect -350 4695 -330 4715
rect -310 4695 -290 4715
rect -270 4695 -250 4715
rect -230 4695 -210 4715
rect -190 4695 -170 4715
rect -150 4695 -130 4715
rect -110 4695 -90 4715
rect -70 4695 -50 4715
rect -30 4695 -10 4715
rect 10 4695 30 4715
rect 50 4695 70 4715
rect 90 4695 110 4715
rect 130 4695 150 4715
rect 170 4695 190 4715
rect 210 4695 230 4715
rect 250 4695 270 4715
rect 290 4695 310 4715
rect 330 4695 350 4715
rect 370 4695 390 4715
rect 410 4695 440 4715
rect -5580 4600 -5550 4620
rect -5530 4600 -5510 4620
rect -5490 4600 -5470 4620
rect -5450 4600 -5430 4620
rect -5410 4600 -5390 4620
rect -5370 4600 -5350 4620
rect -5330 4600 -5310 4620
rect -5290 4600 -5270 4620
rect -5250 4600 -5230 4620
rect -5210 4600 -5190 4620
rect -5170 4600 -5150 4620
rect -5130 4600 -5110 4620
rect -5090 4600 -5070 4620
rect -5050 4600 -5030 4620
rect -5010 4600 -4990 4620
rect -4970 4600 -4950 4620
rect -4930 4600 -4910 4620
rect -4890 4600 -4870 4620
rect -4850 4600 -4830 4620
rect -4810 4600 -4790 4620
rect -4770 4600 -4750 4620
rect -4730 4600 -4710 4620
rect -4690 4600 -4670 4620
rect -4650 4600 -4630 4620
rect -4610 4600 -4590 4620
rect -4570 4600 -4550 4620
rect -4530 4600 -4510 4620
rect -4490 4600 -4470 4620
rect -4450 4600 -4430 4620
rect -4410 4600 -4390 4620
rect -4370 4600 -4350 4620
rect -4330 4600 -4310 4620
rect -4290 4600 -4270 4620
rect -4250 4600 -4230 4620
rect -4210 4600 -4190 4620
rect -4170 4600 -4150 4620
rect -4130 4600 -4110 4620
rect -4090 4600 -4070 4620
rect -4050 4600 -4030 4620
rect -4010 4600 -3990 4620
rect -3970 4600 -3950 4620
rect -3930 4600 -3910 4620
rect -3890 4600 -3870 4620
rect -3850 4600 -3830 4620
rect -3810 4600 -3790 4620
rect -3770 4600 -3750 4620
rect -3730 4600 -3710 4620
rect -3690 4600 -3670 4620
rect -3650 4600 -3630 4620
rect -3610 4600 -3590 4620
rect -3570 4600 -3550 4620
rect -3530 4600 -3510 4620
rect -3490 4600 -3470 4620
rect -3450 4600 -3430 4620
rect -3410 4600 -3390 4620
rect -3370 4600 -3350 4620
rect -3330 4600 -3310 4620
rect -3290 4600 -3270 4620
rect -3250 4600 -3230 4620
rect -3210 4600 -3190 4620
rect -3170 4600 -3150 4620
rect -3130 4600 -3110 4620
rect -2030 4600 -2010 4620
rect -1990 4600 -1970 4620
rect -1950 4600 -1930 4620
rect -1910 4600 -1890 4620
rect -1870 4600 -1850 4620
rect -1830 4600 -1810 4620
rect -1790 4600 -1770 4620
rect -1750 4600 -1730 4620
rect -1710 4600 -1690 4620
rect -1670 4600 -1650 4620
rect -1630 4600 -1610 4620
rect -1590 4600 -1570 4620
rect -1550 4600 -1530 4620
rect -1510 4600 -1490 4620
rect -1470 4600 -1450 4620
rect -1430 4600 -1410 4620
rect -1390 4600 -1370 4620
rect -1350 4600 -1330 4620
rect -1310 4600 -1290 4620
rect -1270 4600 -1250 4620
rect -1230 4600 -1210 4620
rect -1190 4600 -1170 4620
rect -1150 4600 -1130 4620
rect -1110 4600 -1090 4620
rect -1070 4600 -1050 4620
rect -1030 4600 -1010 4620
rect -990 4600 -970 4620
rect -950 4600 -930 4620
rect -910 4600 -890 4620
rect -870 4600 -850 4620
rect -830 4600 -810 4620
rect -790 4600 -770 4620
rect -750 4600 -730 4620
rect -710 4600 -690 4620
rect -670 4600 -650 4620
rect -630 4600 -610 4620
rect -590 4600 -570 4620
rect -550 4600 -530 4620
rect -510 4600 -490 4620
rect -470 4600 -450 4620
rect -430 4600 -410 4620
rect -390 4600 -370 4620
rect -350 4600 -330 4620
rect -310 4600 -290 4620
rect -270 4600 -250 4620
rect -230 4600 -210 4620
rect -190 4600 -170 4620
rect -150 4600 -130 4620
rect -110 4600 -90 4620
rect -70 4600 -50 4620
rect -30 4600 -10 4620
rect 10 4600 30 4620
rect 50 4600 70 4620
rect 90 4600 110 4620
rect 130 4600 150 4620
rect 170 4600 190 4620
rect 210 4600 230 4620
rect 250 4600 270 4620
rect 290 4600 310 4620
rect 330 4600 350 4620
rect 370 4600 390 4620
rect 410 4600 440 4620
rect -5580 4505 -5550 4525
rect -5530 4505 -5510 4525
rect -5490 4505 -5470 4525
rect -5450 4505 -5430 4525
rect -5410 4505 -5390 4525
rect -5370 4505 -5350 4525
rect -5330 4505 -5310 4525
rect -5290 4505 -5270 4525
rect -5250 4505 -5230 4525
rect -5210 4505 -5190 4525
rect -5170 4505 -5150 4525
rect -5130 4505 -5110 4525
rect -5090 4505 -5070 4525
rect -5050 4505 -5030 4525
rect -5010 4505 -4990 4525
rect -4970 4505 -4950 4525
rect -4930 4505 -4910 4525
rect -4890 4505 -4870 4525
rect -4850 4505 -4830 4525
rect -4810 4505 -4790 4525
rect -4770 4505 -4750 4525
rect -4730 4505 -4710 4525
rect -4690 4505 -4670 4525
rect -4650 4505 -4630 4525
rect -4610 4505 -4590 4525
rect -4570 4505 -4550 4525
rect -4530 4505 -4510 4525
rect -4490 4505 -4470 4525
rect -4450 4505 -4430 4525
rect -4410 4505 -4390 4525
rect -4370 4505 -4350 4525
rect -4330 4505 -4310 4525
rect -4290 4505 -4270 4525
rect -4250 4505 -4230 4525
rect -4210 4505 -4190 4525
rect -4170 4505 -4150 4525
rect -4130 4505 -4110 4525
rect -4090 4505 -4070 4525
rect -4050 4505 -4030 4525
rect -4010 4505 -3990 4525
rect -3970 4505 -3950 4525
rect -3930 4505 -3910 4525
rect -3890 4505 -3870 4525
rect -3850 4505 -3830 4525
rect -3810 4505 -3790 4525
rect -3770 4505 -3750 4525
rect -3730 4505 -3710 4525
rect -3690 4505 -3670 4525
rect -3650 4505 -3630 4525
rect -3610 4505 -3590 4525
rect -3570 4505 -3550 4525
rect -3530 4505 -3510 4525
rect -3490 4505 -3470 4525
rect -3450 4505 -3430 4525
rect -3410 4505 -3390 4525
rect -3370 4505 -3350 4525
rect -3330 4505 -3310 4525
rect -3290 4505 -3270 4525
rect -3250 4505 -3230 4525
rect -3210 4505 -3190 4525
rect -3170 4505 -3150 4525
rect -3130 4505 -3110 4525
rect -2030 4505 -2010 4525
rect -1990 4505 -1970 4525
rect -1950 4505 -1930 4525
rect -1910 4505 -1890 4525
rect -1870 4505 -1850 4525
rect -1830 4505 -1810 4525
rect -1790 4505 -1770 4525
rect -1750 4505 -1730 4525
rect -1710 4505 -1690 4525
rect -1670 4505 -1650 4525
rect -1630 4505 -1610 4525
rect -1590 4505 -1570 4525
rect -1550 4505 -1530 4525
rect -1510 4505 -1490 4525
rect -1470 4505 -1450 4525
rect -1430 4505 -1410 4525
rect -1390 4505 -1370 4525
rect -1350 4505 -1330 4525
rect -1310 4505 -1290 4525
rect -1270 4505 -1250 4525
rect -1230 4505 -1210 4525
rect -1190 4505 -1170 4525
rect -1150 4505 -1130 4525
rect -1110 4505 -1090 4525
rect -1070 4505 -1050 4525
rect -1030 4505 -1010 4525
rect -990 4505 -970 4525
rect -950 4505 -930 4525
rect -910 4505 -890 4525
rect -870 4505 -850 4525
rect -830 4505 -810 4525
rect -790 4505 -770 4525
rect -750 4505 -730 4525
rect -710 4505 -690 4525
rect -670 4505 -650 4525
rect -630 4505 -610 4525
rect -590 4505 -570 4525
rect -550 4505 -530 4525
rect -510 4505 -490 4525
rect -470 4505 -450 4525
rect -430 4505 -410 4525
rect -390 4505 -370 4525
rect -350 4505 -330 4525
rect -310 4505 -290 4525
rect -270 4505 -250 4525
rect -230 4505 -210 4525
rect -190 4505 -170 4525
rect -150 4505 -130 4525
rect -110 4505 -90 4525
rect -70 4505 -50 4525
rect -30 4505 -10 4525
rect 10 4505 30 4525
rect 50 4505 70 4525
rect 90 4505 110 4525
rect 130 4505 150 4525
rect 170 4505 190 4525
rect 210 4505 230 4525
rect 250 4505 270 4525
rect 290 4505 310 4525
rect 330 4505 350 4525
rect 370 4505 390 4525
rect 410 4505 440 4525
rect -5580 4410 -5550 4430
rect -5530 4410 -5510 4430
rect -5490 4410 -5470 4430
rect -5450 4410 -5430 4430
rect -5410 4410 -5390 4430
rect -5370 4410 -5350 4430
rect -5330 4410 -5310 4430
rect -5290 4410 -5270 4430
rect -5250 4410 -5230 4430
rect -5210 4410 -5190 4430
rect -5170 4410 -5150 4430
rect -5130 4410 -5110 4430
rect -5090 4410 -5070 4430
rect -5050 4410 -5030 4430
rect -5010 4410 -4990 4430
rect -4970 4410 -4950 4430
rect -4930 4410 -4910 4430
rect -4890 4410 -4870 4430
rect -4850 4410 -4830 4430
rect -4810 4410 -4790 4430
rect -4770 4410 -4750 4430
rect -4730 4410 -4710 4430
rect -4690 4410 -4670 4430
rect -4650 4410 -4630 4430
rect -4610 4410 -4590 4430
rect -4570 4410 -4550 4430
rect -4530 4410 -4510 4430
rect -4490 4410 -4470 4430
rect -4450 4410 -4430 4430
rect -4410 4410 -4390 4430
rect -4370 4410 -4350 4430
rect -4330 4410 -4310 4430
rect -4290 4410 -4270 4430
rect -4250 4410 -4230 4430
rect -4210 4410 -4190 4430
rect -4170 4410 -4150 4430
rect -4130 4410 -4110 4430
rect -4090 4410 -4070 4430
rect -4050 4410 -4030 4430
rect -4010 4410 -3990 4430
rect -3970 4410 -3950 4430
rect -3930 4410 -3910 4430
rect -3890 4410 -3870 4430
rect -3850 4410 -3830 4430
rect -3810 4410 -3790 4430
rect -3770 4410 -3750 4430
rect -3730 4410 -3710 4430
rect -3690 4410 -3670 4430
rect -3650 4410 -3630 4430
rect -3610 4410 -3590 4430
rect -3570 4410 -3550 4430
rect -3530 4410 -3510 4430
rect -3490 4410 -3470 4430
rect -3450 4410 -3430 4430
rect -3410 4410 -3390 4430
rect -3370 4410 -3350 4430
rect -3330 4410 -3310 4430
rect -3290 4410 -3270 4430
rect -3250 4410 -3230 4430
rect -3210 4410 -3190 4430
rect -3170 4410 -3150 4430
rect -3130 4410 -3110 4430
rect -2030 4410 -2010 4430
rect -1990 4410 -1970 4430
rect -1950 4410 -1930 4430
rect -1910 4410 -1890 4430
rect -1870 4410 -1850 4430
rect -1830 4410 -1810 4430
rect -1790 4410 -1770 4430
rect -1750 4410 -1730 4430
rect -1710 4410 -1690 4430
rect -1670 4410 -1650 4430
rect -1630 4410 -1610 4430
rect -1590 4410 -1570 4430
rect -1550 4410 -1530 4430
rect -1510 4410 -1490 4430
rect -1470 4410 -1450 4430
rect -1430 4410 -1410 4430
rect -1390 4410 -1370 4430
rect -1350 4410 -1330 4430
rect -1310 4410 -1290 4430
rect -1270 4410 -1250 4430
rect -1230 4410 -1210 4430
rect -1190 4410 -1170 4430
rect -1150 4410 -1130 4430
rect -1110 4410 -1090 4430
rect -1070 4410 -1050 4430
rect -1030 4410 -1010 4430
rect -990 4410 -970 4430
rect -950 4410 -930 4430
rect -910 4410 -890 4430
rect -870 4410 -850 4430
rect -830 4410 -810 4430
rect -790 4410 -770 4430
rect -750 4410 -730 4430
rect -710 4410 -690 4430
rect -670 4410 -650 4430
rect -630 4410 -610 4430
rect -590 4410 -570 4430
rect -550 4410 -530 4430
rect -510 4410 -490 4430
rect -470 4410 -450 4430
rect -430 4410 -410 4430
rect -390 4410 -370 4430
rect -350 4410 -330 4430
rect -310 4410 -290 4430
rect -270 4410 -250 4430
rect -230 4410 -210 4430
rect -190 4410 -170 4430
rect -150 4410 -130 4430
rect -110 4410 -90 4430
rect -70 4410 -50 4430
rect -30 4410 -10 4430
rect 10 4410 30 4430
rect 50 4410 70 4430
rect 90 4410 110 4430
rect 130 4410 150 4430
rect 170 4410 190 4430
rect 210 4410 230 4430
rect 250 4410 270 4430
rect 290 4410 310 4430
rect 330 4410 350 4430
rect 370 4410 390 4430
rect 410 4410 440 4430
rect -5580 4315 -5550 4335
rect -5530 4315 -5510 4335
rect -5490 4315 -5470 4335
rect -5450 4315 -5430 4335
rect -5410 4315 -5390 4335
rect -5370 4315 -5350 4335
rect -5330 4315 -5310 4335
rect -5290 4315 -5270 4335
rect -5250 4315 -5230 4335
rect -5210 4315 -5190 4335
rect -5170 4315 -5150 4335
rect -5130 4315 -5110 4335
rect -5090 4315 -5070 4335
rect -5050 4315 -5030 4335
rect -5010 4315 -4990 4335
rect -4970 4315 -4950 4335
rect -4930 4315 -4910 4335
rect -4890 4315 -4870 4335
rect -4850 4315 -4830 4335
rect -4810 4315 -4790 4335
rect -4770 4315 -4750 4335
rect -4730 4315 -4710 4335
rect -4690 4315 -4670 4335
rect -4650 4315 -4630 4335
rect -4610 4315 -4590 4335
rect -4570 4315 -4550 4335
rect -4530 4315 -4510 4335
rect -4490 4315 -4470 4335
rect -4450 4315 -4430 4335
rect -4410 4315 -4390 4335
rect -4370 4315 -4350 4335
rect -4330 4315 -4310 4335
rect -4290 4315 -4270 4335
rect -4250 4315 -4230 4335
rect -4210 4315 -4190 4335
rect -4170 4315 -4150 4335
rect -4130 4315 -4110 4335
rect -4090 4315 -4070 4335
rect -4050 4315 -4030 4335
rect -4010 4315 -3990 4335
rect -3970 4315 -3950 4335
rect -3930 4315 -3910 4335
rect -3890 4315 -3870 4335
rect -3850 4315 -3830 4335
rect -3810 4315 -3790 4335
rect -3770 4315 -3750 4335
rect -3730 4315 -3710 4335
rect -3690 4315 -3670 4335
rect -3650 4315 -3630 4335
rect -3610 4315 -3590 4335
rect -3570 4315 -3550 4335
rect -3530 4315 -3510 4335
rect -3490 4315 -3470 4335
rect -3450 4315 -3430 4335
rect -3410 4315 -3390 4335
rect -3370 4315 -3350 4335
rect -3330 4315 -3310 4335
rect -3290 4315 -3270 4335
rect -3250 4315 -3230 4335
rect -3210 4315 -3190 4335
rect -3170 4315 -3150 4335
rect -3130 4315 -3110 4335
rect -2030 4315 -2010 4335
rect -1990 4315 -1970 4335
rect -1950 4315 -1930 4335
rect -1910 4315 -1890 4335
rect -1870 4315 -1850 4335
rect -1830 4315 -1810 4335
rect -1790 4315 -1770 4335
rect -1750 4315 -1730 4335
rect -1710 4315 -1690 4335
rect -1670 4315 -1650 4335
rect -1630 4315 -1610 4335
rect -1590 4315 -1570 4335
rect -1550 4315 -1530 4335
rect -1510 4315 -1490 4335
rect -1470 4315 -1450 4335
rect -1430 4315 -1410 4335
rect -1390 4315 -1370 4335
rect -1350 4315 -1330 4335
rect -1310 4315 -1290 4335
rect -1270 4315 -1250 4335
rect -1230 4315 -1210 4335
rect -1190 4315 -1170 4335
rect -1150 4315 -1130 4335
rect -1110 4315 -1090 4335
rect -1070 4315 -1050 4335
rect -1030 4315 -1010 4335
rect -990 4315 -970 4335
rect -950 4315 -930 4335
rect -910 4315 -890 4335
rect -870 4315 -850 4335
rect -830 4315 -810 4335
rect -790 4315 -770 4335
rect -750 4315 -730 4335
rect -710 4315 -690 4335
rect -670 4315 -650 4335
rect -630 4315 -610 4335
rect -590 4315 -570 4335
rect -550 4315 -530 4335
rect -510 4315 -490 4335
rect -470 4315 -450 4335
rect -430 4315 -410 4335
rect -390 4315 -370 4335
rect -350 4315 -330 4335
rect -310 4315 -290 4335
rect -270 4315 -250 4335
rect -230 4315 -210 4335
rect -190 4315 -170 4335
rect -150 4315 -130 4335
rect -110 4315 -90 4335
rect -70 4315 -50 4335
rect -30 4315 -10 4335
rect 10 4315 30 4335
rect 50 4315 70 4335
rect 90 4315 110 4335
rect 130 4315 150 4335
rect 170 4315 190 4335
rect 210 4315 230 4335
rect 250 4315 270 4335
rect 290 4315 310 4335
rect 330 4315 350 4335
rect 370 4315 390 4335
rect 410 4315 440 4335
rect -5580 4220 -5550 4240
rect -5530 4220 -5510 4240
rect -5490 4220 -5470 4240
rect -5450 4220 -5430 4240
rect -5410 4220 -5390 4240
rect -5370 4220 -5350 4240
rect -5330 4220 -5310 4240
rect -5290 4220 -5270 4240
rect -5250 4220 -5230 4240
rect -5210 4220 -5190 4240
rect -5170 4220 -5150 4240
rect -5130 4220 -5110 4240
rect -5090 4220 -5070 4240
rect -5050 4220 -5030 4240
rect -5010 4220 -4990 4240
rect -4970 4220 -4950 4240
rect -4930 4220 -4910 4240
rect -4890 4220 -4870 4240
rect -4850 4220 -4830 4240
rect -4810 4220 -4790 4240
rect -4770 4220 -4750 4240
rect -4730 4220 -4710 4240
rect -4690 4220 -4670 4240
rect -4650 4220 -4630 4240
rect -4610 4220 -4590 4240
rect -4570 4220 -4550 4240
rect -4530 4220 -4510 4240
rect -4490 4220 -4470 4240
rect -4450 4220 -4430 4240
rect -4410 4220 -4390 4240
rect -4370 4220 -4350 4240
rect -4330 4220 -4310 4240
rect -4290 4220 -4270 4240
rect -4250 4220 -4230 4240
rect -4210 4220 -4190 4240
rect -4170 4220 -4150 4240
rect -4130 4220 -4110 4240
rect -4090 4220 -4070 4240
rect -4050 4220 -4030 4240
rect -4010 4220 -3990 4240
rect -3970 4220 -3950 4240
rect -3930 4220 -3910 4240
rect -3890 4220 -3870 4240
rect -3850 4220 -3830 4240
rect -3810 4220 -3790 4240
rect -3770 4220 -3750 4240
rect -3730 4220 -3710 4240
rect -3690 4220 -3670 4240
rect -3650 4220 -3630 4240
rect -3610 4220 -3590 4240
rect -3570 4220 -3550 4240
rect -3530 4220 -3510 4240
rect -3490 4220 -3470 4240
rect -3450 4220 -3430 4240
rect -3410 4220 -3390 4240
rect -3370 4220 -3350 4240
rect -3330 4220 -3310 4240
rect -3290 4220 -3270 4240
rect -3250 4220 -3230 4240
rect -3210 4220 -3190 4240
rect -3170 4220 -3150 4240
rect -3130 4220 -3110 4240
rect -2030 4220 -2010 4240
rect -1990 4220 -1970 4240
rect -1950 4220 -1930 4240
rect -1910 4220 -1890 4240
rect -1870 4220 -1850 4240
rect -1830 4220 -1810 4240
rect -1790 4220 -1770 4240
rect -1750 4220 -1730 4240
rect -1710 4220 -1690 4240
rect -1670 4220 -1650 4240
rect -1630 4220 -1610 4240
rect -1590 4220 -1570 4240
rect -1550 4220 -1530 4240
rect -1510 4220 -1490 4240
rect -1470 4220 -1450 4240
rect -1430 4220 -1410 4240
rect -1390 4220 -1370 4240
rect -1350 4220 -1330 4240
rect -1310 4220 -1290 4240
rect -1270 4220 -1250 4240
rect -1230 4220 -1210 4240
rect -1190 4220 -1170 4240
rect -1150 4220 -1130 4240
rect -1110 4220 -1090 4240
rect -1070 4220 -1050 4240
rect -1030 4220 -1010 4240
rect -990 4220 -970 4240
rect -950 4220 -930 4240
rect -910 4220 -890 4240
rect -870 4220 -850 4240
rect -830 4220 -810 4240
rect -790 4220 -770 4240
rect -750 4220 -730 4240
rect -710 4220 -690 4240
rect -670 4220 -650 4240
rect -630 4220 -610 4240
rect -590 4220 -570 4240
rect -550 4220 -530 4240
rect -510 4220 -490 4240
rect -470 4220 -450 4240
rect -430 4220 -410 4240
rect -390 4220 -370 4240
rect -350 4220 -330 4240
rect -310 4220 -290 4240
rect -270 4220 -250 4240
rect -230 4220 -210 4240
rect -190 4220 -170 4240
rect -150 4220 -130 4240
rect -110 4220 -90 4240
rect -70 4220 -50 4240
rect -30 4220 -10 4240
rect 10 4220 30 4240
rect 50 4220 70 4240
rect 90 4220 110 4240
rect 130 4220 150 4240
rect 170 4220 190 4240
rect 210 4220 230 4240
rect 250 4220 270 4240
rect 290 4220 310 4240
rect 330 4220 350 4240
rect 370 4220 390 4240
rect 410 4220 440 4240
rect -5580 4125 -5550 4145
rect -5530 4125 -5510 4145
rect -5490 4125 -5470 4145
rect -5450 4125 -5430 4145
rect -5410 4125 -5390 4145
rect -5370 4125 -5350 4145
rect -5330 4125 -5310 4145
rect -5290 4125 -5270 4145
rect -5250 4125 -5230 4145
rect -5210 4125 -5190 4145
rect -5170 4125 -5150 4145
rect -5130 4125 -5110 4145
rect -5090 4125 -5070 4145
rect -5050 4125 -5030 4145
rect -5010 4125 -4990 4145
rect -4970 4125 -4950 4145
rect -4930 4125 -4910 4145
rect -4890 4125 -4870 4145
rect -4850 4125 -4830 4145
rect -4810 4125 -4790 4145
rect -4770 4125 -4750 4145
rect -4730 4125 -4710 4145
rect -4690 4125 -4670 4145
rect -4650 4125 -4630 4145
rect -4610 4125 -4590 4145
rect -4570 4125 -4550 4145
rect -4530 4125 -4510 4145
rect -4490 4125 -4470 4145
rect -4450 4125 -4430 4145
rect -4410 4125 -4390 4145
rect -4370 4125 -4350 4145
rect -4330 4125 -4310 4145
rect -4290 4125 -4270 4145
rect -4250 4125 -4230 4145
rect -4210 4125 -4190 4145
rect -4170 4125 -4150 4145
rect -4130 4125 -4110 4145
rect -4090 4125 -4070 4145
rect -4050 4125 -4030 4145
rect -4010 4125 -3990 4145
rect -3970 4125 -3950 4145
rect -3930 4125 -3910 4145
rect -3890 4125 -3870 4145
rect -3850 4125 -3830 4145
rect -3810 4125 -3790 4145
rect -3770 4125 -3750 4145
rect -3730 4125 -3710 4145
rect -3690 4125 -3670 4145
rect -3650 4125 -3630 4145
rect -3610 4125 -3590 4145
rect -3570 4125 -3550 4145
rect -3530 4125 -3510 4145
rect -3490 4125 -3470 4145
rect -3450 4125 -3430 4145
rect -3410 4125 -3390 4145
rect -3370 4125 -3350 4145
rect -3330 4125 -3310 4145
rect -3290 4125 -3270 4145
rect -3250 4125 -3230 4145
rect -3210 4125 -3190 4145
rect -3170 4125 -3150 4145
rect -3130 4125 -3110 4145
rect -2030 4125 -2010 4145
rect -1990 4125 -1970 4145
rect -1950 4125 -1930 4145
rect -1910 4125 -1890 4145
rect -1870 4125 -1850 4145
rect -1830 4125 -1810 4145
rect -1790 4125 -1770 4145
rect -1750 4125 -1730 4145
rect -1710 4125 -1690 4145
rect -1670 4125 -1650 4145
rect -1630 4125 -1610 4145
rect -1590 4125 -1570 4145
rect -1550 4125 -1530 4145
rect -1510 4125 -1490 4145
rect -1470 4125 -1450 4145
rect -1430 4125 -1410 4145
rect -1390 4125 -1370 4145
rect -1350 4125 -1330 4145
rect -1310 4125 -1290 4145
rect -1270 4125 -1250 4145
rect -1230 4125 -1210 4145
rect -1190 4125 -1170 4145
rect -1150 4125 -1130 4145
rect -1110 4125 -1090 4145
rect -1070 4125 -1050 4145
rect -1030 4125 -1010 4145
rect -990 4125 -970 4145
rect -950 4125 -930 4145
rect -910 4125 -890 4145
rect -870 4125 -850 4145
rect -830 4125 -810 4145
rect -790 4125 -770 4145
rect -750 4125 -730 4145
rect -710 4125 -690 4145
rect -670 4125 -650 4145
rect -630 4125 -610 4145
rect -590 4125 -570 4145
rect -550 4125 -530 4145
rect -510 4125 -490 4145
rect -470 4125 -450 4145
rect -430 4125 -410 4145
rect -390 4125 -370 4145
rect -350 4125 -330 4145
rect -310 4125 -290 4145
rect -270 4125 -250 4145
rect -230 4125 -210 4145
rect -190 4125 -170 4145
rect -150 4125 -130 4145
rect -110 4125 -90 4145
rect -70 4125 -50 4145
rect -30 4125 -10 4145
rect 10 4125 30 4145
rect 50 4125 70 4145
rect 90 4125 110 4145
rect 130 4125 150 4145
rect 170 4125 190 4145
rect 210 4125 230 4145
rect 250 4125 270 4145
rect 290 4125 310 4145
rect 330 4125 350 4145
rect 370 4125 390 4145
rect 410 4125 440 4145
rect -5580 4030 -5550 4050
rect -5530 4030 -5510 4050
rect -5490 4030 -5470 4050
rect -5450 4030 -5430 4050
rect -5410 4030 -5390 4050
rect -5370 4030 -5350 4050
rect -5330 4030 -5310 4050
rect -5290 4030 -5270 4050
rect -5250 4030 -5230 4050
rect -5210 4030 -5190 4050
rect -5170 4030 -5150 4050
rect -5130 4030 -5110 4050
rect -5090 4030 -5070 4050
rect -5050 4030 -5030 4050
rect -5010 4030 -4990 4050
rect -4970 4030 -4950 4050
rect -4930 4030 -4910 4050
rect -4890 4030 -4870 4050
rect -4850 4030 -4830 4050
rect -4810 4030 -4790 4050
rect -4770 4030 -4750 4050
rect -4730 4030 -4710 4050
rect -4690 4030 -4670 4050
rect -4650 4030 -4630 4050
rect -4610 4030 -4590 4050
rect -4570 4030 -4550 4050
rect -4530 4030 -4510 4050
rect -4490 4030 -4470 4050
rect -4450 4030 -4430 4050
rect -4410 4030 -4390 4050
rect -4370 4030 -4350 4050
rect -4330 4030 -4310 4050
rect -4290 4030 -4270 4050
rect -4250 4030 -4230 4050
rect -4210 4030 -4190 4050
rect -4170 4030 -4150 4050
rect -4130 4030 -4110 4050
rect -4090 4030 -4070 4050
rect -4050 4030 -4030 4050
rect -4010 4030 -3990 4050
rect -3970 4030 -3950 4050
rect -3930 4030 -3910 4050
rect -3890 4030 -3870 4050
rect -3850 4030 -3830 4050
rect -3810 4030 -3790 4050
rect -3770 4030 -3750 4050
rect -3730 4030 -3710 4050
rect -3690 4030 -3670 4050
rect -3650 4030 -3630 4050
rect -3610 4030 -3590 4050
rect -3570 4030 -3550 4050
rect -3530 4030 -3510 4050
rect -3490 4030 -3470 4050
rect -3450 4030 -3430 4050
rect -3410 4030 -3390 4050
rect -3370 4030 -3350 4050
rect -3330 4030 -3310 4050
rect -3290 4030 -3270 4050
rect -3250 4030 -3230 4050
rect -3210 4030 -3190 4050
rect -3170 4030 -3150 4050
rect -3130 4030 -3110 4050
rect -2030 4030 -2010 4050
rect -1990 4030 -1970 4050
rect -1950 4030 -1930 4050
rect -1910 4030 -1890 4050
rect -1870 4030 -1850 4050
rect -1830 4030 -1810 4050
rect -1790 4030 -1770 4050
rect -1750 4030 -1730 4050
rect -1710 4030 -1690 4050
rect -1670 4030 -1650 4050
rect -1630 4030 -1610 4050
rect -1590 4030 -1570 4050
rect -1550 4030 -1530 4050
rect -1510 4030 -1490 4050
rect -1470 4030 -1450 4050
rect -1430 4030 -1410 4050
rect -1390 4030 -1370 4050
rect -1350 4030 -1330 4050
rect -1310 4030 -1290 4050
rect -1270 4030 -1250 4050
rect -1230 4030 -1210 4050
rect -1190 4030 -1170 4050
rect -1150 4030 -1130 4050
rect -1110 4030 -1090 4050
rect -1070 4030 -1050 4050
rect -1030 4030 -1010 4050
rect -990 4030 -970 4050
rect -950 4030 -930 4050
rect -910 4030 -890 4050
rect -870 4030 -850 4050
rect -830 4030 -810 4050
rect -790 4030 -770 4050
rect -750 4030 -730 4050
rect -710 4030 -690 4050
rect -670 4030 -650 4050
rect -630 4030 -610 4050
rect -590 4030 -570 4050
rect -550 4030 -530 4050
rect -510 4030 -490 4050
rect -470 4030 -450 4050
rect -430 4030 -410 4050
rect -390 4030 -370 4050
rect -350 4030 -330 4050
rect -310 4030 -290 4050
rect -270 4030 -250 4050
rect -230 4030 -210 4050
rect -190 4030 -170 4050
rect -150 4030 -130 4050
rect -110 4030 -90 4050
rect -70 4030 -50 4050
rect -30 4030 -10 4050
rect 10 4030 30 4050
rect 50 4030 70 4050
rect 90 4030 110 4050
rect 130 4030 150 4050
rect 170 4030 190 4050
rect 210 4030 230 4050
rect 250 4030 270 4050
rect 290 4030 310 4050
rect 330 4030 350 4050
rect 370 4030 390 4050
rect 410 4030 440 4050
rect -5580 3935 -5550 3955
rect -5530 3935 -5510 3955
rect -5490 3935 -5470 3955
rect -5450 3935 -5430 3955
rect -5410 3935 -5390 3955
rect -5370 3935 -5350 3955
rect -5330 3935 -5310 3955
rect -5290 3935 -5270 3955
rect -5250 3935 -5230 3955
rect -5210 3935 -5190 3955
rect -5170 3935 -5150 3955
rect -5130 3935 -5110 3955
rect -5090 3935 -5070 3955
rect -5050 3935 -5030 3955
rect -5010 3935 -4990 3955
rect -4970 3935 -4950 3955
rect -4930 3935 -4910 3955
rect -4890 3935 -4870 3955
rect -4850 3935 -4830 3955
rect -4810 3935 -4790 3955
rect -4770 3935 -4750 3955
rect -4730 3935 -4710 3955
rect -4690 3935 -4670 3955
rect -4650 3935 -4630 3955
rect -4610 3935 -4590 3955
rect -4570 3935 -4550 3955
rect -4530 3935 -4510 3955
rect -4490 3935 -4470 3955
rect -4450 3935 -4430 3955
rect -4410 3935 -4390 3955
rect -4370 3935 -4350 3955
rect -4330 3935 -4310 3955
rect -4290 3935 -4270 3955
rect -4250 3935 -4230 3955
rect -4210 3935 -4190 3955
rect -4170 3935 -4150 3955
rect -4130 3935 -4110 3955
rect -4090 3935 -4070 3955
rect -4050 3935 -4030 3955
rect -4010 3935 -3990 3955
rect -3970 3935 -3950 3955
rect -3930 3935 -3910 3955
rect -3890 3935 -3870 3955
rect -3850 3935 -3830 3955
rect -3810 3935 -3790 3955
rect -3770 3935 -3750 3955
rect -3730 3935 -3710 3955
rect -3690 3935 -3670 3955
rect -3650 3935 -3630 3955
rect -3610 3935 -3590 3955
rect -3570 3935 -3550 3955
rect -3530 3935 -3510 3955
rect -3490 3935 -3470 3955
rect -3450 3935 -3430 3955
rect -3410 3935 -3390 3955
rect -3370 3935 -3350 3955
rect -3330 3935 -3310 3955
rect -3290 3935 -3270 3955
rect -3250 3935 -3230 3955
rect -3210 3935 -3190 3955
rect -3170 3935 -3150 3955
rect -3130 3935 -3110 3955
rect -2030 3935 -2010 3955
rect -1990 3935 -1970 3955
rect -1950 3935 -1930 3955
rect -1910 3935 -1890 3955
rect -1870 3935 -1850 3955
rect -1830 3935 -1810 3955
rect -1790 3935 -1770 3955
rect -1750 3935 -1730 3955
rect -1710 3935 -1690 3955
rect -1670 3935 -1650 3955
rect -1630 3935 -1610 3955
rect -1590 3935 -1570 3955
rect -1550 3935 -1530 3955
rect -1510 3935 -1490 3955
rect -1470 3935 -1450 3955
rect -1430 3935 -1410 3955
rect -1390 3935 -1370 3955
rect -1350 3935 -1330 3955
rect -1310 3935 -1290 3955
rect -1270 3935 -1250 3955
rect -1230 3935 -1210 3955
rect -1190 3935 -1170 3955
rect -1150 3935 -1130 3955
rect -1110 3935 -1090 3955
rect -1070 3935 -1050 3955
rect -1030 3935 -1010 3955
rect -990 3935 -970 3955
rect -950 3935 -930 3955
rect -910 3935 -890 3955
rect -870 3935 -850 3955
rect -830 3935 -810 3955
rect -790 3935 -770 3955
rect -750 3935 -730 3955
rect -710 3935 -690 3955
rect -670 3935 -650 3955
rect -630 3935 -610 3955
rect -590 3935 -570 3955
rect -550 3935 -530 3955
rect -510 3935 -490 3955
rect -470 3935 -450 3955
rect -430 3935 -410 3955
rect -390 3935 -370 3955
rect -350 3935 -330 3955
rect -310 3935 -290 3955
rect -270 3935 -250 3955
rect -230 3935 -210 3955
rect -190 3935 -170 3955
rect -150 3935 -130 3955
rect -110 3935 -90 3955
rect -70 3935 -50 3955
rect -30 3935 -10 3955
rect 10 3935 30 3955
rect 50 3935 70 3955
rect 90 3935 110 3955
rect 130 3935 150 3955
rect 170 3935 190 3955
rect 210 3935 230 3955
rect 250 3935 270 3955
rect 290 3935 310 3955
rect 330 3935 350 3955
rect 370 3935 390 3955
rect 410 3935 440 3955
rect -5580 3840 -5550 3860
rect -5530 3840 -5510 3860
rect -5490 3840 -5470 3860
rect -5450 3840 -5430 3860
rect -5410 3840 -5390 3860
rect -5370 3840 -5350 3860
rect -5330 3840 -5310 3860
rect -5290 3840 -5270 3860
rect -5250 3840 -5230 3860
rect -5210 3840 -5190 3860
rect -5170 3840 -5150 3860
rect -5130 3840 -5110 3860
rect -5090 3840 -5070 3860
rect -5050 3840 -5030 3860
rect -5010 3840 -4990 3860
rect -4970 3840 -4950 3860
rect -4930 3840 -4910 3860
rect -4890 3840 -4870 3860
rect -4850 3840 -4830 3860
rect -4810 3840 -4790 3860
rect -4770 3840 -4750 3860
rect -4730 3840 -4710 3860
rect -4690 3840 -4670 3860
rect -4650 3840 -4630 3860
rect -4610 3840 -4590 3860
rect -4570 3840 -4550 3860
rect -4530 3840 -4510 3860
rect -4490 3840 -4470 3860
rect -4450 3840 -4430 3860
rect -4410 3840 -4390 3860
rect -4370 3840 -4350 3860
rect -4330 3840 -4310 3860
rect -4290 3840 -4270 3860
rect -4250 3840 -4230 3860
rect -4210 3840 -4190 3860
rect -4170 3840 -4150 3860
rect -4130 3840 -4110 3860
rect -4090 3840 -4070 3860
rect -4050 3840 -4030 3860
rect -4010 3840 -3990 3860
rect -3970 3840 -3950 3860
rect -3930 3840 -3910 3860
rect -3890 3840 -3870 3860
rect -3850 3840 -3830 3860
rect -3810 3840 -3790 3860
rect -3770 3840 -3750 3860
rect -3730 3840 -3710 3860
rect -3690 3840 -3670 3860
rect -3650 3840 -3630 3860
rect -3610 3840 -3590 3860
rect -3570 3840 -3550 3860
rect -3530 3840 -3510 3860
rect -3490 3840 -3470 3860
rect -3450 3840 -3430 3860
rect -3410 3840 -3390 3860
rect -3370 3840 -3350 3860
rect -3330 3840 -3310 3860
rect -3290 3840 -3270 3860
rect -3250 3840 -3230 3860
rect -3210 3840 -3190 3860
rect -3170 3840 -3150 3860
rect -3130 3840 -3110 3860
rect -2030 3840 -2010 3860
rect -1990 3840 -1970 3860
rect -1950 3840 -1930 3860
rect -1910 3840 -1890 3860
rect -1870 3840 -1850 3860
rect -1830 3840 -1810 3860
rect -1790 3840 -1770 3860
rect -1750 3840 -1730 3860
rect -1710 3840 -1690 3860
rect -1670 3840 -1650 3860
rect -1630 3840 -1610 3860
rect -1590 3840 -1570 3860
rect -1550 3840 -1530 3860
rect -1510 3840 -1490 3860
rect -1470 3840 -1450 3860
rect -1430 3840 -1410 3860
rect -1390 3840 -1370 3860
rect -1350 3840 -1330 3860
rect -1310 3840 -1290 3860
rect -1270 3840 -1250 3860
rect -1230 3840 -1210 3860
rect -1190 3840 -1170 3860
rect -1150 3840 -1130 3860
rect -1110 3840 -1090 3860
rect -1070 3840 -1050 3860
rect -1030 3840 -1010 3860
rect -990 3840 -970 3860
rect -950 3840 -930 3860
rect -910 3840 -890 3860
rect -870 3840 -850 3860
rect -830 3840 -810 3860
rect -790 3840 -770 3860
rect -750 3840 -730 3860
rect -710 3840 -690 3860
rect -670 3840 -650 3860
rect -630 3840 -610 3860
rect -590 3840 -570 3860
rect -550 3840 -530 3860
rect -510 3840 -490 3860
rect -470 3840 -450 3860
rect -430 3840 -410 3860
rect -390 3840 -370 3860
rect -350 3840 -330 3860
rect -310 3840 -290 3860
rect -270 3840 -250 3860
rect -230 3840 -210 3860
rect -190 3840 -170 3860
rect -150 3840 -130 3860
rect -110 3840 -90 3860
rect -70 3840 -50 3860
rect -30 3840 -10 3860
rect 10 3840 30 3860
rect 50 3840 70 3860
rect 90 3840 110 3860
rect 130 3840 150 3860
rect 170 3840 190 3860
rect 210 3840 230 3860
rect 250 3840 270 3860
rect 290 3840 310 3860
rect 330 3840 350 3860
rect 370 3840 390 3860
rect 410 3840 440 3860
rect -5580 3745 -5550 3765
rect -5530 3745 -5510 3765
rect -5490 3745 -5470 3765
rect -5450 3745 -5430 3765
rect -5410 3745 -5390 3765
rect -5370 3745 -5350 3765
rect -5330 3745 -5310 3765
rect -5290 3745 -5270 3765
rect -5250 3745 -5230 3765
rect -5210 3745 -5190 3765
rect -5170 3745 -5150 3765
rect -5130 3745 -5110 3765
rect -5090 3745 -5070 3765
rect -5050 3745 -5030 3765
rect -5010 3745 -4990 3765
rect -4970 3745 -4950 3765
rect -4930 3745 -4910 3765
rect -4890 3745 -4870 3765
rect -4850 3745 -4830 3765
rect -4810 3745 -4790 3765
rect -4770 3745 -4750 3765
rect -4730 3745 -4710 3765
rect -4690 3745 -4670 3765
rect -4650 3745 -4630 3765
rect -4610 3745 -4590 3765
rect -4570 3745 -4550 3765
rect -4530 3745 -4510 3765
rect -4490 3745 -4470 3765
rect -4450 3745 -4430 3765
rect -4410 3745 -4390 3765
rect -4370 3745 -4350 3765
rect -4330 3745 -4310 3765
rect -4290 3745 -4270 3765
rect -4250 3745 -4230 3765
rect -4210 3745 -4190 3765
rect -4170 3745 -4150 3765
rect -4130 3745 -4110 3765
rect -4090 3745 -4070 3765
rect -4050 3745 -4030 3765
rect -4010 3745 -3990 3765
rect -3970 3745 -3950 3765
rect -3930 3745 -3910 3765
rect -3890 3745 -3870 3765
rect -3850 3745 -3830 3765
rect -3810 3745 -3790 3765
rect -3770 3745 -3750 3765
rect -3730 3745 -3710 3765
rect -3690 3745 -3670 3765
rect -3650 3745 -3630 3765
rect -3610 3745 -3590 3765
rect -3570 3745 -3550 3765
rect -3530 3745 -3510 3765
rect -3490 3745 -3470 3765
rect -3450 3745 -3430 3765
rect -3410 3745 -3390 3765
rect -3370 3745 -3350 3765
rect -3330 3745 -3310 3765
rect -3290 3745 -3270 3765
rect -3250 3745 -3230 3765
rect -3210 3745 -3190 3765
rect -3170 3745 -3150 3765
rect -3130 3745 -3110 3765
rect -2030 3745 -2010 3765
rect -1990 3745 -1970 3765
rect -1950 3745 -1930 3765
rect -1910 3745 -1890 3765
rect -1870 3745 -1850 3765
rect -1830 3745 -1810 3765
rect -1790 3745 -1770 3765
rect -1750 3745 -1730 3765
rect -1710 3745 -1690 3765
rect -1670 3745 -1650 3765
rect -1630 3745 -1610 3765
rect -1590 3745 -1570 3765
rect -1550 3745 -1530 3765
rect -1510 3745 -1490 3765
rect -1470 3745 -1450 3765
rect -1430 3745 -1410 3765
rect -1390 3745 -1370 3765
rect -1350 3745 -1330 3765
rect -1310 3745 -1290 3765
rect -1270 3745 -1250 3765
rect -1230 3745 -1210 3765
rect -1190 3745 -1170 3765
rect -1150 3745 -1130 3765
rect -1110 3745 -1090 3765
rect -1070 3745 -1050 3765
rect -1030 3745 -1010 3765
rect -990 3745 -970 3765
rect -950 3745 -930 3765
rect -910 3745 -890 3765
rect -870 3745 -850 3765
rect -830 3745 -810 3765
rect -790 3745 -770 3765
rect -750 3745 -730 3765
rect -710 3745 -690 3765
rect -670 3745 -650 3765
rect -630 3745 -610 3765
rect -590 3745 -570 3765
rect -550 3745 -530 3765
rect -510 3745 -490 3765
rect -470 3745 -450 3765
rect -430 3745 -410 3765
rect -390 3745 -370 3765
rect -350 3745 -330 3765
rect -310 3745 -290 3765
rect -270 3745 -250 3765
rect -230 3745 -210 3765
rect -190 3745 -170 3765
rect -150 3745 -130 3765
rect -110 3745 -90 3765
rect -70 3745 -50 3765
rect -30 3745 -10 3765
rect 10 3745 30 3765
rect 50 3745 70 3765
rect 90 3745 110 3765
rect 130 3745 150 3765
rect 170 3745 190 3765
rect 210 3745 230 3765
rect 250 3745 270 3765
rect 290 3745 310 3765
rect 330 3745 350 3765
rect 370 3745 390 3765
rect 410 3745 440 3765
rect -5580 3650 -5550 3670
rect -5530 3650 -5510 3670
rect -5490 3650 -5470 3670
rect -5450 3650 -5430 3670
rect -5410 3650 -5390 3670
rect -5370 3650 -5350 3670
rect -5330 3650 -5310 3670
rect -5290 3650 -5270 3670
rect -5250 3650 -5230 3670
rect -5210 3650 -5190 3670
rect -5170 3650 -5150 3670
rect -5130 3650 -5110 3670
rect -5090 3650 -5070 3670
rect -5050 3650 -5030 3670
rect -5010 3650 -4990 3670
rect -4970 3650 -4950 3670
rect -4930 3650 -4910 3670
rect -4890 3650 -4870 3670
rect -4850 3650 -4830 3670
rect -4810 3650 -4790 3670
rect -4770 3650 -4750 3670
rect -4730 3650 -4710 3670
rect -4690 3650 -4670 3670
rect -4650 3650 -4630 3670
rect -4610 3650 -4590 3670
rect -4570 3650 -4550 3670
rect -4530 3650 -4510 3670
rect -4490 3650 -4470 3670
rect -4450 3650 -4430 3670
rect -4410 3650 -4390 3670
rect -4370 3650 -4350 3670
rect -4330 3650 -4310 3670
rect -4290 3650 -4270 3670
rect -4250 3650 -4230 3670
rect -4210 3650 -4190 3670
rect -4170 3650 -4150 3670
rect -4130 3650 -4110 3670
rect -4090 3650 -4070 3670
rect -4050 3650 -4030 3670
rect -4010 3650 -3990 3670
rect -3970 3650 -3950 3670
rect -3930 3650 -3910 3670
rect -3890 3650 -3870 3670
rect -3850 3650 -3830 3670
rect -3810 3650 -3790 3670
rect -3770 3650 -3750 3670
rect -3730 3650 -3710 3670
rect -3690 3650 -3670 3670
rect -3650 3650 -3630 3670
rect -3610 3650 -3590 3670
rect -3570 3650 -3550 3670
rect -3530 3650 -3510 3670
rect -3490 3650 -3470 3670
rect -3450 3650 -3430 3670
rect -3410 3650 -3390 3670
rect -3370 3650 -3350 3670
rect -3330 3650 -3310 3670
rect -3290 3650 -3270 3670
rect -3250 3650 -3230 3670
rect -3210 3650 -3190 3670
rect -3170 3650 -3150 3670
rect -3130 3650 -3110 3670
rect -2030 3650 -2010 3670
rect -1990 3650 -1970 3670
rect -1950 3650 -1930 3670
rect -1910 3650 -1890 3670
rect -1870 3650 -1850 3670
rect -1830 3650 -1810 3670
rect -1790 3650 -1770 3670
rect -1750 3650 -1730 3670
rect -1710 3650 -1690 3670
rect -1670 3650 -1650 3670
rect -1630 3650 -1610 3670
rect -1590 3650 -1570 3670
rect -1550 3650 -1530 3670
rect -1510 3650 -1490 3670
rect -1470 3650 -1450 3670
rect -1430 3650 -1410 3670
rect -1390 3650 -1370 3670
rect -1350 3650 -1330 3670
rect -1310 3650 -1290 3670
rect -1270 3650 -1250 3670
rect -1230 3650 -1210 3670
rect -1190 3650 -1170 3670
rect -1150 3650 -1130 3670
rect -1110 3650 -1090 3670
rect -1070 3650 -1050 3670
rect -1030 3650 -1010 3670
rect -990 3650 -970 3670
rect -950 3650 -930 3670
rect -910 3650 -890 3670
rect -870 3650 -850 3670
rect -830 3650 -810 3670
rect -790 3650 -770 3670
rect -750 3650 -730 3670
rect -710 3650 -690 3670
rect -670 3650 -650 3670
rect -630 3650 -610 3670
rect -590 3650 -570 3670
rect -550 3650 -530 3670
rect -510 3650 -490 3670
rect -470 3650 -450 3670
rect -430 3650 -410 3670
rect -390 3650 -370 3670
rect -350 3650 -330 3670
rect -310 3650 -290 3670
rect -270 3650 -250 3670
rect -230 3650 -210 3670
rect -190 3650 -170 3670
rect -150 3650 -130 3670
rect -110 3650 -90 3670
rect -70 3650 -50 3670
rect -30 3650 -10 3670
rect 10 3650 30 3670
rect 50 3650 70 3670
rect 90 3650 110 3670
rect 130 3650 150 3670
rect 170 3650 190 3670
rect 210 3650 230 3670
rect 250 3650 270 3670
rect 290 3650 310 3670
rect 330 3650 350 3670
rect 370 3650 390 3670
rect 410 3650 440 3670
rect -5580 3555 -5550 3575
rect -5530 3555 -5510 3575
rect -5490 3555 -5470 3575
rect -5450 3555 -5430 3575
rect -5410 3555 -5390 3575
rect -5370 3555 -5350 3575
rect -5330 3555 -5310 3575
rect -5290 3555 -5270 3575
rect -5250 3555 -5230 3575
rect -5210 3555 -5190 3575
rect -5170 3555 -5150 3575
rect -5130 3555 -5110 3575
rect -5090 3555 -5070 3575
rect -5050 3555 -5030 3575
rect -5010 3555 -4990 3575
rect -4970 3555 -4950 3575
rect -4930 3555 -4910 3575
rect -4890 3555 -4870 3575
rect -4850 3555 -4830 3575
rect -4810 3555 -4790 3575
rect -4770 3555 -4750 3575
rect -4730 3555 -4710 3575
rect -4690 3555 -4670 3575
rect -4650 3555 -4630 3575
rect -4610 3555 -4590 3575
rect -4570 3555 -4550 3575
rect -4530 3555 -4510 3575
rect -4490 3555 -4470 3575
rect -4450 3555 -4430 3575
rect -4410 3555 -4390 3575
rect -4370 3555 -4350 3575
rect -4330 3555 -4310 3575
rect -4290 3555 -4270 3575
rect -4250 3555 -4230 3575
rect -4210 3555 -4190 3575
rect -4170 3555 -4150 3575
rect -4130 3555 -4110 3575
rect -4090 3555 -4070 3575
rect -4050 3555 -4030 3575
rect -4010 3555 -3990 3575
rect -3970 3555 -3950 3575
rect -3930 3555 -3910 3575
rect -3890 3555 -3870 3575
rect -3850 3555 -3830 3575
rect -3810 3555 -3790 3575
rect -3770 3555 -3750 3575
rect -3730 3555 -3710 3575
rect -3690 3555 -3670 3575
rect -3650 3555 -3630 3575
rect -3610 3555 -3590 3575
rect -3570 3555 -3550 3575
rect -3530 3555 -3510 3575
rect -3490 3555 -3470 3575
rect -3450 3555 -3430 3575
rect -3410 3555 -3390 3575
rect -3370 3555 -3350 3575
rect -3330 3555 -3310 3575
rect -3290 3555 -3270 3575
rect -3250 3555 -3230 3575
rect -3210 3555 -3190 3575
rect -3170 3555 -3150 3575
rect -3130 3555 -3110 3575
rect -2030 3555 -2010 3575
rect -1990 3555 -1970 3575
rect -1950 3555 -1930 3575
rect -1910 3555 -1890 3575
rect -1870 3555 -1850 3575
rect -1830 3555 -1810 3575
rect -1790 3555 -1770 3575
rect -1750 3555 -1730 3575
rect -1710 3555 -1690 3575
rect -1670 3555 -1650 3575
rect -1630 3555 -1610 3575
rect -1590 3555 -1570 3575
rect -1550 3555 -1530 3575
rect -1510 3555 -1490 3575
rect -1470 3555 -1450 3575
rect -1430 3555 -1410 3575
rect -1390 3555 -1370 3575
rect -1350 3555 -1330 3575
rect -1310 3555 -1290 3575
rect -1270 3555 -1250 3575
rect -1230 3555 -1210 3575
rect -1190 3555 -1170 3575
rect -1150 3555 -1130 3575
rect -1110 3555 -1090 3575
rect -1070 3555 -1050 3575
rect -1030 3555 -1010 3575
rect -990 3555 -970 3575
rect -950 3555 -930 3575
rect -910 3555 -890 3575
rect -870 3555 -850 3575
rect -830 3555 -810 3575
rect -790 3555 -770 3575
rect -750 3555 -730 3575
rect -710 3555 -690 3575
rect -670 3555 -650 3575
rect -630 3555 -610 3575
rect -590 3555 -570 3575
rect -550 3555 -530 3575
rect -510 3555 -490 3575
rect -470 3555 -450 3575
rect -430 3555 -410 3575
rect -390 3555 -370 3575
rect -350 3555 -330 3575
rect -310 3555 -290 3575
rect -270 3555 -250 3575
rect -230 3555 -210 3575
rect -190 3555 -170 3575
rect -150 3555 -130 3575
rect -110 3555 -90 3575
rect -70 3555 -50 3575
rect -30 3555 -10 3575
rect 10 3555 30 3575
rect 50 3555 70 3575
rect 90 3555 110 3575
rect 130 3555 150 3575
rect 170 3555 190 3575
rect 210 3555 230 3575
rect 250 3555 270 3575
rect 290 3555 310 3575
rect 330 3555 350 3575
rect 370 3555 390 3575
rect 410 3555 440 3575
<< psubdiff >>
rect -5665 8520 -3165 8530
rect -5665 8500 -5650 8520
rect -5630 8500 -5610 8520
rect -5590 8500 -5570 8520
rect -5550 8500 -5530 8520
rect -5510 8500 -5490 8520
rect -5470 8500 -5450 8520
rect -5430 8500 -5410 8520
rect -5390 8500 -5370 8520
rect -5350 8500 -5330 8520
rect -5310 8500 -5290 8520
rect -5270 8500 -5250 8520
rect -5230 8500 -5210 8520
rect -5190 8500 -5170 8520
rect -5150 8500 -5130 8520
rect -5110 8500 -5090 8520
rect -5070 8500 -5050 8520
rect -5030 8500 -5010 8520
rect -4990 8500 -4970 8520
rect -4950 8500 -4930 8520
rect -4910 8500 -4890 8520
rect -4870 8500 -4850 8520
rect -4830 8500 -4810 8520
rect -4790 8500 -4770 8520
rect -4750 8500 -4730 8520
rect -4710 8500 -4690 8520
rect -4670 8500 -4650 8520
rect -4630 8500 -4610 8520
rect -4590 8500 -4570 8520
rect -4550 8500 -4530 8520
rect -4510 8500 -4490 8520
rect -4470 8500 -4450 8520
rect -4430 8500 -4410 8520
rect -4390 8500 -4370 8520
rect -4350 8500 -4330 8520
rect -4310 8500 -4290 8520
rect -4270 8500 -4250 8520
rect -4230 8500 -4210 8520
rect -4190 8500 -4170 8520
rect -4150 8500 -4130 8520
rect -4110 8500 -4090 8520
rect -4070 8500 -4050 8520
rect -4030 8500 -4010 8520
rect -3990 8500 -3970 8520
rect -3950 8500 -3930 8520
rect -3910 8500 -3890 8520
rect -3870 8500 -3850 8520
rect -3830 8500 -3810 8520
rect -3790 8500 -3770 8520
rect -3750 8500 -3730 8520
rect -3710 8500 -3690 8520
rect -3670 8500 -3650 8520
rect -3630 8500 -3610 8520
rect -3590 8500 -3570 8520
rect -3550 8500 -3530 8520
rect -3510 8500 -3490 8520
rect -3470 8500 -3450 8520
rect -3430 8500 -3410 8520
rect -3390 8500 -3370 8520
rect -3350 8500 -3330 8520
rect -3310 8500 -3290 8520
rect -3270 8500 -3250 8520
rect -3230 8500 -3210 8520
rect -3190 8500 -3165 8520
rect -5665 8490 -3165 8500
rect -5665 6305 -3165 6315
rect -5665 6285 -5650 6305
rect -5630 6285 -5610 6305
rect -5590 6285 -5570 6305
rect -5550 6285 -5530 6305
rect -5510 6285 -5490 6305
rect -5470 6285 -5450 6305
rect -5430 6285 -5410 6305
rect -5390 6285 -5370 6305
rect -5350 6285 -5330 6305
rect -5310 6285 -5290 6305
rect -5270 6285 -5250 6305
rect -5230 6285 -5210 6305
rect -5190 6285 -5170 6305
rect -5150 6285 -5130 6305
rect -5110 6285 -5090 6305
rect -5070 6285 -5050 6305
rect -5030 6285 -5010 6305
rect -4990 6285 -4970 6305
rect -4950 6285 -4930 6305
rect -4910 6285 -4890 6305
rect -4870 6285 -4850 6305
rect -4830 6285 -4810 6305
rect -4790 6285 -4770 6305
rect -4750 6285 -4730 6305
rect -4710 6285 -4690 6305
rect -4670 6285 -4650 6305
rect -4630 6285 -4610 6305
rect -4590 6285 -4570 6305
rect -4550 6285 -4530 6305
rect -4510 6285 -4490 6305
rect -4470 6285 -4450 6305
rect -4430 6285 -4410 6305
rect -4390 6285 -4370 6305
rect -4350 6285 -4330 6305
rect -4310 6285 -4290 6305
rect -4270 6285 -4250 6305
rect -4230 6285 -4210 6305
rect -4190 6285 -4170 6305
rect -4150 6285 -4130 6305
rect -4110 6285 -4090 6305
rect -4070 6285 -4050 6305
rect -4030 6285 -4010 6305
rect -3990 6285 -3970 6305
rect -3950 6285 -3930 6305
rect -3910 6285 -3890 6305
rect -3870 6285 -3850 6305
rect -3830 6285 -3810 6305
rect -3790 6285 -3770 6305
rect -3750 6285 -3730 6305
rect -3710 6285 -3690 6305
rect -3670 6285 -3650 6305
rect -3630 6285 -3610 6305
rect -3590 6285 -3570 6305
rect -3550 6285 -3530 6305
rect -3510 6285 -3490 6305
rect -3470 6285 -3450 6305
rect -3430 6285 -3410 6305
rect -3390 6285 -3370 6305
rect -3350 6285 -3330 6305
rect -3310 6285 -3290 6305
rect -3270 6285 -3250 6305
rect -3230 6285 -3210 6305
rect -3190 6285 -3165 6305
rect -5665 6275 -3165 6285
rect -1975 8520 525 8530
rect -1975 8500 -1950 8520
rect -1930 8500 -1910 8520
rect -1890 8500 -1870 8520
rect -1850 8500 -1830 8520
rect -1810 8500 -1790 8520
rect -1770 8500 -1750 8520
rect -1730 8500 -1710 8520
rect -1690 8500 -1670 8520
rect -1650 8500 -1630 8520
rect -1610 8500 -1590 8520
rect -1570 8500 -1550 8520
rect -1530 8500 -1510 8520
rect -1490 8500 -1470 8520
rect -1450 8500 -1430 8520
rect -1410 8500 -1390 8520
rect -1370 8500 -1350 8520
rect -1330 8500 -1310 8520
rect -1290 8500 -1270 8520
rect -1250 8500 -1230 8520
rect -1210 8500 -1190 8520
rect -1170 8500 -1150 8520
rect -1130 8500 -1110 8520
rect -1090 8500 -1070 8520
rect -1050 8500 -1030 8520
rect -1010 8500 -990 8520
rect -970 8500 -950 8520
rect -930 8500 -910 8520
rect -890 8500 -870 8520
rect -850 8500 -830 8520
rect -810 8500 -790 8520
rect -770 8500 -750 8520
rect -730 8500 -710 8520
rect -690 8500 -670 8520
rect -650 8500 -630 8520
rect -610 8500 -590 8520
rect -570 8500 -550 8520
rect -530 8500 -510 8520
rect -490 8500 -470 8520
rect -450 8500 -430 8520
rect -410 8500 -390 8520
rect -370 8500 -350 8520
rect -330 8500 -310 8520
rect -290 8500 -270 8520
rect -250 8500 -230 8520
rect -210 8500 -190 8520
rect -170 8500 -150 8520
rect -130 8500 -110 8520
rect -90 8500 -70 8520
rect -50 8500 -30 8520
rect -10 8500 10 8520
rect 30 8500 50 8520
rect 70 8500 90 8520
rect 110 8500 130 8520
rect 150 8500 170 8520
rect 190 8500 210 8520
rect 230 8500 250 8520
rect 270 8500 290 8520
rect 310 8500 330 8520
rect 350 8500 370 8520
rect 390 8500 410 8520
rect 430 8500 450 8520
rect 470 8500 490 8520
rect 510 8500 525 8520
rect -1975 8490 525 8500
rect -1975 6305 525 6315
rect -1975 6285 -1950 6305
rect -1930 6285 -1910 6305
rect -1890 6285 -1870 6305
rect -1850 6285 -1830 6305
rect -1810 6285 -1790 6305
rect -1770 6285 -1750 6305
rect -1730 6285 -1710 6305
rect -1690 6285 -1670 6305
rect -1650 6285 -1630 6305
rect -1610 6285 -1590 6305
rect -1570 6285 -1550 6305
rect -1530 6285 -1510 6305
rect -1490 6285 -1470 6305
rect -1450 6285 -1430 6305
rect -1410 6285 -1390 6305
rect -1370 6285 -1350 6305
rect -1330 6285 -1310 6305
rect -1290 6285 -1270 6305
rect -1250 6285 -1230 6305
rect -1210 6285 -1190 6305
rect -1170 6285 -1150 6305
rect -1130 6285 -1110 6305
rect -1090 6285 -1070 6305
rect -1050 6285 -1030 6305
rect -1010 6285 -990 6305
rect -970 6285 -950 6305
rect -930 6285 -910 6305
rect -890 6285 -870 6305
rect -850 6285 -830 6305
rect -810 6285 -790 6305
rect -770 6285 -750 6305
rect -730 6285 -710 6305
rect -690 6285 -670 6305
rect -650 6285 -630 6305
rect -610 6285 -590 6305
rect -570 6285 -550 6305
rect -530 6285 -510 6305
rect -490 6285 -470 6305
rect -450 6285 -430 6305
rect -410 6285 -390 6305
rect -370 6285 -350 6305
rect -330 6285 -310 6305
rect -290 6285 -270 6305
rect -250 6285 -230 6305
rect -210 6285 -190 6305
rect -170 6285 -150 6305
rect -130 6285 -110 6305
rect -90 6285 -70 6305
rect -50 6285 -30 6305
rect -10 6285 10 6305
rect 30 6285 50 6305
rect 70 6285 90 6305
rect 110 6285 130 6305
rect 150 6285 170 6305
rect 190 6285 210 6305
rect 230 6285 250 6305
rect 270 6285 290 6305
rect 310 6285 330 6305
rect 350 6285 370 6305
rect 390 6285 410 6305
rect 430 6285 450 6305
rect 470 6285 490 6305
rect 510 6285 525 6305
rect -1975 6275 525 6285
rect -5595 6085 -3095 6095
rect -5595 6065 -5580 6085
rect -5550 6065 -5530 6085
rect -5510 6065 -5490 6085
rect -5470 6065 -5450 6085
rect -5430 6065 -5410 6085
rect -5390 6065 -5370 6085
rect -5350 6065 -5330 6085
rect -5310 6065 -5290 6085
rect -5270 6065 -5250 6085
rect -5230 6065 -5210 6085
rect -5190 6065 -5170 6085
rect -5150 6065 -5130 6085
rect -5110 6065 -5090 6085
rect -5070 6065 -5050 6085
rect -5030 6065 -5010 6085
rect -4990 6065 -4970 6085
rect -4950 6065 -4930 6085
rect -4910 6065 -4890 6085
rect -4870 6065 -4850 6085
rect -4830 6065 -4810 6085
rect -4790 6065 -4770 6085
rect -4750 6065 -4730 6085
rect -4710 6065 -4690 6085
rect -4670 6065 -4650 6085
rect -4630 6065 -4610 6085
rect -4590 6065 -4570 6085
rect -4550 6065 -4530 6085
rect -4510 6065 -4490 6085
rect -4470 6065 -4450 6085
rect -4430 6065 -4410 6085
rect -4390 6065 -4370 6085
rect -4350 6065 -4330 6085
rect -4310 6065 -4290 6085
rect -4270 6065 -4250 6085
rect -4230 6065 -4210 6085
rect -4190 6065 -4170 6085
rect -4150 6065 -4130 6085
rect -4110 6065 -4090 6085
rect -4070 6065 -4050 6085
rect -4030 6065 -4010 6085
rect -3990 6065 -3970 6085
rect -3950 6065 -3930 6085
rect -3910 6065 -3890 6085
rect -3870 6065 -3850 6085
rect -3830 6065 -3810 6085
rect -3790 6065 -3770 6085
rect -3750 6065 -3730 6085
rect -3710 6065 -3690 6085
rect -3670 6065 -3650 6085
rect -3630 6065 -3610 6085
rect -3590 6065 -3570 6085
rect -3550 6065 -3530 6085
rect -3510 6065 -3490 6085
rect -3470 6065 -3450 6085
rect -3430 6065 -3410 6085
rect -3390 6065 -3370 6085
rect -3350 6065 -3330 6085
rect -3310 6065 -3290 6085
rect -3270 6065 -3250 6085
rect -3230 6065 -3210 6085
rect -3190 6065 -3170 6085
rect -3150 6065 -3130 6085
rect -3110 6065 -3095 6085
rect -5595 6055 -3095 6065
rect -2045 6085 455 6095
rect -2045 6065 -2030 6085
rect -2010 6065 -1990 6085
rect -1970 6065 -1950 6085
rect -1930 6065 -1910 6085
rect -1890 6065 -1870 6085
rect -1850 6065 -1830 6085
rect -1810 6065 -1790 6085
rect -1770 6065 -1750 6085
rect -1730 6065 -1710 6085
rect -1690 6065 -1670 6085
rect -1650 6065 -1630 6085
rect -1610 6065 -1590 6085
rect -1570 6065 -1550 6085
rect -1530 6065 -1510 6085
rect -1490 6065 -1470 6085
rect -1450 6065 -1430 6085
rect -1410 6065 -1390 6085
rect -1370 6065 -1350 6085
rect -1330 6065 -1310 6085
rect -1290 6065 -1270 6085
rect -1250 6065 -1230 6085
rect -1210 6065 -1190 6085
rect -1170 6065 -1150 6085
rect -1130 6065 -1110 6085
rect -1090 6065 -1070 6085
rect -1050 6065 -1030 6085
rect -1010 6065 -990 6085
rect -970 6065 -950 6085
rect -930 6065 -910 6085
rect -890 6065 -870 6085
rect -850 6065 -830 6085
rect -810 6065 -790 6085
rect -770 6065 -750 6085
rect -730 6065 -710 6085
rect -690 6065 -670 6085
rect -650 6065 -630 6085
rect -610 6065 -590 6085
rect -570 6065 -550 6085
rect -530 6065 -510 6085
rect -490 6065 -470 6085
rect -450 6065 -430 6085
rect -410 6065 -390 6085
rect -370 6065 -350 6085
rect -330 6065 -310 6085
rect -290 6065 -270 6085
rect -250 6065 -230 6085
rect -210 6065 -190 6085
rect -170 6065 -150 6085
rect -130 6065 -110 6085
rect -90 6065 -70 6085
rect -50 6065 -30 6085
rect -10 6065 10 6085
rect 30 6065 50 6085
rect 70 6065 90 6085
rect 110 6065 130 6085
rect 150 6065 170 6085
rect 190 6065 210 6085
rect 230 6065 250 6085
rect 270 6065 290 6085
rect 310 6065 330 6085
rect 350 6065 370 6085
rect 390 6065 410 6085
rect 440 6065 455 6085
rect -2045 6055 455 6065
rect -5595 3535 -3095 3545
rect -5595 3515 -5580 3535
rect -5550 3515 -5530 3535
rect -5510 3515 -5490 3535
rect -5470 3515 -5450 3535
rect -5430 3515 -5410 3535
rect -5390 3515 -5370 3535
rect -5350 3515 -5330 3535
rect -5310 3515 -5290 3535
rect -5270 3515 -5250 3535
rect -5230 3515 -5210 3535
rect -5190 3515 -5170 3535
rect -5150 3515 -5130 3535
rect -5110 3515 -5090 3535
rect -5070 3515 -5050 3535
rect -5030 3515 -5010 3535
rect -4990 3515 -4970 3535
rect -4950 3515 -4930 3535
rect -4910 3515 -4890 3535
rect -4870 3515 -4850 3535
rect -4830 3515 -4810 3535
rect -4790 3515 -4770 3535
rect -4750 3515 -4730 3535
rect -4710 3515 -4690 3535
rect -4670 3515 -4650 3535
rect -4630 3515 -4610 3535
rect -4590 3515 -4570 3535
rect -4550 3515 -4530 3535
rect -4510 3515 -4490 3535
rect -4470 3515 -4450 3535
rect -4430 3515 -4410 3535
rect -4390 3515 -4370 3535
rect -4350 3515 -4330 3535
rect -4310 3515 -4290 3535
rect -4270 3515 -4250 3535
rect -4230 3515 -4210 3535
rect -4190 3515 -4170 3535
rect -4150 3515 -4130 3535
rect -4110 3515 -4090 3535
rect -4070 3515 -4050 3535
rect -4030 3515 -4010 3535
rect -3990 3515 -3970 3535
rect -3950 3515 -3930 3535
rect -3910 3515 -3890 3535
rect -3870 3515 -3850 3535
rect -3830 3515 -3810 3535
rect -3790 3515 -3770 3535
rect -3750 3515 -3730 3535
rect -3710 3515 -3690 3535
rect -3670 3515 -3650 3535
rect -3630 3515 -3610 3535
rect -3590 3515 -3570 3535
rect -3550 3515 -3530 3535
rect -3510 3515 -3490 3535
rect -3470 3515 -3450 3535
rect -3430 3515 -3410 3535
rect -3390 3515 -3370 3535
rect -3350 3515 -3330 3535
rect -3310 3515 -3290 3535
rect -3270 3515 -3250 3535
rect -3230 3515 -3210 3535
rect -3190 3515 -3170 3535
rect -3150 3515 -3130 3535
rect -3110 3515 -3095 3535
rect -5595 3505 -3095 3515
rect -2045 3535 455 3545
rect -2045 3515 -2030 3535
rect -2010 3515 -1990 3535
rect -1970 3515 -1950 3535
rect -1930 3515 -1910 3535
rect -1890 3515 -1870 3535
rect -1850 3515 -1830 3535
rect -1810 3515 -1790 3535
rect -1770 3515 -1750 3535
rect -1730 3515 -1710 3535
rect -1690 3515 -1670 3535
rect -1650 3515 -1630 3535
rect -1610 3515 -1590 3535
rect -1570 3515 -1550 3535
rect -1530 3515 -1510 3535
rect -1490 3515 -1470 3535
rect -1450 3515 -1430 3535
rect -1410 3515 -1390 3535
rect -1370 3515 -1350 3535
rect -1330 3515 -1310 3535
rect -1290 3515 -1270 3535
rect -1250 3515 -1230 3535
rect -1210 3515 -1190 3535
rect -1170 3515 -1150 3535
rect -1130 3515 -1110 3535
rect -1090 3515 -1070 3535
rect -1050 3515 -1030 3535
rect -1010 3515 -990 3535
rect -970 3515 -950 3535
rect -930 3515 -910 3535
rect -890 3515 -870 3535
rect -850 3515 -830 3535
rect -810 3515 -790 3535
rect -770 3515 -750 3535
rect -730 3515 -710 3535
rect -690 3515 -670 3535
rect -650 3515 -630 3535
rect -610 3515 -590 3535
rect -570 3515 -550 3535
rect -530 3515 -510 3535
rect -490 3515 -470 3535
rect -450 3515 -430 3535
rect -410 3515 -390 3535
rect -370 3515 -350 3535
rect -330 3515 -310 3535
rect -290 3515 -270 3535
rect -250 3515 -230 3535
rect -210 3515 -190 3535
rect -170 3515 -150 3535
rect -130 3515 -110 3535
rect -90 3515 -70 3535
rect -50 3515 -30 3535
rect -10 3515 10 3535
rect 30 3515 50 3535
rect 70 3515 90 3535
rect 110 3515 130 3535
rect 150 3515 170 3535
rect 190 3515 210 3535
rect 230 3515 250 3535
rect 270 3515 290 3535
rect 310 3515 330 3535
rect 350 3515 370 3535
rect 390 3515 410 3535
rect 440 3515 455 3535
rect -2045 3505 455 3515
<< nsubdiff >>
rect -5775 8605 -2915 8620
rect -5775 8585 -5710 8605
rect -5690 8585 -5670 8605
rect -5650 8585 -5630 8605
rect -5610 8585 -5590 8605
rect -5570 8585 -5550 8605
rect -5530 8585 -5510 8605
rect -5490 8585 -5470 8605
rect -5450 8585 -5430 8605
rect -5410 8585 -5390 8605
rect -5370 8585 -5350 8605
rect -5330 8585 -5310 8605
rect -5290 8585 -5270 8605
rect -5250 8585 -5230 8605
rect -5210 8585 -5190 8605
rect -5170 8585 -5150 8605
rect -5130 8585 -5110 8605
rect -5090 8585 -5070 8605
rect -5050 8585 -5030 8605
rect -5010 8585 -4990 8605
rect -4970 8585 -4950 8605
rect -4930 8585 -4910 8605
rect -4890 8585 -4870 8605
rect -4850 8585 -4830 8605
rect -4810 8585 -4790 8605
rect -4770 8585 -4750 8605
rect -4730 8585 -4710 8605
rect -4690 8585 -4670 8605
rect -4650 8585 -4630 8605
rect -4610 8585 -4590 8605
rect -4570 8585 -4550 8605
rect -4530 8585 -4510 8605
rect -4490 8585 -4470 8605
rect -4450 8585 -4430 8605
rect -4410 8585 -4390 8605
rect -4370 8585 -4350 8605
rect -4330 8585 -4310 8605
rect -4290 8585 -4270 8605
rect -4250 8585 -4230 8605
rect -4210 8585 -4190 8605
rect -4170 8585 -4150 8605
rect -4130 8585 -4110 8605
rect -4090 8585 -4070 8605
rect -4050 8585 -4030 8605
rect -4010 8585 -3990 8605
rect -3970 8585 -3950 8605
rect -3930 8585 -3910 8605
rect -3890 8585 -3870 8605
rect -3850 8585 -3830 8605
rect -3810 8585 -3790 8605
rect -3770 8585 -3750 8605
rect -3730 8585 -3710 8605
rect -3690 8585 -3670 8605
rect -3650 8585 -3630 8605
rect -3610 8585 -3590 8605
rect -3570 8585 -3550 8605
rect -3530 8585 -3510 8605
rect -3490 8585 -3470 8605
rect -3450 8585 -3430 8605
rect -3410 8585 -3390 8605
rect -3370 8585 -3350 8605
rect -3330 8585 -3310 8605
rect -3290 8585 -3270 8605
rect -3250 8585 -3230 8605
rect -3210 8585 -3190 8605
rect -3170 8585 -3150 8605
rect -3130 8585 -3110 8605
rect -3090 8585 -3070 8605
rect -3050 8585 -3030 8605
rect -3010 8585 -2990 8605
rect -2970 8585 -2915 8605
rect -5775 8570 -2915 8585
rect -5775 8550 -5760 8570
rect -5740 8550 -5725 8570
rect -5775 8530 -5725 8550
rect -2965 8550 -2950 8570
rect -2930 8550 -2915 8570
rect -2965 8530 -2915 8550
rect -5775 8510 -5760 8530
rect -5740 8510 -5725 8530
rect -5775 8490 -5725 8510
rect -5775 8470 -5760 8490
rect -5740 8470 -5725 8490
rect -5775 8450 -5725 8470
rect -5775 8430 -5760 8450
rect -5740 8430 -5725 8450
rect -2965 8510 -2950 8530
rect -2930 8510 -2915 8530
rect -2965 8490 -2915 8510
rect -2965 8470 -2950 8490
rect -2930 8470 -2915 8490
rect -2965 8450 -2915 8470
rect -5775 8410 -5725 8430
rect -5775 8390 -5760 8410
rect -5740 8390 -5725 8410
rect -5775 8370 -5725 8390
rect -5775 8350 -5760 8370
rect -5740 8350 -5725 8370
rect -2965 8430 -2950 8450
rect -2930 8430 -2915 8450
rect -2965 8410 -2915 8430
rect -2965 8390 -2950 8410
rect -2930 8390 -2915 8410
rect -2965 8370 -2915 8390
rect -5775 8330 -5725 8350
rect -5775 8310 -5760 8330
rect -5740 8310 -5725 8330
rect -5775 8290 -5725 8310
rect -5775 8270 -5760 8290
rect -5740 8270 -5725 8290
rect -2965 8350 -2950 8370
rect -2930 8350 -2915 8370
rect -2965 8330 -2915 8350
rect -2965 8310 -2950 8330
rect -2930 8310 -2915 8330
rect -2965 8290 -2915 8310
rect -5775 8250 -5725 8270
rect -5775 8230 -5760 8250
rect -5740 8230 -5725 8250
rect -5775 8210 -5725 8230
rect -5775 8190 -5760 8210
rect -5740 8190 -5725 8210
rect -2965 8270 -2950 8290
rect -2930 8270 -2915 8290
rect -2965 8250 -2915 8270
rect -2965 8230 -2950 8250
rect -2930 8230 -2915 8250
rect -2965 8210 -2915 8230
rect -5775 8170 -5725 8190
rect -5775 8150 -5760 8170
rect -5740 8150 -5725 8170
rect -5775 8130 -5725 8150
rect -5775 8110 -5760 8130
rect -5740 8110 -5725 8130
rect -2965 8190 -2950 8210
rect -2930 8190 -2915 8210
rect -2965 8170 -2915 8190
rect -2965 8150 -2950 8170
rect -2930 8150 -2915 8170
rect -2965 8130 -2915 8150
rect -5775 8090 -5725 8110
rect -5775 8070 -5760 8090
rect -5740 8070 -5725 8090
rect -5775 8050 -5725 8070
rect -5775 8030 -5760 8050
rect -5740 8030 -5725 8050
rect -2965 8110 -2950 8130
rect -2930 8110 -2915 8130
rect -2965 8090 -2915 8110
rect -2965 8070 -2950 8090
rect -2930 8070 -2915 8090
rect -2965 8050 -2915 8070
rect -5775 8010 -5725 8030
rect -5775 7990 -5760 8010
rect -5740 7990 -5725 8010
rect -5775 7970 -5725 7990
rect -5775 7950 -5760 7970
rect -5740 7950 -5725 7970
rect -2965 8030 -2950 8050
rect -2930 8030 -2915 8050
rect -2965 8010 -2915 8030
rect -2965 7990 -2950 8010
rect -2930 7990 -2915 8010
rect -2965 7970 -2915 7990
rect -5775 7930 -5725 7950
rect -5775 7910 -5760 7930
rect -5740 7910 -5725 7930
rect -5775 7890 -5725 7910
rect -5775 7870 -5760 7890
rect -5740 7870 -5725 7890
rect -5775 7850 -5725 7870
rect -2965 7950 -2950 7970
rect -2930 7950 -2915 7970
rect -2965 7930 -2915 7950
rect -2965 7910 -2950 7930
rect -2930 7910 -2915 7930
rect -2965 7890 -2915 7910
rect -2965 7870 -2950 7890
rect -2930 7870 -2915 7890
rect -5775 7830 -5760 7850
rect -5740 7830 -5725 7850
rect -5775 7810 -5725 7830
rect -5775 7790 -5760 7810
rect -5740 7790 -5725 7810
rect -5775 7770 -5725 7790
rect -2965 7850 -2915 7870
rect -2965 7830 -2950 7850
rect -2930 7830 -2915 7850
rect -2965 7810 -2915 7830
rect -2965 7790 -2950 7810
rect -2930 7790 -2915 7810
rect -5775 7750 -5760 7770
rect -5740 7750 -5725 7770
rect -5775 7730 -5725 7750
rect -5775 7710 -5760 7730
rect -5740 7710 -5725 7730
rect -5775 7690 -5725 7710
rect -2965 7770 -2915 7790
rect -2965 7750 -2950 7770
rect -2930 7750 -2915 7770
rect -2965 7730 -2915 7750
rect -2965 7710 -2950 7730
rect -2930 7710 -2915 7730
rect -5775 7670 -5760 7690
rect -5740 7670 -5725 7690
rect -5775 7650 -5725 7670
rect -5775 7630 -5760 7650
rect -5740 7630 -5725 7650
rect -5775 7610 -5725 7630
rect -2965 7690 -2915 7710
rect -2965 7670 -2950 7690
rect -2930 7670 -2915 7690
rect -2965 7650 -2915 7670
rect -2965 7630 -2950 7650
rect -2930 7630 -2915 7650
rect -5775 7590 -5760 7610
rect -5740 7590 -5725 7610
rect -5775 7570 -5725 7590
rect -5775 7550 -5760 7570
rect -5740 7550 -5725 7570
rect -5775 7530 -5725 7550
rect -2965 7610 -2915 7630
rect -2965 7590 -2950 7610
rect -2930 7590 -2915 7610
rect -2965 7570 -2915 7590
rect -2965 7550 -2950 7570
rect -2930 7550 -2915 7570
rect -5775 7510 -5760 7530
rect -5740 7510 -5725 7530
rect -5775 7490 -5725 7510
rect -5775 7470 -5760 7490
rect -5740 7470 -5725 7490
rect -5775 7450 -5725 7470
rect -2965 7530 -2915 7550
rect -2965 7510 -2950 7530
rect -2930 7510 -2915 7530
rect -2965 7490 -2915 7510
rect -2965 7470 -2950 7490
rect -2930 7470 -2915 7490
rect -5775 7430 -5760 7450
rect -5740 7430 -5725 7450
rect -5775 7410 -5725 7430
rect -5775 7390 -5760 7410
rect -5740 7390 -5725 7410
rect -5775 7370 -5725 7390
rect -2965 7450 -2915 7470
rect -2965 7430 -2950 7450
rect -2930 7430 -2915 7450
rect -2965 7410 -2915 7430
rect -2965 7390 -2950 7410
rect -2930 7390 -2915 7410
rect -5775 7350 -5760 7370
rect -5740 7350 -5725 7370
rect -5775 7330 -5725 7350
rect -5775 7310 -5760 7330
rect -5740 7310 -5725 7330
rect -5775 7290 -5725 7310
rect -2965 7370 -2915 7390
rect -2965 7350 -2950 7370
rect -2930 7350 -2915 7370
rect -2965 7330 -2915 7350
rect -2965 7310 -2950 7330
rect -2930 7310 -2915 7330
rect -5775 7270 -5760 7290
rect -5740 7270 -5725 7290
rect -5775 7250 -5725 7270
rect -5775 7230 -5760 7250
rect -5740 7230 -5725 7250
rect -5775 7210 -5725 7230
rect -2965 7290 -2915 7310
rect -2965 7270 -2950 7290
rect -2930 7270 -2915 7290
rect -2965 7250 -2915 7270
rect -2965 7230 -2950 7250
rect -2930 7230 -2915 7250
rect -5775 7190 -5760 7210
rect -5740 7190 -5725 7210
rect -5775 7170 -5725 7190
rect -5775 7150 -5760 7170
rect -5740 7150 -5725 7170
rect -5775 7130 -5725 7150
rect -2965 7210 -2915 7230
rect -2965 7190 -2950 7210
rect -2930 7190 -2915 7210
rect -2965 7170 -2915 7190
rect -2965 7150 -2950 7170
rect -2930 7150 -2915 7170
rect -5775 7110 -5760 7130
rect -5740 7110 -5725 7130
rect -5775 7090 -5725 7110
rect -5775 7070 -5760 7090
rect -5740 7070 -5725 7090
rect -5775 7050 -5725 7070
rect -5775 7030 -5760 7050
rect -5740 7030 -5725 7050
rect -2965 7130 -2915 7150
rect -2965 7110 -2950 7130
rect -2930 7110 -2915 7130
rect -2965 7090 -2915 7110
rect -2965 7070 -2950 7090
rect -2930 7070 -2915 7090
rect -2965 7050 -2915 7070
rect -5775 7010 -5725 7030
rect -5775 6990 -5760 7010
rect -5740 6990 -5725 7010
rect -5775 6970 -5725 6990
rect -5775 6950 -5760 6970
rect -5740 6950 -5725 6970
rect -2965 7030 -2950 7050
rect -2930 7030 -2915 7050
rect -2965 7010 -2915 7030
rect -2965 6990 -2950 7010
rect -2930 6990 -2915 7010
rect -2965 6970 -2915 6990
rect -5775 6930 -5725 6950
rect -5775 6910 -5760 6930
rect -5740 6910 -5725 6930
rect -5775 6890 -5725 6910
rect -5775 6870 -5760 6890
rect -5740 6870 -5725 6890
rect -2965 6950 -2950 6970
rect -2930 6950 -2915 6970
rect -2965 6930 -2915 6950
rect -2965 6910 -2950 6930
rect -2930 6910 -2915 6930
rect -2965 6890 -2915 6910
rect -5775 6850 -5725 6870
rect -5775 6830 -5760 6850
rect -5740 6830 -5725 6850
rect -5775 6810 -5725 6830
rect -5775 6790 -5760 6810
rect -5740 6790 -5725 6810
rect -2965 6870 -2950 6890
rect -2930 6870 -2915 6890
rect -2965 6850 -2915 6870
rect -2965 6830 -2950 6850
rect -2930 6830 -2915 6850
rect -2965 6810 -2915 6830
rect -5775 6770 -5725 6790
rect -5775 6750 -5760 6770
rect -5740 6750 -5725 6770
rect -5775 6730 -5725 6750
rect -5775 6710 -5760 6730
rect -5740 6710 -5725 6730
rect -2965 6790 -2950 6810
rect -2930 6790 -2915 6810
rect -2965 6770 -2915 6790
rect -2965 6750 -2950 6770
rect -2930 6750 -2915 6770
rect -2965 6730 -2915 6750
rect -5775 6690 -5725 6710
rect -5775 6670 -5760 6690
rect -5740 6670 -5725 6690
rect -5775 6650 -5725 6670
rect -5775 6630 -5760 6650
rect -5740 6630 -5725 6650
rect -2965 6710 -2950 6730
rect -2930 6710 -2915 6730
rect -2965 6690 -2915 6710
rect -2965 6670 -2950 6690
rect -2930 6670 -2915 6690
rect -2965 6650 -2915 6670
rect -5775 6610 -5725 6630
rect -5775 6590 -5760 6610
rect -5740 6590 -5725 6610
rect -5775 6570 -5725 6590
rect -5775 6550 -5760 6570
rect -5740 6550 -5725 6570
rect -2965 6630 -2950 6650
rect -2930 6630 -2915 6650
rect -2965 6610 -2915 6630
rect -2965 6590 -2950 6610
rect -2930 6590 -2915 6610
rect -2965 6570 -2915 6590
rect -5775 6530 -5725 6550
rect -5775 6510 -5760 6530
rect -5740 6510 -5725 6530
rect -5775 6490 -5725 6510
rect -5775 6470 -5760 6490
rect -5740 6470 -5725 6490
rect -2965 6550 -2950 6570
rect -2930 6550 -2915 6570
rect -2965 6530 -2915 6550
rect -2965 6510 -2950 6530
rect -2930 6510 -2915 6530
rect -2965 6490 -2915 6510
rect -5775 6450 -5725 6470
rect -5775 6430 -5760 6450
rect -5740 6430 -5725 6450
rect -5775 6410 -5725 6430
rect -5775 6390 -5760 6410
rect -5740 6390 -5725 6410
rect -2965 6470 -2950 6490
rect -2930 6470 -2915 6490
rect -2965 6450 -2915 6470
rect -2965 6430 -2950 6450
rect -2930 6430 -2915 6450
rect -2965 6410 -2915 6430
rect -5775 6370 -5725 6390
rect -5775 6350 -5760 6370
rect -5740 6350 -5725 6370
rect -2965 6390 -2950 6410
rect -2930 6390 -2915 6410
rect -2965 6370 -2915 6390
rect -5775 6330 -5725 6350
rect -5775 6310 -5760 6330
rect -5740 6310 -5725 6330
rect -5775 6290 -5725 6310
rect -5775 6270 -5760 6290
rect -5740 6270 -5725 6290
rect -2965 6350 -2950 6370
rect -2930 6350 -2915 6370
rect -2965 6330 -2915 6350
rect -2965 6310 -2950 6330
rect -2930 6310 -2915 6330
rect -2965 6290 -2915 6310
rect -5775 6250 -5725 6270
rect -5775 6230 -5760 6250
rect -5740 6235 -5725 6250
rect -2965 6270 -2950 6290
rect -2930 6270 -2915 6290
rect -2965 6250 -2915 6270
rect -2965 6235 -2950 6250
rect -5740 6230 -2950 6235
rect -2930 6230 -2915 6250
rect -5775 6220 -2915 6230
rect -5775 6200 -5710 6220
rect -5690 6200 -5670 6220
rect -5650 6200 -5630 6220
rect -5610 6200 -5590 6220
rect -5570 6200 -5550 6220
rect -5530 6200 -5510 6220
rect -5490 6200 -5470 6220
rect -5450 6200 -5430 6220
rect -5410 6200 -5390 6220
rect -5370 6200 -5350 6220
rect -5330 6200 -5310 6220
rect -5290 6200 -5270 6220
rect -5250 6200 -5230 6220
rect -5210 6200 -5190 6220
rect -5170 6200 -5150 6220
rect -5130 6200 -5110 6220
rect -5090 6200 -5070 6220
rect -5050 6200 -5030 6220
rect -5010 6200 -4990 6220
rect -4970 6200 -4950 6220
rect -4930 6200 -4910 6220
rect -4890 6200 -4870 6220
rect -4850 6200 -4830 6220
rect -4810 6200 -4790 6220
rect -4770 6200 -4750 6220
rect -4730 6200 -4710 6220
rect -4690 6200 -4670 6220
rect -4650 6200 -4630 6220
rect -4610 6200 -4590 6220
rect -4570 6200 -4550 6220
rect -4530 6200 -4510 6220
rect -4490 6200 -4470 6220
rect -4450 6200 -4430 6220
rect -4410 6200 -4390 6220
rect -4370 6200 -4350 6220
rect -4330 6200 -4310 6220
rect -4290 6200 -4270 6220
rect -4250 6200 -4230 6220
rect -4210 6200 -4190 6220
rect -4170 6200 -4150 6220
rect -4130 6200 -4110 6220
rect -4090 6200 -4070 6220
rect -4050 6200 -4030 6220
rect -4010 6200 -3990 6220
rect -3970 6200 -3950 6220
rect -3930 6200 -3910 6220
rect -3890 6200 -3870 6220
rect -3850 6200 -3830 6220
rect -3810 6200 -3790 6220
rect -3770 6200 -3750 6220
rect -3730 6200 -3710 6220
rect -3690 6200 -3670 6220
rect -3650 6200 -3630 6220
rect -3610 6200 -3590 6220
rect -3570 6200 -3550 6220
rect -3530 6200 -3510 6220
rect -3490 6200 -3470 6220
rect -3450 6200 -3430 6220
rect -3410 6200 -3390 6220
rect -3370 6200 -3350 6220
rect -3330 6200 -3310 6220
rect -3290 6200 -3270 6220
rect -3250 6200 -3230 6220
rect -3210 6200 -3190 6220
rect -3170 6200 -3150 6220
rect -3130 6200 -3110 6220
rect -3090 6200 -3070 6220
rect -3050 6200 -3030 6220
rect -3010 6200 -2990 6220
rect -2970 6200 -2915 6220
rect -5775 6185 -2915 6200
rect -2225 8605 635 8620
rect -2225 8585 -2170 8605
rect -2150 8585 -2130 8605
rect -2110 8585 -2090 8605
rect -2070 8585 -2050 8605
rect -2030 8585 -2010 8605
rect -1990 8585 -1970 8605
rect -1950 8585 -1930 8605
rect -1910 8585 -1890 8605
rect -1870 8585 -1850 8605
rect -1830 8585 -1810 8605
rect -1790 8585 -1770 8605
rect -1750 8585 -1730 8605
rect -1710 8585 -1690 8605
rect -1670 8585 -1650 8605
rect -1630 8585 -1610 8605
rect -1590 8585 -1570 8605
rect -1550 8585 -1530 8605
rect -1510 8585 -1490 8605
rect -1470 8585 -1450 8605
rect -1430 8585 -1410 8605
rect -1390 8585 -1370 8605
rect -1350 8585 -1330 8605
rect -1310 8585 -1290 8605
rect -1270 8585 -1250 8605
rect -1230 8585 -1210 8605
rect -1190 8585 -1170 8605
rect -1150 8585 -1130 8605
rect -1110 8585 -1090 8605
rect -1070 8585 -1050 8605
rect -1030 8585 -1010 8605
rect -990 8585 -970 8605
rect -950 8585 -930 8605
rect -910 8585 -890 8605
rect -870 8585 -850 8605
rect -830 8585 -810 8605
rect -790 8585 -770 8605
rect -750 8585 -730 8605
rect -710 8585 -690 8605
rect -670 8585 -650 8605
rect -630 8585 -610 8605
rect -590 8585 -570 8605
rect -550 8585 -530 8605
rect -510 8585 -490 8605
rect -470 8585 -450 8605
rect -430 8585 -410 8605
rect -390 8585 -370 8605
rect -350 8585 -330 8605
rect -310 8585 -290 8605
rect -270 8585 -250 8605
rect -230 8585 -210 8605
rect -190 8585 -170 8605
rect -150 8585 -130 8605
rect -110 8585 -90 8605
rect -70 8585 -50 8605
rect -30 8585 -10 8605
rect 10 8585 30 8605
rect 50 8585 70 8605
rect 90 8585 110 8605
rect 130 8585 150 8605
rect 170 8585 190 8605
rect 210 8585 230 8605
rect 250 8585 270 8605
rect 290 8585 310 8605
rect 330 8585 350 8605
rect 370 8585 390 8605
rect 410 8585 430 8605
rect 450 8585 470 8605
rect 490 8585 510 8605
rect 530 8585 550 8605
rect 570 8585 635 8605
rect -2225 8570 635 8585
rect -2225 8550 -2210 8570
rect -2190 8550 -2175 8570
rect -2225 8530 -2175 8550
rect 585 8550 600 8570
rect 620 8550 635 8570
rect 585 8530 635 8550
rect -2225 8510 -2210 8530
rect -2190 8510 -2175 8530
rect -2225 8490 -2175 8510
rect -2225 8470 -2210 8490
rect -2190 8470 -2175 8490
rect -2225 8450 -2175 8470
rect -2225 8430 -2210 8450
rect -2190 8430 -2175 8450
rect -2225 8410 -2175 8430
rect -2225 8390 -2210 8410
rect -2190 8390 -2175 8410
rect 585 8510 600 8530
rect 620 8510 635 8530
rect 585 8490 635 8510
rect 585 8470 600 8490
rect 620 8470 635 8490
rect 585 8450 635 8470
rect 585 8430 600 8450
rect 620 8430 635 8450
rect 585 8410 635 8430
rect -2225 8370 -2175 8390
rect -2225 8350 -2210 8370
rect -2190 8350 -2175 8370
rect -2225 8330 -2175 8350
rect -2225 8310 -2210 8330
rect -2190 8310 -2175 8330
rect 585 8390 600 8410
rect 620 8390 635 8410
rect 585 8370 635 8390
rect 585 8350 600 8370
rect 620 8350 635 8370
rect 585 8330 635 8350
rect -2225 8290 -2175 8310
rect -2225 8270 -2210 8290
rect -2190 8270 -2175 8290
rect -2225 8250 -2175 8270
rect -2225 8230 -2210 8250
rect -2190 8230 -2175 8250
rect 585 8310 600 8330
rect 620 8310 635 8330
rect 585 8290 635 8310
rect 585 8270 600 8290
rect 620 8270 635 8290
rect 585 8250 635 8270
rect -2225 8210 -2175 8230
rect -2225 8190 -2210 8210
rect -2190 8190 -2175 8210
rect -2225 8170 -2175 8190
rect -2225 8150 -2210 8170
rect -2190 8150 -2175 8170
rect 585 8230 600 8250
rect 620 8230 635 8250
rect 585 8210 635 8230
rect 585 8190 600 8210
rect 620 8190 635 8210
rect 585 8170 635 8190
rect -2225 8130 -2175 8150
rect -2225 8110 -2210 8130
rect -2190 8110 -2175 8130
rect -2225 8090 -2175 8110
rect -2225 8070 -2210 8090
rect -2190 8070 -2175 8090
rect 585 8150 600 8170
rect 620 8150 635 8170
rect 585 8130 635 8150
rect 585 8110 600 8130
rect 620 8110 635 8130
rect 585 8090 635 8110
rect -2225 8050 -2175 8070
rect -2225 8030 -2210 8050
rect -2190 8030 -2175 8050
rect -2225 8010 -2175 8030
rect -2225 7990 -2210 8010
rect -2190 7990 -2175 8010
rect 585 8070 600 8090
rect 620 8070 635 8090
rect 585 8050 635 8070
rect 585 8030 600 8050
rect 620 8030 635 8050
rect 585 8010 635 8030
rect -2225 7970 -2175 7990
rect -2225 7950 -2210 7970
rect -2190 7950 -2175 7970
rect -2225 7930 -2175 7950
rect -2225 7910 -2210 7930
rect -2190 7910 -2175 7930
rect 585 7990 600 8010
rect 620 7990 635 8010
rect 585 7970 635 7990
rect 585 7950 600 7970
rect 620 7950 635 7970
rect 585 7930 635 7950
rect -2225 7890 -2175 7910
rect -2225 7870 -2210 7890
rect -2190 7870 -2175 7890
rect -2225 7850 -2175 7870
rect -2225 7830 -2210 7850
rect -2190 7830 -2175 7850
rect 585 7910 600 7930
rect 620 7910 635 7930
rect 585 7890 635 7910
rect 585 7870 600 7890
rect 620 7870 635 7890
rect 585 7850 635 7870
rect -2225 7810 -2175 7830
rect -2225 7790 -2210 7810
rect -2190 7790 -2175 7810
rect -2225 7770 -2175 7790
rect -2225 7750 -2210 7770
rect -2190 7750 -2175 7770
rect 585 7830 600 7850
rect 620 7830 635 7850
rect 585 7810 635 7830
rect 585 7790 600 7810
rect 620 7790 635 7810
rect 585 7770 635 7790
rect -2225 7730 -2175 7750
rect -2225 7710 -2210 7730
rect -2190 7710 -2175 7730
rect -2225 7690 -2175 7710
rect -2225 7670 -2210 7690
rect -2190 7670 -2175 7690
rect 585 7750 600 7770
rect 620 7750 635 7770
rect 585 7730 635 7750
rect 585 7710 600 7730
rect 620 7710 635 7730
rect 585 7690 635 7710
rect -2225 7650 -2175 7670
rect -2225 7630 -2210 7650
rect -2190 7630 -2175 7650
rect -2225 7610 -2175 7630
rect -2225 7590 -2210 7610
rect -2190 7590 -2175 7610
rect -2225 7570 -2175 7590
rect 585 7670 600 7690
rect 620 7670 635 7690
rect 585 7650 635 7670
rect 585 7630 600 7650
rect 620 7630 635 7650
rect 585 7610 635 7630
rect 585 7590 600 7610
rect 620 7590 635 7610
rect -2225 7550 -2210 7570
rect -2190 7550 -2175 7570
rect -2225 7530 -2175 7550
rect -2225 7510 -2210 7530
rect -2190 7510 -2175 7530
rect -2225 7490 -2175 7510
rect 585 7570 635 7590
rect 585 7550 600 7570
rect 620 7550 635 7570
rect 585 7530 635 7550
rect 585 7510 600 7530
rect 620 7510 635 7530
rect -2225 7470 -2210 7490
rect -2190 7470 -2175 7490
rect -2225 7450 -2175 7470
rect -2225 7430 -2210 7450
rect -2190 7430 -2175 7450
rect -2225 7410 -2175 7430
rect 585 7490 635 7510
rect 585 7470 600 7490
rect 620 7470 635 7490
rect 585 7450 635 7470
rect 585 7430 600 7450
rect 620 7430 635 7450
rect -2225 7390 -2210 7410
rect -2190 7390 -2175 7410
rect -2225 7370 -2175 7390
rect -2225 7350 -2210 7370
rect -2190 7350 -2175 7370
rect -2225 7330 -2175 7350
rect 585 7410 635 7430
rect 585 7390 600 7410
rect 620 7390 635 7410
rect 585 7370 635 7390
rect 585 7350 600 7370
rect 620 7350 635 7370
rect -2225 7310 -2210 7330
rect -2190 7310 -2175 7330
rect -2225 7290 -2175 7310
rect -2225 7270 -2210 7290
rect -2190 7270 -2175 7290
rect -2225 7250 -2175 7270
rect 585 7330 635 7350
rect 585 7310 600 7330
rect 620 7310 635 7330
rect 585 7290 635 7310
rect 585 7270 600 7290
rect 620 7270 635 7290
rect -2225 7230 -2210 7250
rect -2190 7230 -2175 7250
rect -2225 7210 -2175 7230
rect -2225 7190 -2210 7210
rect -2190 7190 -2175 7210
rect -2225 7170 -2175 7190
rect 585 7250 635 7270
rect 585 7230 600 7250
rect 620 7230 635 7250
rect 585 7210 635 7230
rect 585 7190 600 7210
rect 620 7190 635 7210
rect -2225 7150 -2210 7170
rect -2190 7150 -2175 7170
rect -2225 7130 -2175 7150
rect -2225 7110 -2210 7130
rect -2190 7110 -2175 7130
rect -2225 7090 -2175 7110
rect 585 7170 635 7190
rect 585 7150 600 7170
rect 620 7150 635 7170
rect 585 7130 635 7150
rect 585 7110 600 7130
rect 620 7110 635 7130
rect -2225 7070 -2210 7090
rect -2190 7070 -2175 7090
rect -2225 7050 -2175 7070
rect -2225 7030 -2210 7050
rect -2190 7030 -2175 7050
rect -2225 7010 -2175 7030
rect 585 7090 635 7110
rect 585 7070 600 7090
rect 620 7070 635 7090
rect 585 7050 635 7070
rect 585 7030 600 7050
rect 620 7030 635 7050
rect -2225 6990 -2210 7010
rect -2190 6990 -2175 7010
rect -2225 6970 -2175 6990
rect -2225 6950 -2210 6970
rect -2190 6950 -2175 6970
rect -2225 6930 -2175 6950
rect 585 7010 635 7030
rect 585 6990 600 7010
rect 620 6990 635 7010
rect 585 6970 635 6990
rect 585 6950 600 6970
rect 620 6950 635 6970
rect -2225 6910 -2210 6930
rect -2190 6910 -2175 6930
rect -2225 6890 -2175 6910
rect -2225 6870 -2210 6890
rect -2190 6870 -2175 6890
rect -2225 6850 -2175 6870
rect 585 6930 635 6950
rect 585 6910 600 6930
rect 620 6910 635 6930
rect 585 6890 635 6910
rect 585 6870 600 6890
rect 620 6870 635 6890
rect -2225 6830 -2210 6850
rect -2190 6830 -2175 6850
rect -2225 6810 -2175 6830
rect -2225 6790 -2210 6810
rect -2190 6790 -2175 6810
rect -2225 6770 -2175 6790
rect -2225 6750 -2210 6770
rect -2190 6750 -2175 6770
rect 585 6850 635 6870
rect 585 6830 600 6850
rect 620 6830 635 6850
rect 585 6810 635 6830
rect 585 6790 600 6810
rect 620 6790 635 6810
rect 585 6770 635 6790
rect -2225 6730 -2175 6750
rect -2225 6710 -2210 6730
rect -2190 6710 -2175 6730
rect -2225 6690 -2175 6710
rect -2225 6670 -2210 6690
rect -2190 6670 -2175 6690
rect 585 6750 600 6770
rect 620 6750 635 6770
rect 585 6730 635 6750
rect 585 6710 600 6730
rect 620 6710 635 6730
rect 585 6690 635 6710
rect -2225 6650 -2175 6670
rect -2225 6630 -2210 6650
rect -2190 6630 -2175 6650
rect -2225 6610 -2175 6630
rect -2225 6590 -2210 6610
rect -2190 6590 -2175 6610
rect 585 6670 600 6690
rect 620 6670 635 6690
rect 585 6650 635 6670
rect 585 6630 600 6650
rect 620 6630 635 6650
rect 585 6610 635 6630
rect -2225 6570 -2175 6590
rect -2225 6550 -2210 6570
rect -2190 6550 -2175 6570
rect -2225 6530 -2175 6550
rect -2225 6510 -2210 6530
rect -2190 6510 -2175 6530
rect 585 6590 600 6610
rect 620 6590 635 6610
rect 585 6570 635 6590
rect 585 6550 600 6570
rect 620 6550 635 6570
rect 585 6530 635 6550
rect -2225 6490 -2175 6510
rect -2225 6470 -2210 6490
rect -2190 6470 -2175 6490
rect -2225 6450 -2175 6470
rect -2225 6430 -2210 6450
rect -2190 6430 -2175 6450
rect 585 6510 600 6530
rect 620 6510 635 6530
rect 585 6490 635 6510
rect 585 6470 600 6490
rect 620 6470 635 6490
rect 585 6450 635 6470
rect -2225 6410 -2175 6430
rect -2225 6390 -2210 6410
rect -2190 6390 -2175 6410
rect -2225 6370 -2175 6390
rect -2225 6350 -2210 6370
rect -2190 6350 -2175 6370
rect 585 6430 600 6450
rect 620 6430 635 6450
rect 585 6410 635 6430
rect 585 6390 600 6410
rect 620 6390 635 6410
rect 585 6370 635 6390
rect -2225 6330 -2175 6350
rect -2225 6310 -2210 6330
rect -2190 6310 -2175 6330
rect -2225 6290 -2175 6310
rect -2225 6270 -2210 6290
rect -2190 6270 -2175 6290
rect 585 6350 600 6370
rect 620 6350 635 6370
rect 585 6330 635 6350
rect 585 6310 600 6330
rect 620 6310 635 6330
rect 585 6290 635 6310
rect -2225 6250 -2175 6270
rect -2225 6230 -2210 6250
rect -2190 6235 -2175 6250
rect 585 6270 600 6290
rect 620 6270 635 6290
rect 585 6250 635 6270
rect 585 6235 600 6250
rect -2190 6230 600 6235
rect 620 6230 635 6250
rect -2225 6220 635 6230
rect -2225 6200 -2170 6220
rect -2150 6200 -2130 6220
rect -2110 6200 -2090 6220
rect -2070 6200 -2050 6220
rect -2030 6200 -2010 6220
rect -1990 6200 -1970 6220
rect -1950 6200 -1930 6220
rect -1910 6200 -1890 6220
rect -1870 6200 -1850 6220
rect -1830 6200 -1810 6220
rect -1790 6200 -1770 6220
rect -1750 6200 -1730 6220
rect -1710 6200 -1690 6220
rect -1670 6200 -1650 6220
rect -1630 6200 -1610 6220
rect -1590 6200 -1570 6220
rect -1550 6200 -1530 6220
rect -1510 6200 -1490 6220
rect -1470 6200 -1450 6220
rect -1430 6200 -1410 6220
rect -1390 6200 -1370 6220
rect -1350 6200 -1330 6220
rect -1310 6200 -1290 6220
rect -1270 6200 -1250 6220
rect -1230 6200 -1210 6220
rect -1190 6200 -1170 6220
rect -1150 6200 -1130 6220
rect -1110 6200 -1090 6220
rect -1070 6200 -1050 6220
rect -1030 6200 -1010 6220
rect -990 6200 -970 6220
rect -950 6200 -930 6220
rect -910 6200 -890 6220
rect -870 6200 -850 6220
rect -830 6200 -810 6220
rect -790 6200 -770 6220
rect -750 6200 -730 6220
rect -710 6200 -690 6220
rect -670 6200 -650 6220
rect -630 6200 -610 6220
rect -590 6200 -570 6220
rect -550 6200 -530 6220
rect -510 6200 -490 6220
rect -470 6200 -450 6220
rect -430 6200 -410 6220
rect -390 6200 -370 6220
rect -350 6200 -330 6220
rect -310 6200 -290 6220
rect -270 6200 -250 6220
rect -230 6200 -210 6220
rect -190 6200 -170 6220
rect -150 6200 -130 6220
rect -110 6200 -90 6220
rect -70 6200 -50 6220
rect -30 6200 -10 6220
rect 10 6200 30 6220
rect 50 6200 70 6220
rect 90 6200 110 6220
rect 130 6200 150 6220
rect 170 6200 190 6220
rect 210 6200 230 6220
rect 250 6200 270 6220
rect 290 6200 310 6220
rect 330 6200 350 6220
rect 370 6200 390 6220
rect 410 6200 430 6220
rect 450 6200 470 6220
rect 490 6200 510 6220
rect 530 6200 550 6220
rect 570 6200 635 6220
rect -2225 6185 635 6200
<< psubdiffcont >>
rect -5650 8500 -5630 8520
rect -5610 8500 -5590 8520
rect -5570 8500 -5550 8520
rect -5530 8500 -5510 8520
rect -5490 8500 -5470 8520
rect -5450 8500 -5430 8520
rect -5410 8500 -5390 8520
rect -5370 8500 -5350 8520
rect -5330 8500 -5310 8520
rect -5290 8500 -5270 8520
rect -5250 8500 -5230 8520
rect -5210 8500 -5190 8520
rect -5170 8500 -5150 8520
rect -5130 8500 -5110 8520
rect -5090 8500 -5070 8520
rect -5050 8500 -5030 8520
rect -5010 8500 -4990 8520
rect -4970 8500 -4950 8520
rect -4930 8500 -4910 8520
rect -4890 8500 -4870 8520
rect -4850 8500 -4830 8520
rect -4810 8500 -4790 8520
rect -4770 8500 -4750 8520
rect -4730 8500 -4710 8520
rect -4690 8500 -4670 8520
rect -4650 8500 -4630 8520
rect -4610 8500 -4590 8520
rect -4570 8500 -4550 8520
rect -4530 8500 -4510 8520
rect -4490 8500 -4470 8520
rect -4450 8500 -4430 8520
rect -4410 8500 -4390 8520
rect -4370 8500 -4350 8520
rect -4330 8500 -4310 8520
rect -4290 8500 -4270 8520
rect -4250 8500 -4230 8520
rect -4210 8500 -4190 8520
rect -4170 8500 -4150 8520
rect -4130 8500 -4110 8520
rect -4090 8500 -4070 8520
rect -4050 8500 -4030 8520
rect -4010 8500 -3990 8520
rect -3970 8500 -3950 8520
rect -3930 8500 -3910 8520
rect -3890 8500 -3870 8520
rect -3850 8500 -3830 8520
rect -3810 8500 -3790 8520
rect -3770 8500 -3750 8520
rect -3730 8500 -3710 8520
rect -3690 8500 -3670 8520
rect -3650 8500 -3630 8520
rect -3610 8500 -3590 8520
rect -3570 8500 -3550 8520
rect -3530 8500 -3510 8520
rect -3490 8500 -3470 8520
rect -3450 8500 -3430 8520
rect -3410 8500 -3390 8520
rect -3370 8500 -3350 8520
rect -3330 8500 -3310 8520
rect -3290 8500 -3270 8520
rect -3250 8500 -3230 8520
rect -3210 8500 -3190 8520
rect -5650 6285 -5630 6305
rect -5610 6285 -5590 6305
rect -5570 6285 -5550 6305
rect -5530 6285 -5510 6305
rect -5490 6285 -5470 6305
rect -5450 6285 -5430 6305
rect -5410 6285 -5390 6305
rect -5370 6285 -5350 6305
rect -5330 6285 -5310 6305
rect -5290 6285 -5270 6305
rect -5250 6285 -5230 6305
rect -5210 6285 -5190 6305
rect -5170 6285 -5150 6305
rect -5130 6285 -5110 6305
rect -5090 6285 -5070 6305
rect -5050 6285 -5030 6305
rect -5010 6285 -4990 6305
rect -4970 6285 -4950 6305
rect -4930 6285 -4910 6305
rect -4890 6285 -4870 6305
rect -4850 6285 -4830 6305
rect -4810 6285 -4790 6305
rect -4770 6285 -4750 6305
rect -4730 6285 -4710 6305
rect -4690 6285 -4670 6305
rect -4650 6285 -4630 6305
rect -4610 6285 -4590 6305
rect -4570 6285 -4550 6305
rect -4530 6285 -4510 6305
rect -4490 6285 -4470 6305
rect -4450 6285 -4430 6305
rect -4410 6285 -4390 6305
rect -4370 6285 -4350 6305
rect -4330 6285 -4310 6305
rect -4290 6285 -4270 6305
rect -4250 6285 -4230 6305
rect -4210 6285 -4190 6305
rect -4170 6285 -4150 6305
rect -4130 6285 -4110 6305
rect -4090 6285 -4070 6305
rect -4050 6285 -4030 6305
rect -4010 6285 -3990 6305
rect -3970 6285 -3950 6305
rect -3930 6285 -3910 6305
rect -3890 6285 -3870 6305
rect -3850 6285 -3830 6305
rect -3810 6285 -3790 6305
rect -3770 6285 -3750 6305
rect -3730 6285 -3710 6305
rect -3690 6285 -3670 6305
rect -3650 6285 -3630 6305
rect -3610 6285 -3590 6305
rect -3570 6285 -3550 6305
rect -3530 6285 -3510 6305
rect -3490 6285 -3470 6305
rect -3450 6285 -3430 6305
rect -3410 6285 -3390 6305
rect -3370 6285 -3350 6305
rect -3330 6285 -3310 6305
rect -3290 6285 -3270 6305
rect -3250 6285 -3230 6305
rect -3210 6285 -3190 6305
rect -1950 8500 -1930 8520
rect -1910 8500 -1890 8520
rect -1870 8500 -1850 8520
rect -1830 8500 -1810 8520
rect -1790 8500 -1770 8520
rect -1750 8500 -1730 8520
rect -1710 8500 -1690 8520
rect -1670 8500 -1650 8520
rect -1630 8500 -1610 8520
rect -1590 8500 -1570 8520
rect -1550 8500 -1530 8520
rect -1510 8500 -1490 8520
rect -1470 8500 -1450 8520
rect -1430 8500 -1410 8520
rect -1390 8500 -1370 8520
rect -1350 8500 -1330 8520
rect -1310 8500 -1290 8520
rect -1270 8500 -1250 8520
rect -1230 8500 -1210 8520
rect -1190 8500 -1170 8520
rect -1150 8500 -1130 8520
rect -1110 8500 -1090 8520
rect -1070 8500 -1050 8520
rect -1030 8500 -1010 8520
rect -990 8500 -970 8520
rect -950 8500 -930 8520
rect -910 8500 -890 8520
rect -870 8500 -850 8520
rect -830 8500 -810 8520
rect -790 8500 -770 8520
rect -750 8500 -730 8520
rect -710 8500 -690 8520
rect -670 8500 -650 8520
rect -630 8500 -610 8520
rect -590 8500 -570 8520
rect -550 8500 -530 8520
rect -510 8500 -490 8520
rect -470 8500 -450 8520
rect -430 8500 -410 8520
rect -390 8500 -370 8520
rect -350 8500 -330 8520
rect -310 8500 -290 8520
rect -270 8500 -250 8520
rect -230 8500 -210 8520
rect -190 8500 -170 8520
rect -150 8500 -130 8520
rect -110 8500 -90 8520
rect -70 8500 -50 8520
rect -30 8500 -10 8520
rect 10 8500 30 8520
rect 50 8500 70 8520
rect 90 8500 110 8520
rect 130 8500 150 8520
rect 170 8500 190 8520
rect 210 8500 230 8520
rect 250 8500 270 8520
rect 290 8500 310 8520
rect 330 8500 350 8520
rect 370 8500 390 8520
rect 410 8500 430 8520
rect 450 8500 470 8520
rect 490 8500 510 8520
rect -1950 6285 -1930 6305
rect -1910 6285 -1890 6305
rect -1870 6285 -1850 6305
rect -1830 6285 -1810 6305
rect -1790 6285 -1770 6305
rect -1750 6285 -1730 6305
rect -1710 6285 -1690 6305
rect -1670 6285 -1650 6305
rect -1630 6285 -1610 6305
rect -1590 6285 -1570 6305
rect -1550 6285 -1530 6305
rect -1510 6285 -1490 6305
rect -1470 6285 -1450 6305
rect -1430 6285 -1410 6305
rect -1390 6285 -1370 6305
rect -1350 6285 -1330 6305
rect -1310 6285 -1290 6305
rect -1270 6285 -1250 6305
rect -1230 6285 -1210 6305
rect -1190 6285 -1170 6305
rect -1150 6285 -1130 6305
rect -1110 6285 -1090 6305
rect -1070 6285 -1050 6305
rect -1030 6285 -1010 6305
rect -990 6285 -970 6305
rect -950 6285 -930 6305
rect -910 6285 -890 6305
rect -870 6285 -850 6305
rect -830 6285 -810 6305
rect -790 6285 -770 6305
rect -750 6285 -730 6305
rect -710 6285 -690 6305
rect -670 6285 -650 6305
rect -630 6285 -610 6305
rect -590 6285 -570 6305
rect -550 6285 -530 6305
rect -510 6285 -490 6305
rect -470 6285 -450 6305
rect -430 6285 -410 6305
rect -390 6285 -370 6305
rect -350 6285 -330 6305
rect -310 6285 -290 6305
rect -270 6285 -250 6305
rect -230 6285 -210 6305
rect -190 6285 -170 6305
rect -150 6285 -130 6305
rect -110 6285 -90 6305
rect -70 6285 -50 6305
rect -30 6285 -10 6305
rect 10 6285 30 6305
rect 50 6285 70 6305
rect 90 6285 110 6305
rect 130 6285 150 6305
rect 170 6285 190 6305
rect 210 6285 230 6305
rect 250 6285 270 6305
rect 290 6285 310 6305
rect 330 6285 350 6305
rect 370 6285 390 6305
rect 410 6285 430 6305
rect 450 6285 470 6305
rect 490 6285 510 6305
rect -5580 6065 -5550 6085
rect -5530 6065 -5510 6085
rect -5490 6065 -5470 6085
rect -5450 6065 -5430 6085
rect -5410 6065 -5390 6085
rect -5370 6065 -5350 6085
rect -5330 6065 -5310 6085
rect -5290 6065 -5270 6085
rect -5250 6065 -5230 6085
rect -5210 6065 -5190 6085
rect -5170 6065 -5150 6085
rect -5130 6065 -5110 6085
rect -5090 6065 -5070 6085
rect -5050 6065 -5030 6085
rect -5010 6065 -4990 6085
rect -4970 6065 -4950 6085
rect -4930 6065 -4910 6085
rect -4890 6065 -4870 6085
rect -4850 6065 -4830 6085
rect -4810 6065 -4790 6085
rect -4770 6065 -4750 6085
rect -4730 6065 -4710 6085
rect -4690 6065 -4670 6085
rect -4650 6065 -4630 6085
rect -4610 6065 -4590 6085
rect -4570 6065 -4550 6085
rect -4530 6065 -4510 6085
rect -4490 6065 -4470 6085
rect -4450 6065 -4430 6085
rect -4410 6065 -4390 6085
rect -4370 6065 -4350 6085
rect -4330 6065 -4310 6085
rect -4290 6065 -4270 6085
rect -4250 6065 -4230 6085
rect -4210 6065 -4190 6085
rect -4170 6065 -4150 6085
rect -4130 6065 -4110 6085
rect -4090 6065 -4070 6085
rect -4050 6065 -4030 6085
rect -4010 6065 -3990 6085
rect -3970 6065 -3950 6085
rect -3930 6065 -3910 6085
rect -3890 6065 -3870 6085
rect -3850 6065 -3830 6085
rect -3810 6065 -3790 6085
rect -3770 6065 -3750 6085
rect -3730 6065 -3710 6085
rect -3690 6065 -3670 6085
rect -3650 6065 -3630 6085
rect -3610 6065 -3590 6085
rect -3570 6065 -3550 6085
rect -3530 6065 -3510 6085
rect -3490 6065 -3470 6085
rect -3450 6065 -3430 6085
rect -3410 6065 -3390 6085
rect -3370 6065 -3350 6085
rect -3330 6065 -3310 6085
rect -3290 6065 -3270 6085
rect -3250 6065 -3230 6085
rect -3210 6065 -3190 6085
rect -3170 6065 -3150 6085
rect -3130 6065 -3110 6085
rect -2030 6065 -2010 6085
rect -1990 6065 -1970 6085
rect -1950 6065 -1930 6085
rect -1910 6065 -1890 6085
rect -1870 6065 -1850 6085
rect -1830 6065 -1810 6085
rect -1790 6065 -1770 6085
rect -1750 6065 -1730 6085
rect -1710 6065 -1690 6085
rect -1670 6065 -1650 6085
rect -1630 6065 -1610 6085
rect -1590 6065 -1570 6085
rect -1550 6065 -1530 6085
rect -1510 6065 -1490 6085
rect -1470 6065 -1450 6085
rect -1430 6065 -1410 6085
rect -1390 6065 -1370 6085
rect -1350 6065 -1330 6085
rect -1310 6065 -1290 6085
rect -1270 6065 -1250 6085
rect -1230 6065 -1210 6085
rect -1190 6065 -1170 6085
rect -1150 6065 -1130 6085
rect -1110 6065 -1090 6085
rect -1070 6065 -1050 6085
rect -1030 6065 -1010 6085
rect -990 6065 -970 6085
rect -950 6065 -930 6085
rect -910 6065 -890 6085
rect -870 6065 -850 6085
rect -830 6065 -810 6085
rect -790 6065 -770 6085
rect -750 6065 -730 6085
rect -710 6065 -690 6085
rect -670 6065 -650 6085
rect -630 6065 -610 6085
rect -590 6065 -570 6085
rect -550 6065 -530 6085
rect -510 6065 -490 6085
rect -470 6065 -450 6085
rect -430 6065 -410 6085
rect -390 6065 -370 6085
rect -350 6065 -330 6085
rect -310 6065 -290 6085
rect -270 6065 -250 6085
rect -230 6065 -210 6085
rect -190 6065 -170 6085
rect -150 6065 -130 6085
rect -110 6065 -90 6085
rect -70 6065 -50 6085
rect -30 6065 -10 6085
rect 10 6065 30 6085
rect 50 6065 70 6085
rect 90 6065 110 6085
rect 130 6065 150 6085
rect 170 6065 190 6085
rect 210 6065 230 6085
rect 250 6065 270 6085
rect 290 6065 310 6085
rect 330 6065 350 6085
rect 370 6065 390 6085
rect 410 6065 440 6085
rect -5580 3515 -5550 3535
rect -5530 3515 -5510 3535
rect -5490 3515 -5470 3535
rect -5450 3515 -5430 3535
rect -5410 3515 -5390 3535
rect -5370 3515 -5350 3535
rect -5330 3515 -5310 3535
rect -5290 3515 -5270 3535
rect -5250 3515 -5230 3535
rect -5210 3515 -5190 3535
rect -5170 3515 -5150 3535
rect -5130 3515 -5110 3535
rect -5090 3515 -5070 3535
rect -5050 3515 -5030 3535
rect -5010 3515 -4990 3535
rect -4970 3515 -4950 3535
rect -4930 3515 -4910 3535
rect -4890 3515 -4870 3535
rect -4850 3515 -4830 3535
rect -4810 3515 -4790 3535
rect -4770 3515 -4750 3535
rect -4730 3515 -4710 3535
rect -4690 3515 -4670 3535
rect -4650 3515 -4630 3535
rect -4610 3515 -4590 3535
rect -4570 3515 -4550 3535
rect -4530 3515 -4510 3535
rect -4490 3515 -4470 3535
rect -4450 3515 -4430 3535
rect -4410 3515 -4390 3535
rect -4370 3515 -4350 3535
rect -4330 3515 -4310 3535
rect -4290 3515 -4270 3535
rect -4250 3515 -4230 3535
rect -4210 3515 -4190 3535
rect -4170 3515 -4150 3535
rect -4130 3515 -4110 3535
rect -4090 3515 -4070 3535
rect -4050 3515 -4030 3535
rect -4010 3515 -3990 3535
rect -3970 3515 -3950 3535
rect -3930 3515 -3910 3535
rect -3890 3515 -3870 3535
rect -3850 3515 -3830 3535
rect -3810 3515 -3790 3535
rect -3770 3515 -3750 3535
rect -3730 3515 -3710 3535
rect -3690 3515 -3670 3535
rect -3650 3515 -3630 3535
rect -3610 3515 -3590 3535
rect -3570 3515 -3550 3535
rect -3530 3515 -3510 3535
rect -3490 3515 -3470 3535
rect -3450 3515 -3430 3535
rect -3410 3515 -3390 3535
rect -3370 3515 -3350 3535
rect -3330 3515 -3310 3535
rect -3290 3515 -3270 3535
rect -3250 3515 -3230 3535
rect -3210 3515 -3190 3535
rect -3170 3515 -3150 3535
rect -3130 3515 -3110 3535
rect -2030 3515 -2010 3535
rect -1990 3515 -1970 3535
rect -1950 3515 -1930 3535
rect -1910 3515 -1890 3535
rect -1870 3515 -1850 3535
rect -1830 3515 -1810 3535
rect -1790 3515 -1770 3535
rect -1750 3515 -1730 3535
rect -1710 3515 -1690 3535
rect -1670 3515 -1650 3535
rect -1630 3515 -1610 3535
rect -1590 3515 -1570 3535
rect -1550 3515 -1530 3535
rect -1510 3515 -1490 3535
rect -1470 3515 -1450 3535
rect -1430 3515 -1410 3535
rect -1390 3515 -1370 3535
rect -1350 3515 -1330 3535
rect -1310 3515 -1290 3535
rect -1270 3515 -1250 3535
rect -1230 3515 -1210 3535
rect -1190 3515 -1170 3535
rect -1150 3515 -1130 3535
rect -1110 3515 -1090 3535
rect -1070 3515 -1050 3535
rect -1030 3515 -1010 3535
rect -990 3515 -970 3535
rect -950 3515 -930 3535
rect -910 3515 -890 3535
rect -870 3515 -850 3535
rect -830 3515 -810 3535
rect -790 3515 -770 3535
rect -750 3515 -730 3535
rect -710 3515 -690 3535
rect -670 3515 -650 3535
rect -630 3515 -610 3535
rect -590 3515 -570 3535
rect -550 3515 -530 3535
rect -510 3515 -490 3535
rect -470 3515 -450 3535
rect -430 3515 -410 3535
rect -390 3515 -370 3535
rect -350 3515 -330 3535
rect -310 3515 -290 3535
rect -270 3515 -250 3535
rect -230 3515 -210 3535
rect -190 3515 -170 3535
rect -150 3515 -130 3535
rect -110 3515 -90 3535
rect -70 3515 -50 3535
rect -30 3515 -10 3535
rect 10 3515 30 3535
rect 50 3515 70 3535
rect 90 3515 110 3535
rect 130 3515 150 3535
rect 170 3515 190 3535
rect 210 3515 230 3535
rect 250 3515 270 3535
rect 290 3515 310 3535
rect 330 3515 350 3535
rect 370 3515 390 3535
rect 410 3515 440 3535
<< nsubdiffcont >>
rect -5710 8585 -5690 8605
rect -5670 8585 -5650 8605
rect -5630 8585 -5610 8605
rect -5590 8585 -5570 8605
rect -5550 8585 -5530 8605
rect -5510 8585 -5490 8605
rect -5470 8585 -5450 8605
rect -5430 8585 -5410 8605
rect -5390 8585 -5370 8605
rect -5350 8585 -5330 8605
rect -5310 8585 -5290 8605
rect -5270 8585 -5250 8605
rect -5230 8585 -5210 8605
rect -5190 8585 -5170 8605
rect -5150 8585 -5130 8605
rect -5110 8585 -5090 8605
rect -5070 8585 -5050 8605
rect -5030 8585 -5010 8605
rect -4990 8585 -4970 8605
rect -4950 8585 -4930 8605
rect -4910 8585 -4890 8605
rect -4870 8585 -4850 8605
rect -4830 8585 -4810 8605
rect -4790 8585 -4770 8605
rect -4750 8585 -4730 8605
rect -4710 8585 -4690 8605
rect -4670 8585 -4650 8605
rect -4630 8585 -4610 8605
rect -4590 8585 -4570 8605
rect -4550 8585 -4530 8605
rect -4510 8585 -4490 8605
rect -4470 8585 -4450 8605
rect -4430 8585 -4410 8605
rect -4390 8585 -4370 8605
rect -4350 8585 -4330 8605
rect -4310 8585 -4290 8605
rect -4270 8585 -4250 8605
rect -4230 8585 -4210 8605
rect -4190 8585 -4170 8605
rect -4150 8585 -4130 8605
rect -4110 8585 -4090 8605
rect -4070 8585 -4050 8605
rect -4030 8585 -4010 8605
rect -3990 8585 -3970 8605
rect -3950 8585 -3930 8605
rect -3910 8585 -3890 8605
rect -3870 8585 -3850 8605
rect -3830 8585 -3810 8605
rect -3790 8585 -3770 8605
rect -3750 8585 -3730 8605
rect -3710 8585 -3690 8605
rect -3670 8585 -3650 8605
rect -3630 8585 -3610 8605
rect -3590 8585 -3570 8605
rect -3550 8585 -3530 8605
rect -3510 8585 -3490 8605
rect -3470 8585 -3450 8605
rect -3430 8585 -3410 8605
rect -3390 8585 -3370 8605
rect -3350 8585 -3330 8605
rect -3310 8585 -3290 8605
rect -3270 8585 -3250 8605
rect -3230 8585 -3210 8605
rect -3190 8585 -3170 8605
rect -3150 8585 -3130 8605
rect -3110 8585 -3090 8605
rect -3070 8585 -3050 8605
rect -3030 8585 -3010 8605
rect -2990 8585 -2970 8605
rect -5760 8550 -5740 8570
rect -2950 8550 -2930 8570
rect -5760 8510 -5740 8530
rect -5760 8470 -5740 8490
rect -5760 8430 -5740 8450
rect -2950 8510 -2930 8530
rect -2950 8470 -2930 8490
rect -5760 8390 -5740 8410
rect -5760 8350 -5740 8370
rect -2950 8430 -2930 8450
rect -2950 8390 -2930 8410
rect -5760 8310 -5740 8330
rect -5760 8270 -5740 8290
rect -2950 8350 -2930 8370
rect -2950 8310 -2930 8330
rect -5760 8230 -5740 8250
rect -5760 8190 -5740 8210
rect -2950 8270 -2930 8290
rect -2950 8230 -2930 8250
rect -5760 8150 -5740 8170
rect -5760 8110 -5740 8130
rect -2950 8190 -2930 8210
rect -2950 8150 -2930 8170
rect -5760 8070 -5740 8090
rect -5760 8030 -5740 8050
rect -2950 8110 -2930 8130
rect -2950 8070 -2930 8090
rect -5760 7990 -5740 8010
rect -5760 7950 -5740 7970
rect -2950 8030 -2930 8050
rect -2950 7990 -2930 8010
rect -5760 7910 -5740 7930
rect -5760 7870 -5740 7890
rect -2950 7950 -2930 7970
rect -2950 7910 -2930 7930
rect -2950 7870 -2930 7890
rect -5760 7830 -5740 7850
rect -5760 7790 -5740 7810
rect -2950 7830 -2930 7850
rect -2950 7790 -2930 7810
rect -5760 7750 -5740 7770
rect -5760 7710 -5740 7730
rect -2950 7750 -2930 7770
rect -2950 7710 -2930 7730
rect -5760 7670 -5740 7690
rect -5760 7630 -5740 7650
rect -2950 7670 -2930 7690
rect -2950 7630 -2930 7650
rect -5760 7590 -5740 7610
rect -5760 7550 -5740 7570
rect -2950 7590 -2930 7610
rect -2950 7550 -2930 7570
rect -5760 7510 -5740 7530
rect -5760 7470 -5740 7490
rect -2950 7510 -2930 7530
rect -2950 7470 -2930 7490
rect -5760 7430 -5740 7450
rect -5760 7390 -5740 7410
rect -2950 7430 -2930 7450
rect -2950 7390 -2930 7410
rect -5760 7350 -5740 7370
rect -5760 7310 -5740 7330
rect -2950 7350 -2930 7370
rect -2950 7310 -2930 7330
rect -5760 7270 -5740 7290
rect -5760 7230 -5740 7250
rect -2950 7270 -2930 7290
rect -2950 7230 -2930 7250
rect -5760 7190 -5740 7210
rect -5760 7150 -5740 7170
rect -2950 7190 -2930 7210
rect -2950 7150 -2930 7170
rect -5760 7110 -5740 7130
rect -5760 7070 -5740 7090
rect -5760 7030 -5740 7050
rect -2950 7110 -2930 7130
rect -2950 7070 -2930 7090
rect -5760 6990 -5740 7010
rect -5760 6950 -5740 6970
rect -2950 7030 -2930 7050
rect -2950 6990 -2930 7010
rect -5760 6910 -5740 6930
rect -5760 6870 -5740 6890
rect -2950 6950 -2930 6970
rect -2950 6910 -2930 6930
rect -5760 6830 -5740 6850
rect -5760 6790 -5740 6810
rect -2950 6870 -2930 6890
rect -2950 6830 -2930 6850
rect -5760 6750 -5740 6770
rect -5760 6710 -5740 6730
rect -2950 6790 -2930 6810
rect -2950 6750 -2930 6770
rect -5760 6670 -5740 6690
rect -5760 6630 -5740 6650
rect -2950 6710 -2930 6730
rect -2950 6670 -2930 6690
rect -5760 6590 -5740 6610
rect -5760 6550 -5740 6570
rect -2950 6630 -2930 6650
rect -2950 6590 -2930 6610
rect -5760 6510 -5740 6530
rect -5760 6470 -5740 6490
rect -2950 6550 -2930 6570
rect -2950 6510 -2930 6530
rect -5760 6430 -5740 6450
rect -5760 6390 -5740 6410
rect -2950 6470 -2930 6490
rect -2950 6430 -2930 6450
rect -5760 6350 -5740 6370
rect -2950 6390 -2930 6410
rect -5760 6310 -5740 6330
rect -5760 6270 -5740 6290
rect -2950 6350 -2930 6370
rect -2950 6310 -2930 6330
rect -5760 6230 -5740 6250
rect -2950 6270 -2930 6290
rect -2950 6230 -2930 6250
rect -5710 6200 -5690 6220
rect -5670 6200 -5650 6220
rect -5630 6200 -5610 6220
rect -5590 6200 -5570 6220
rect -5550 6200 -5530 6220
rect -5510 6200 -5490 6220
rect -5470 6200 -5450 6220
rect -5430 6200 -5410 6220
rect -5390 6200 -5370 6220
rect -5350 6200 -5330 6220
rect -5310 6200 -5290 6220
rect -5270 6200 -5250 6220
rect -5230 6200 -5210 6220
rect -5190 6200 -5170 6220
rect -5150 6200 -5130 6220
rect -5110 6200 -5090 6220
rect -5070 6200 -5050 6220
rect -5030 6200 -5010 6220
rect -4990 6200 -4970 6220
rect -4950 6200 -4930 6220
rect -4910 6200 -4890 6220
rect -4870 6200 -4850 6220
rect -4830 6200 -4810 6220
rect -4790 6200 -4770 6220
rect -4750 6200 -4730 6220
rect -4710 6200 -4690 6220
rect -4670 6200 -4650 6220
rect -4630 6200 -4610 6220
rect -4590 6200 -4570 6220
rect -4550 6200 -4530 6220
rect -4510 6200 -4490 6220
rect -4470 6200 -4450 6220
rect -4430 6200 -4410 6220
rect -4390 6200 -4370 6220
rect -4350 6200 -4330 6220
rect -4310 6200 -4290 6220
rect -4270 6200 -4250 6220
rect -4230 6200 -4210 6220
rect -4190 6200 -4170 6220
rect -4150 6200 -4130 6220
rect -4110 6200 -4090 6220
rect -4070 6200 -4050 6220
rect -4030 6200 -4010 6220
rect -3990 6200 -3970 6220
rect -3950 6200 -3930 6220
rect -3910 6200 -3890 6220
rect -3870 6200 -3850 6220
rect -3830 6200 -3810 6220
rect -3790 6200 -3770 6220
rect -3750 6200 -3730 6220
rect -3710 6200 -3690 6220
rect -3670 6200 -3650 6220
rect -3630 6200 -3610 6220
rect -3590 6200 -3570 6220
rect -3550 6200 -3530 6220
rect -3510 6200 -3490 6220
rect -3470 6200 -3450 6220
rect -3430 6200 -3410 6220
rect -3390 6200 -3370 6220
rect -3350 6200 -3330 6220
rect -3310 6200 -3290 6220
rect -3270 6200 -3250 6220
rect -3230 6200 -3210 6220
rect -3190 6200 -3170 6220
rect -3150 6200 -3130 6220
rect -3110 6200 -3090 6220
rect -3070 6200 -3050 6220
rect -3030 6200 -3010 6220
rect -2990 6200 -2970 6220
rect -2170 8585 -2150 8605
rect -2130 8585 -2110 8605
rect -2090 8585 -2070 8605
rect -2050 8585 -2030 8605
rect -2010 8585 -1990 8605
rect -1970 8585 -1950 8605
rect -1930 8585 -1910 8605
rect -1890 8585 -1870 8605
rect -1850 8585 -1830 8605
rect -1810 8585 -1790 8605
rect -1770 8585 -1750 8605
rect -1730 8585 -1710 8605
rect -1690 8585 -1670 8605
rect -1650 8585 -1630 8605
rect -1610 8585 -1590 8605
rect -1570 8585 -1550 8605
rect -1530 8585 -1510 8605
rect -1490 8585 -1470 8605
rect -1450 8585 -1430 8605
rect -1410 8585 -1390 8605
rect -1370 8585 -1350 8605
rect -1330 8585 -1310 8605
rect -1290 8585 -1270 8605
rect -1250 8585 -1230 8605
rect -1210 8585 -1190 8605
rect -1170 8585 -1150 8605
rect -1130 8585 -1110 8605
rect -1090 8585 -1070 8605
rect -1050 8585 -1030 8605
rect -1010 8585 -990 8605
rect -970 8585 -950 8605
rect -930 8585 -910 8605
rect -890 8585 -870 8605
rect -850 8585 -830 8605
rect -810 8585 -790 8605
rect -770 8585 -750 8605
rect -730 8585 -710 8605
rect -690 8585 -670 8605
rect -650 8585 -630 8605
rect -610 8585 -590 8605
rect -570 8585 -550 8605
rect -530 8585 -510 8605
rect -490 8585 -470 8605
rect -450 8585 -430 8605
rect -410 8585 -390 8605
rect -370 8585 -350 8605
rect -330 8585 -310 8605
rect -290 8585 -270 8605
rect -250 8585 -230 8605
rect -210 8585 -190 8605
rect -170 8585 -150 8605
rect -130 8585 -110 8605
rect -90 8585 -70 8605
rect -50 8585 -30 8605
rect -10 8585 10 8605
rect 30 8585 50 8605
rect 70 8585 90 8605
rect 110 8585 130 8605
rect 150 8585 170 8605
rect 190 8585 210 8605
rect 230 8585 250 8605
rect 270 8585 290 8605
rect 310 8585 330 8605
rect 350 8585 370 8605
rect 390 8585 410 8605
rect 430 8585 450 8605
rect 470 8585 490 8605
rect 510 8585 530 8605
rect 550 8585 570 8605
rect -2210 8550 -2190 8570
rect 600 8550 620 8570
rect -2210 8510 -2190 8530
rect -2210 8470 -2190 8490
rect -2210 8430 -2190 8450
rect -2210 8390 -2190 8410
rect 600 8510 620 8530
rect 600 8470 620 8490
rect 600 8430 620 8450
rect -2210 8350 -2190 8370
rect -2210 8310 -2190 8330
rect 600 8390 620 8410
rect 600 8350 620 8370
rect -2210 8270 -2190 8290
rect -2210 8230 -2190 8250
rect 600 8310 620 8330
rect 600 8270 620 8290
rect -2210 8190 -2190 8210
rect -2210 8150 -2190 8170
rect 600 8230 620 8250
rect 600 8190 620 8210
rect -2210 8110 -2190 8130
rect -2210 8070 -2190 8090
rect 600 8150 620 8170
rect 600 8110 620 8130
rect -2210 8030 -2190 8050
rect -2210 7990 -2190 8010
rect 600 8070 620 8090
rect 600 8030 620 8050
rect -2210 7950 -2190 7970
rect -2210 7910 -2190 7930
rect 600 7990 620 8010
rect 600 7950 620 7970
rect -2210 7870 -2190 7890
rect -2210 7830 -2190 7850
rect 600 7910 620 7930
rect 600 7870 620 7890
rect -2210 7790 -2190 7810
rect -2210 7750 -2190 7770
rect 600 7830 620 7850
rect 600 7790 620 7810
rect -2210 7710 -2190 7730
rect -2210 7670 -2190 7690
rect 600 7750 620 7770
rect 600 7710 620 7730
rect -2210 7630 -2190 7650
rect -2210 7590 -2190 7610
rect 600 7670 620 7690
rect 600 7630 620 7650
rect 600 7590 620 7610
rect -2210 7550 -2190 7570
rect -2210 7510 -2190 7530
rect 600 7550 620 7570
rect 600 7510 620 7530
rect -2210 7470 -2190 7490
rect -2210 7430 -2190 7450
rect 600 7470 620 7490
rect 600 7430 620 7450
rect -2210 7390 -2190 7410
rect -2210 7350 -2190 7370
rect 600 7390 620 7410
rect 600 7350 620 7370
rect -2210 7310 -2190 7330
rect -2210 7270 -2190 7290
rect 600 7310 620 7330
rect 600 7270 620 7290
rect -2210 7230 -2190 7250
rect -2210 7190 -2190 7210
rect 600 7230 620 7250
rect 600 7190 620 7210
rect -2210 7150 -2190 7170
rect -2210 7110 -2190 7130
rect 600 7150 620 7170
rect 600 7110 620 7130
rect -2210 7070 -2190 7090
rect -2210 7030 -2190 7050
rect 600 7070 620 7090
rect 600 7030 620 7050
rect -2210 6990 -2190 7010
rect -2210 6950 -2190 6970
rect 600 6990 620 7010
rect 600 6950 620 6970
rect -2210 6910 -2190 6930
rect -2210 6870 -2190 6890
rect 600 6910 620 6930
rect 600 6870 620 6890
rect -2210 6830 -2190 6850
rect -2210 6790 -2190 6810
rect -2210 6750 -2190 6770
rect 600 6830 620 6850
rect 600 6790 620 6810
rect -2210 6710 -2190 6730
rect -2210 6670 -2190 6690
rect 600 6750 620 6770
rect 600 6710 620 6730
rect -2210 6630 -2190 6650
rect -2210 6590 -2190 6610
rect 600 6670 620 6690
rect 600 6630 620 6650
rect -2210 6550 -2190 6570
rect -2210 6510 -2190 6530
rect 600 6590 620 6610
rect 600 6550 620 6570
rect -2210 6470 -2190 6490
rect -2210 6430 -2190 6450
rect 600 6510 620 6530
rect 600 6470 620 6490
rect -2210 6390 -2190 6410
rect -2210 6350 -2190 6370
rect 600 6430 620 6450
rect 600 6390 620 6410
rect -2210 6310 -2190 6330
rect -2210 6270 -2190 6290
rect 600 6350 620 6370
rect 600 6310 620 6330
rect -2210 6230 -2190 6250
rect 600 6270 620 6290
rect 600 6230 620 6250
rect -2170 6200 -2150 6220
rect -2130 6200 -2110 6220
rect -2090 6200 -2070 6220
rect -2050 6200 -2030 6220
rect -2010 6200 -1990 6220
rect -1970 6200 -1950 6220
rect -1930 6200 -1910 6220
rect -1890 6200 -1870 6220
rect -1850 6200 -1830 6220
rect -1810 6200 -1790 6220
rect -1770 6200 -1750 6220
rect -1730 6200 -1710 6220
rect -1690 6200 -1670 6220
rect -1650 6200 -1630 6220
rect -1610 6200 -1590 6220
rect -1570 6200 -1550 6220
rect -1530 6200 -1510 6220
rect -1490 6200 -1470 6220
rect -1450 6200 -1430 6220
rect -1410 6200 -1390 6220
rect -1370 6200 -1350 6220
rect -1330 6200 -1310 6220
rect -1290 6200 -1270 6220
rect -1250 6200 -1230 6220
rect -1210 6200 -1190 6220
rect -1170 6200 -1150 6220
rect -1130 6200 -1110 6220
rect -1090 6200 -1070 6220
rect -1050 6200 -1030 6220
rect -1010 6200 -990 6220
rect -970 6200 -950 6220
rect -930 6200 -910 6220
rect -890 6200 -870 6220
rect -850 6200 -830 6220
rect -810 6200 -790 6220
rect -770 6200 -750 6220
rect -730 6200 -710 6220
rect -690 6200 -670 6220
rect -650 6200 -630 6220
rect -610 6200 -590 6220
rect -570 6200 -550 6220
rect -530 6200 -510 6220
rect -490 6200 -470 6220
rect -450 6200 -430 6220
rect -410 6200 -390 6220
rect -370 6200 -350 6220
rect -330 6200 -310 6220
rect -290 6200 -270 6220
rect -250 6200 -230 6220
rect -210 6200 -190 6220
rect -170 6200 -150 6220
rect -130 6200 -110 6220
rect -90 6200 -70 6220
rect -50 6200 -30 6220
rect -10 6200 10 6220
rect 30 6200 50 6220
rect 70 6200 90 6220
rect 110 6200 130 6220
rect 150 6200 170 6220
rect 190 6200 210 6220
rect 230 6200 250 6220
rect 270 6200 290 6220
rect 310 6200 330 6220
rect 350 6200 370 6220
rect 390 6200 410 6220
rect 430 6200 450 6220
rect 470 6200 490 6220
rect 510 6200 530 6220
rect 550 6200 570 6220
<< poly >>
rect -3155 8442 -2990 8445
rect -5680 8410 -5665 8442
rect -3165 8435 -2990 8442
rect -3165 8415 -3145 8435
rect -3120 8415 -3100 8435
rect -3080 8415 -3060 8435
rect -3040 8415 -3020 8435
rect -3000 8415 -2990 8435
rect -3165 8410 -2990 8415
rect -3155 8405 -2990 8410
rect -3155 8360 -2990 8365
rect -5680 8328 -5665 8360
rect -3165 8355 -2990 8360
rect -3165 8335 -3145 8355
rect -3120 8335 -3100 8355
rect -3080 8335 -3060 8355
rect -3040 8335 -3020 8355
rect -3000 8335 -2990 8355
rect -3165 8328 -2990 8335
rect -3155 8325 -2990 8328
rect -3155 8278 -2990 8280
rect -5680 8246 -5665 8278
rect -3165 8270 -2990 8278
rect -3165 8250 -3145 8270
rect -3120 8250 -3100 8270
rect -3080 8250 -3060 8270
rect -3040 8250 -3020 8270
rect -3000 8250 -2990 8270
rect -3165 8246 -2990 8250
rect -3155 8240 -2990 8246
rect -3155 8196 -2990 8200
rect -5680 8164 -5665 8196
rect -3165 8190 -2990 8196
rect -3165 8170 -3145 8190
rect -3120 8170 -3100 8190
rect -3080 8170 -3060 8190
rect -3040 8170 -3020 8190
rect -3000 8170 -2990 8190
rect -3165 8164 -2990 8170
rect -3155 8160 -2990 8164
rect -3155 8114 -2990 8120
rect -5680 8082 -5665 8114
rect -3165 8110 -2990 8114
rect -3165 8090 -3145 8110
rect -3120 8090 -3100 8110
rect -3080 8090 -3060 8110
rect -3040 8090 -3020 8110
rect -3000 8090 -2990 8110
rect -3165 8082 -2990 8090
rect -3155 8080 -2990 8082
rect -3155 8032 -2990 8035
rect -5680 8000 -5665 8032
rect -3165 8025 -2990 8032
rect -3165 8005 -3145 8025
rect -3120 8005 -3100 8025
rect -3080 8005 -3060 8025
rect -3040 8005 -3020 8025
rect -3000 8005 -2990 8025
rect -3165 8000 -2990 8005
rect -3155 7995 -2990 8000
rect -3155 7950 -2990 7955
rect -5680 7918 -5665 7950
rect -3165 7945 -2990 7950
rect -3165 7925 -3145 7945
rect -3120 7925 -3100 7945
rect -3080 7925 -3060 7945
rect -3040 7925 -3020 7945
rect -3000 7925 -2990 7945
rect -3165 7918 -2990 7925
rect -3155 7915 -2990 7918
rect -3155 7868 -2990 7870
rect -5680 7836 -5665 7868
rect -3165 7860 -2990 7868
rect -3165 7840 -3145 7860
rect -3120 7840 -3100 7860
rect -3080 7840 -3060 7860
rect -3040 7840 -3020 7860
rect -3000 7840 -2990 7860
rect -3165 7836 -2990 7840
rect -3155 7830 -2990 7836
rect -3155 7786 -2990 7790
rect -5680 7754 -5665 7786
rect -3165 7780 -2990 7786
rect -3165 7760 -3145 7780
rect -3120 7760 -3100 7780
rect -3080 7760 -3060 7780
rect -3040 7760 -3020 7780
rect -3000 7760 -2990 7780
rect -3165 7754 -2990 7760
rect -3155 7750 -2990 7754
rect -3155 7704 -2990 7710
rect -5680 7672 -5665 7704
rect -3165 7700 -2990 7704
rect -3165 7680 -3145 7700
rect -3120 7680 -3100 7700
rect -3080 7680 -3060 7700
rect -3040 7680 -3020 7700
rect -3000 7680 -2990 7700
rect -3165 7672 -2990 7680
rect -3155 7670 -2990 7672
rect -3155 7622 -2990 7625
rect -5680 7590 -5665 7622
rect -3165 7615 -2990 7622
rect -3165 7595 -3145 7615
rect -3120 7595 -3100 7615
rect -3080 7595 -3060 7615
rect -3040 7595 -3020 7615
rect -3000 7595 -2990 7615
rect -3165 7590 -2990 7595
rect -3155 7585 -2990 7590
rect -3155 7540 -2990 7545
rect -5680 7508 -5665 7540
rect -3165 7535 -2990 7540
rect -3165 7515 -3145 7535
rect -3120 7515 -3100 7535
rect -3080 7515 -3060 7535
rect -3040 7515 -3020 7535
rect -3000 7515 -2990 7535
rect -3165 7508 -2990 7515
rect -3155 7505 -2990 7508
rect -3155 7458 -2990 7460
rect -5680 7426 -5665 7458
rect -3165 7450 -2990 7458
rect -3165 7430 -3145 7450
rect -3120 7430 -3100 7450
rect -3080 7430 -3060 7450
rect -3040 7430 -3020 7450
rect -3000 7430 -2990 7450
rect -3165 7426 -2990 7430
rect -3155 7420 -2990 7426
rect -3155 7376 -2990 7380
rect -5680 7344 -5665 7376
rect -3165 7370 -2990 7376
rect -3165 7350 -3145 7370
rect -3120 7350 -3100 7370
rect -3080 7350 -3060 7370
rect -3040 7350 -3020 7370
rect -3000 7350 -2990 7370
rect -3165 7344 -2990 7350
rect -3155 7340 -2990 7344
rect -3155 7294 -2990 7300
rect -5680 7262 -5665 7294
rect -3165 7290 -2990 7294
rect -3165 7270 -3145 7290
rect -3120 7270 -3100 7290
rect -3080 7270 -3060 7290
rect -3040 7270 -3020 7290
rect -3000 7270 -2990 7290
rect -3165 7262 -2990 7270
rect -3155 7260 -2990 7262
rect -3155 7212 -2990 7215
rect -5680 7180 -5665 7212
rect -3165 7205 -2990 7212
rect -3165 7185 -3145 7205
rect -3120 7185 -3100 7205
rect -3080 7185 -3060 7205
rect -3040 7185 -3020 7205
rect -3000 7185 -2990 7205
rect -3165 7180 -2990 7185
rect -3155 7175 -2990 7180
rect -3155 7130 -2990 7135
rect -5680 7098 -5665 7130
rect -3165 7125 -2990 7130
rect -3165 7105 -3145 7125
rect -3120 7105 -3100 7125
rect -3080 7105 -3060 7125
rect -3040 7105 -3020 7125
rect -3000 7105 -2990 7125
rect -3165 7098 -2990 7105
rect -3155 7095 -2990 7098
rect -3155 7048 -2990 7050
rect -5680 7016 -5665 7048
rect -3165 7040 -2990 7048
rect -3165 7020 -3145 7040
rect -3120 7020 -3100 7040
rect -3080 7020 -3060 7040
rect -3040 7020 -3020 7040
rect -3000 7020 -2990 7040
rect -3165 7016 -2990 7020
rect -3155 7010 -2990 7016
rect -3155 6966 -2990 6970
rect -5680 6934 -5665 6966
rect -3165 6960 -2990 6966
rect -3165 6940 -3145 6960
rect -3120 6940 -3100 6960
rect -3080 6940 -3060 6960
rect -3040 6940 -3020 6960
rect -3000 6940 -2990 6960
rect -3165 6934 -2990 6940
rect -3155 6930 -2990 6934
rect -3155 6884 -2990 6890
rect -5680 6852 -5665 6884
rect -3165 6880 -2990 6884
rect -3165 6860 -3145 6880
rect -3120 6860 -3100 6880
rect -3080 6860 -3060 6880
rect -3040 6860 -3020 6880
rect -3000 6860 -2990 6880
rect -3165 6852 -2990 6860
rect -3155 6850 -2990 6852
rect -3155 6802 -2990 6805
rect -5680 6770 -5665 6802
rect -3165 6795 -2990 6802
rect -3165 6775 -3145 6795
rect -3120 6775 -3100 6795
rect -3080 6775 -3060 6795
rect -3040 6775 -3020 6795
rect -3000 6775 -2990 6795
rect -3165 6770 -2990 6775
rect -3155 6765 -2990 6770
rect -3155 6720 -2990 6725
rect -5680 6688 -5665 6720
rect -3165 6715 -2990 6720
rect -3165 6695 -3145 6715
rect -3120 6695 -3100 6715
rect -3080 6695 -3060 6715
rect -3040 6695 -3020 6715
rect -3000 6695 -2990 6715
rect -3165 6688 -2990 6695
rect -3155 6685 -2990 6688
rect -3155 6638 -2990 6645
rect -5680 6606 -5665 6638
rect -3165 6635 -2990 6638
rect -3165 6615 -3145 6635
rect -3120 6615 -3100 6635
rect -3080 6615 -3060 6635
rect -3040 6615 -3020 6635
rect -3000 6615 -2990 6635
rect -3165 6606 -2990 6615
rect -3155 6605 -2990 6606
rect -3155 6556 -2990 6560
rect -5680 6524 -5665 6556
rect -3165 6550 -2990 6556
rect -3165 6530 -3145 6550
rect -3120 6530 -3100 6550
rect -3080 6530 -3060 6550
rect -3040 6530 -3020 6550
rect -3000 6530 -2990 6550
rect -3165 6524 -2990 6530
rect -3155 6520 -2990 6524
rect -3155 6474 -2990 6480
rect -5680 6442 -5665 6474
rect -3165 6470 -2990 6474
rect -3165 6450 -3145 6470
rect -3120 6450 -3100 6470
rect -3080 6450 -3060 6470
rect -3040 6450 -3020 6470
rect -3000 6450 -2990 6470
rect -3165 6442 -2990 6450
rect -3155 6440 -2990 6442
rect -3155 6392 -2990 6400
rect -5680 6360 -5665 6392
rect -3165 6390 -2990 6392
rect -3165 6370 -3145 6390
rect -3120 6370 -3100 6390
rect -3080 6370 -3060 6390
rect -3040 6370 -3020 6390
rect -3000 6370 -2990 6390
rect -3165 6360 -2990 6370
rect -2150 8442 -1985 8445
rect -2150 8435 -1975 8442
rect -2150 8415 -2140 8435
rect -2120 8415 -2100 8435
rect -2080 8415 -2060 8435
rect -2040 8415 -2020 8435
rect -1995 8415 -1975 8435
rect -2150 8410 -1975 8415
rect 525 8410 540 8442
rect -2150 8405 -1985 8410
rect -2150 8360 -1985 8365
rect -2150 8355 -1975 8360
rect -2150 8335 -2140 8355
rect -2120 8335 -2100 8355
rect -2080 8335 -2060 8355
rect -2040 8335 -2020 8355
rect -1995 8335 -1975 8355
rect -2150 8328 -1975 8335
rect 525 8328 540 8360
rect -2150 8325 -1985 8328
rect -2150 8278 -1985 8280
rect -2150 8270 -1975 8278
rect -2150 8250 -2140 8270
rect -2120 8250 -2100 8270
rect -2080 8250 -2060 8270
rect -2040 8250 -2020 8270
rect -1995 8250 -1975 8270
rect -2150 8246 -1975 8250
rect 525 8246 540 8278
rect -2150 8240 -1985 8246
rect -2150 8196 -1985 8200
rect -2150 8190 -1975 8196
rect -2150 8170 -2140 8190
rect -2120 8170 -2100 8190
rect -2080 8170 -2060 8190
rect -2040 8170 -2020 8190
rect -1995 8170 -1975 8190
rect -2150 8164 -1975 8170
rect 525 8164 540 8196
rect -2150 8160 -1985 8164
rect -2150 8114 -1985 8120
rect -2150 8110 -1975 8114
rect -2150 8090 -2140 8110
rect -2120 8090 -2100 8110
rect -2080 8090 -2060 8110
rect -2040 8090 -2020 8110
rect -1995 8090 -1975 8110
rect -2150 8082 -1975 8090
rect 525 8082 540 8114
rect -2150 8080 -1985 8082
rect -2150 8032 -1985 8035
rect -2150 8025 -1975 8032
rect -2150 8005 -2140 8025
rect -2120 8005 -2100 8025
rect -2080 8005 -2060 8025
rect -2040 8005 -2020 8025
rect -1995 8005 -1975 8025
rect -2150 8000 -1975 8005
rect 525 8000 540 8032
rect -2150 7995 -1985 8000
rect -2150 7950 -1985 7955
rect -2150 7945 -1975 7950
rect -2150 7925 -2140 7945
rect -2120 7925 -2100 7945
rect -2080 7925 -2060 7945
rect -2040 7925 -2020 7945
rect -1995 7925 -1975 7945
rect -2150 7918 -1975 7925
rect 525 7918 540 7950
rect -2150 7915 -1985 7918
rect -2150 7868 -1985 7870
rect -2150 7860 -1975 7868
rect -2150 7840 -2140 7860
rect -2120 7840 -2100 7860
rect -2080 7840 -2060 7860
rect -2040 7840 -2020 7860
rect -1995 7840 -1975 7860
rect -2150 7836 -1975 7840
rect 525 7836 540 7868
rect -2150 7830 -1985 7836
rect -2150 7786 -1985 7790
rect -2150 7780 -1975 7786
rect -2150 7760 -2140 7780
rect -2120 7760 -2100 7780
rect -2080 7760 -2060 7780
rect -2040 7760 -2020 7780
rect -1995 7760 -1975 7780
rect -2150 7754 -1975 7760
rect 525 7754 540 7786
rect -2150 7750 -1985 7754
rect -2150 7704 -1985 7710
rect -2150 7700 -1975 7704
rect -2150 7680 -2140 7700
rect -2120 7680 -2100 7700
rect -2080 7680 -2060 7700
rect -2040 7680 -2020 7700
rect -1995 7680 -1975 7700
rect -2150 7672 -1975 7680
rect 525 7672 540 7704
rect -2150 7670 -1985 7672
rect -2150 7622 -1985 7625
rect -2150 7615 -1975 7622
rect -2150 7595 -2140 7615
rect -2120 7595 -2100 7615
rect -2080 7595 -2060 7615
rect -2040 7595 -2020 7615
rect -1995 7595 -1975 7615
rect -2150 7590 -1975 7595
rect 525 7590 540 7622
rect -2150 7585 -1985 7590
rect -2150 7540 -1985 7545
rect -2150 7535 -1975 7540
rect -2150 7515 -2140 7535
rect -2120 7515 -2100 7535
rect -2080 7515 -2060 7535
rect -2040 7515 -2020 7535
rect -1995 7515 -1975 7535
rect -2150 7508 -1975 7515
rect 525 7508 540 7540
rect -2150 7505 -1985 7508
rect -2150 7458 -1985 7460
rect -2150 7450 -1975 7458
rect -2150 7430 -2140 7450
rect -2120 7430 -2100 7450
rect -2080 7430 -2060 7450
rect -2040 7430 -2020 7450
rect -1995 7430 -1975 7450
rect -2150 7426 -1975 7430
rect 525 7426 540 7458
rect -2150 7420 -1985 7426
rect -2150 7376 -1985 7380
rect -2150 7370 -1975 7376
rect -2150 7350 -2140 7370
rect -2120 7350 -2100 7370
rect -2080 7350 -2060 7370
rect -2040 7350 -2020 7370
rect -1995 7350 -1975 7370
rect -2150 7344 -1975 7350
rect 525 7344 540 7376
rect -2150 7340 -1985 7344
rect -2150 7294 -1985 7300
rect -2150 7290 -1975 7294
rect -2150 7270 -2140 7290
rect -2120 7270 -2100 7290
rect -2080 7270 -2060 7290
rect -2040 7270 -2020 7290
rect -1995 7270 -1975 7290
rect -2150 7262 -1975 7270
rect 525 7262 540 7294
rect -2150 7260 -1985 7262
rect -2150 7212 -1985 7215
rect -2150 7205 -1975 7212
rect -2150 7185 -2140 7205
rect -2120 7185 -2100 7205
rect -2080 7185 -2060 7205
rect -2040 7185 -2020 7205
rect -1995 7185 -1975 7205
rect -2150 7180 -1975 7185
rect 525 7180 540 7212
rect -2150 7175 -1985 7180
rect -2150 7130 -1985 7135
rect -2150 7125 -1975 7130
rect -2150 7105 -2140 7125
rect -2120 7105 -2100 7125
rect -2080 7105 -2060 7125
rect -2040 7105 -2020 7125
rect -1995 7105 -1975 7125
rect -2150 7098 -1975 7105
rect 525 7098 540 7130
rect -2150 7095 -1985 7098
rect -2150 7048 -1985 7050
rect -2150 7040 -1975 7048
rect -2150 7020 -2140 7040
rect -2120 7020 -2100 7040
rect -2080 7020 -2060 7040
rect -2040 7020 -2020 7040
rect -1995 7020 -1975 7040
rect -2150 7016 -1975 7020
rect 525 7016 540 7048
rect -2150 7010 -1985 7016
rect -2150 6966 -1985 6970
rect -2150 6960 -1975 6966
rect -2150 6940 -2140 6960
rect -2120 6940 -2100 6960
rect -2080 6940 -2060 6960
rect -2040 6940 -2020 6960
rect -1995 6940 -1975 6960
rect -2150 6934 -1975 6940
rect 525 6934 540 6966
rect -2150 6930 -1985 6934
rect -2150 6884 -1985 6890
rect -2150 6880 -1975 6884
rect -2150 6860 -2140 6880
rect -2120 6860 -2100 6880
rect -2080 6860 -2060 6880
rect -2040 6860 -2020 6880
rect -1995 6860 -1975 6880
rect -2150 6852 -1975 6860
rect 525 6852 540 6884
rect -2150 6850 -1985 6852
rect -2150 6802 -1985 6805
rect -2150 6795 -1975 6802
rect -2150 6775 -2140 6795
rect -2120 6775 -2100 6795
rect -2080 6775 -2060 6795
rect -2040 6775 -2020 6795
rect -1995 6775 -1975 6795
rect -2150 6770 -1975 6775
rect 525 6770 540 6802
rect -2150 6765 -1985 6770
rect -2150 6720 -1985 6725
rect -2150 6715 -1975 6720
rect -2150 6695 -2140 6715
rect -2120 6695 -2100 6715
rect -2080 6695 -2060 6715
rect -2040 6695 -2020 6715
rect -1995 6695 -1975 6715
rect -2150 6688 -1975 6695
rect 525 6688 540 6720
rect -2150 6685 -1985 6688
rect -2150 6638 -1985 6645
rect -2150 6635 -1975 6638
rect -2150 6615 -2140 6635
rect -2120 6615 -2100 6635
rect -2080 6615 -2060 6635
rect -2040 6615 -2020 6635
rect -1995 6615 -1975 6635
rect -2150 6606 -1975 6615
rect 525 6606 540 6638
rect -2150 6605 -1985 6606
rect -2150 6556 -1985 6560
rect -2150 6550 -1975 6556
rect -2150 6530 -2140 6550
rect -2120 6530 -2100 6550
rect -2080 6530 -2060 6550
rect -2040 6530 -2020 6550
rect -1995 6530 -1975 6550
rect -2150 6524 -1975 6530
rect 525 6524 540 6556
rect -2150 6520 -1985 6524
rect -2150 6474 -1985 6480
rect -2150 6470 -1975 6474
rect -2150 6450 -2140 6470
rect -2120 6450 -2100 6470
rect -2080 6450 -2060 6470
rect -2040 6450 -2020 6470
rect -1995 6450 -1975 6470
rect -2150 6442 -1975 6450
rect 525 6442 540 6474
rect -2150 6440 -1985 6442
rect -2150 6392 -1985 6400
rect -2150 6390 -1975 6392
rect -2150 6370 -2140 6390
rect -2120 6370 -2100 6390
rect -2080 6370 -2060 6390
rect -2040 6370 -2020 6390
rect -1995 6370 -1975 6390
rect -2150 6360 -1975 6370
rect 525 6360 540 6392
rect -5610 5965 -5595 6010
rect -3095 6000 -2920 6010
rect -3095 5975 -3075 6000
rect -3050 5975 -3030 6000
rect -3010 5975 -2990 6000
rect -2970 5975 -2950 6000
rect -2930 5975 -2920 6000
rect -3095 5965 -2920 5975
rect -2220 6000 -2045 6010
rect -2220 5975 -2210 6000
rect -2190 5975 -2170 6000
rect -2150 5975 -2130 6000
rect -2110 5975 -2090 6000
rect -2065 5975 -2045 6000
rect -2220 5965 -2045 5975
rect 455 5965 470 6010
rect -5610 5870 -5595 5915
rect -3095 5905 -2920 5915
rect -3095 5880 -3075 5905
rect -3050 5880 -3030 5905
rect -3010 5880 -2990 5905
rect -2970 5880 -2950 5905
rect -2930 5880 -2920 5905
rect -3095 5870 -2920 5880
rect -2220 5905 -2045 5915
rect -2220 5880 -2210 5905
rect -2190 5880 -2170 5905
rect -2150 5880 -2130 5905
rect -2110 5880 -2090 5905
rect -2065 5880 -2045 5905
rect -2220 5870 -2045 5880
rect 455 5870 470 5915
rect -5610 5775 -5595 5820
rect -3095 5810 -2920 5820
rect -3095 5785 -3075 5810
rect -3050 5785 -3030 5810
rect -3010 5785 -2990 5810
rect -2970 5785 -2950 5810
rect -2930 5785 -2920 5810
rect -3095 5775 -2920 5785
rect -2220 5810 -2045 5820
rect -2220 5785 -2210 5810
rect -2190 5785 -2170 5810
rect -2150 5785 -2130 5810
rect -2110 5785 -2090 5810
rect -2065 5785 -2045 5810
rect -2220 5775 -2045 5785
rect 455 5775 470 5820
rect -5610 5680 -5595 5725
rect -3095 5715 -2920 5725
rect -3095 5690 -3075 5715
rect -3050 5690 -3030 5715
rect -3010 5690 -2990 5715
rect -2970 5690 -2950 5715
rect -2930 5690 -2920 5715
rect -3095 5680 -2920 5690
rect -2220 5715 -2045 5725
rect -2220 5690 -2210 5715
rect -2190 5690 -2170 5715
rect -2150 5690 -2130 5715
rect -2110 5690 -2090 5715
rect -2065 5690 -2045 5715
rect -2220 5680 -2045 5690
rect 455 5680 470 5725
rect -5610 5585 -5595 5630
rect -3095 5620 -2920 5630
rect -3095 5595 -3075 5620
rect -3050 5595 -3030 5620
rect -3010 5595 -2990 5620
rect -2970 5595 -2950 5620
rect -2930 5595 -2920 5620
rect -3095 5585 -2920 5595
rect -2220 5620 -2045 5630
rect -2220 5595 -2210 5620
rect -2190 5595 -2170 5620
rect -2150 5595 -2130 5620
rect -2110 5595 -2090 5620
rect -2065 5595 -2045 5620
rect -2220 5585 -2045 5595
rect 455 5585 470 5630
rect -5610 5490 -5595 5535
rect -3095 5525 -2920 5535
rect -3095 5500 -3075 5525
rect -3050 5500 -3030 5525
rect -3010 5500 -2990 5525
rect -2970 5500 -2950 5525
rect -2930 5500 -2920 5525
rect -3095 5490 -2920 5500
rect -2220 5525 -2045 5535
rect -2220 5500 -2210 5525
rect -2190 5500 -2170 5525
rect -2150 5500 -2130 5525
rect -2110 5500 -2090 5525
rect -2065 5500 -2045 5525
rect -2220 5490 -2045 5500
rect 455 5490 470 5535
rect -5610 5395 -5595 5440
rect -3095 5430 -2920 5440
rect -3095 5405 -3075 5430
rect -3050 5405 -3030 5430
rect -3010 5405 -2990 5430
rect -2970 5405 -2950 5430
rect -2930 5405 -2920 5430
rect -3095 5395 -2920 5405
rect -2220 5430 -2045 5440
rect -2220 5405 -2210 5430
rect -2190 5405 -2170 5430
rect -2150 5405 -2130 5430
rect -2110 5405 -2090 5430
rect -2065 5405 -2045 5430
rect -2220 5395 -2045 5405
rect 455 5395 470 5440
rect -5610 5300 -5595 5345
rect -3095 5335 -2920 5345
rect -3095 5310 -3075 5335
rect -3050 5310 -3030 5335
rect -3010 5310 -2990 5335
rect -2970 5310 -2950 5335
rect -2930 5310 -2920 5335
rect -3095 5300 -2920 5310
rect -2220 5335 -2045 5345
rect -2220 5310 -2210 5335
rect -2190 5310 -2170 5335
rect -2150 5310 -2130 5335
rect -2110 5310 -2090 5335
rect -2065 5310 -2045 5335
rect -2220 5300 -2045 5310
rect 455 5300 470 5345
rect -5610 5205 -5595 5250
rect -3095 5240 -2920 5250
rect -3095 5215 -3075 5240
rect -3050 5215 -3030 5240
rect -3010 5215 -2990 5240
rect -2970 5215 -2950 5240
rect -2930 5215 -2920 5240
rect -3095 5205 -2920 5215
rect -2220 5240 -2045 5250
rect -2220 5215 -2210 5240
rect -2190 5215 -2170 5240
rect -2150 5215 -2130 5240
rect -2110 5215 -2090 5240
rect -2065 5215 -2045 5240
rect -2220 5205 -2045 5215
rect 455 5205 470 5250
rect -5610 5110 -5595 5155
rect -3095 5145 -2920 5155
rect -3095 5120 -3075 5145
rect -3050 5120 -3030 5145
rect -3010 5120 -2990 5145
rect -2970 5120 -2950 5145
rect -2930 5120 -2920 5145
rect -3095 5110 -2920 5120
rect -2220 5145 -2045 5155
rect -2220 5120 -2210 5145
rect -2190 5120 -2170 5145
rect -2150 5120 -2130 5145
rect -2110 5120 -2090 5145
rect -2065 5120 -2045 5145
rect -2220 5110 -2045 5120
rect 455 5110 470 5155
rect -5610 5015 -5595 5060
rect -3095 5050 -2920 5060
rect -3095 5025 -3075 5050
rect -3050 5025 -3030 5050
rect -3010 5025 -2990 5050
rect -2970 5025 -2950 5050
rect -2930 5025 -2920 5050
rect -3095 5015 -2920 5025
rect -2220 5050 -2045 5060
rect -2220 5025 -2210 5050
rect -2190 5025 -2170 5050
rect -2150 5025 -2130 5050
rect -2110 5025 -2090 5050
rect -2065 5025 -2045 5050
rect -2220 5015 -2045 5025
rect 455 5015 470 5060
rect -5610 4920 -5595 4965
rect -3095 4955 -2920 4965
rect -3095 4930 -3075 4955
rect -3050 4930 -3030 4955
rect -3010 4930 -2990 4955
rect -2970 4930 -2950 4955
rect -2930 4930 -2920 4955
rect -3095 4920 -2920 4930
rect -2220 4955 -2045 4965
rect -2220 4930 -2210 4955
rect -2190 4930 -2170 4955
rect -2150 4930 -2130 4955
rect -2110 4930 -2090 4955
rect -2065 4930 -2045 4955
rect -2220 4920 -2045 4930
rect 455 4920 470 4965
rect -5610 4825 -5595 4870
rect -3095 4860 -2920 4870
rect -3095 4835 -3075 4860
rect -3050 4835 -3030 4860
rect -3010 4835 -2990 4860
rect -2970 4835 -2950 4860
rect -2930 4835 -2920 4860
rect -3095 4825 -2920 4835
rect -2220 4860 -2045 4870
rect -2220 4835 -2210 4860
rect -2190 4835 -2170 4860
rect -2150 4835 -2130 4860
rect -2110 4835 -2090 4860
rect -2065 4835 -2045 4860
rect -2220 4825 -2045 4835
rect 455 4825 470 4870
rect -5610 4730 -5595 4775
rect -3095 4765 -2920 4775
rect -3095 4740 -3075 4765
rect -3050 4740 -3030 4765
rect -3010 4740 -2990 4765
rect -2970 4740 -2950 4765
rect -2930 4740 -2920 4765
rect -3095 4730 -2920 4740
rect -2220 4765 -2045 4775
rect -2220 4740 -2210 4765
rect -2190 4740 -2170 4765
rect -2150 4740 -2130 4765
rect -2110 4740 -2090 4765
rect -2065 4740 -2045 4765
rect -2220 4730 -2045 4740
rect 455 4730 470 4775
rect -5610 4635 -5595 4680
rect -3095 4670 -2920 4680
rect -3095 4645 -3075 4670
rect -3050 4645 -3030 4670
rect -3010 4645 -2990 4670
rect -2970 4645 -2950 4670
rect -2930 4645 -2920 4670
rect -3095 4635 -2920 4645
rect -2220 4670 -2045 4680
rect -2220 4645 -2210 4670
rect -2190 4645 -2170 4670
rect -2150 4645 -2130 4670
rect -2110 4645 -2090 4670
rect -2065 4645 -2045 4670
rect -2220 4635 -2045 4645
rect 455 4635 470 4680
rect -5610 4540 -5595 4585
rect -3095 4575 -2920 4585
rect -3095 4550 -3075 4575
rect -3050 4550 -3030 4575
rect -3010 4550 -2990 4575
rect -2970 4550 -2950 4575
rect -2930 4550 -2920 4575
rect -3095 4540 -2920 4550
rect -2220 4575 -2045 4585
rect -2220 4550 -2210 4575
rect -2190 4550 -2170 4575
rect -2150 4550 -2130 4575
rect -2110 4550 -2090 4575
rect -2065 4550 -2045 4575
rect -2220 4540 -2045 4550
rect 455 4540 470 4585
rect -5610 4445 -5595 4490
rect -3095 4480 -2920 4490
rect -3095 4455 -3075 4480
rect -3050 4455 -3030 4480
rect -3010 4455 -2990 4480
rect -2970 4455 -2950 4480
rect -2930 4455 -2920 4480
rect -3095 4445 -2920 4455
rect -2220 4480 -2045 4490
rect -2220 4455 -2210 4480
rect -2190 4455 -2170 4480
rect -2150 4455 -2130 4480
rect -2110 4455 -2090 4480
rect -2065 4455 -2045 4480
rect -2220 4445 -2045 4455
rect 455 4445 470 4490
rect -5610 4350 -5595 4395
rect -3095 4385 -2920 4395
rect -3095 4360 -3075 4385
rect -3050 4360 -3030 4385
rect -3010 4360 -2990 4385
rect -2970 4360 -2950 4385
rect -2930 4360 -2920 4385
rect -3095 4350 -2920 4360
rect -2220 4385 -2045 4395
rect -2220 4360 -2210 4385
rect -2190 4360 -2170 4385
rect -2150 4360 -2130 4385
rect -2110 4360 -2090 4385
rect -2065 4360 -2045 4385
rect -2220 4350 -2045 4360
rect 455 4350 470 4395
rect -5610 4255 -5595 4300
rect -3095 4290 -2920 4300
rect -3095 4265 -3075 4290
rect -3050 4265 -3030 4290
rect -3010 4265 -2990 4290
rect -2970 4265 -2950 4290
rect -2930 4265 -2920 4290
rect -3095 4255 -2920 4265
rect -2220 4290 -2045 4300
rect -2220 4265 -2210 4290
rect -2190 4265 -2170 4290
rect -2150 4265 -2130 4290
rect -2110 4265 -2090 4290
rect -2065 4265 -2045 4290
rect -2220 4255 -2045 4265
rect 455 4255 470 4300
rect -5610 4160 -5595 4205
rect -3095 4195 -2920 4205
rect -3095 4170 -3075 4195
rect -3050 4170 -3030 4195
rect -3010 4170 -2990 4195
rect -2970 4170 -2950 4195
rect -2930 4170 -2920 4195
rect -3095 4160 -2920 4170
rect -2220 4195 -2045 4205
rect -2220 4170 -2210 4195
rect -2190 4170 -2170 4195
rect -2150 4170 -2130 4195
rect -2110 4170 -2090 4195
rect -2065 4170 -2045 4195
rect -2220 4160 -2045 4170
rect 455 4160 470 4205
rect -5610 4065 -5595 4110
rect -3095 4100 -2920 4110
rect -3095 4075 -3075 4100
rect -3050 4075 -3030 4100
rect -3010 4075 -2990 4100
rect -2970 4075 -2950 4100
rect -2930 4075 -2920 4100
rect -3095 4065 -2920 4075
rect -2220 4100 -2045 4110
rect -2220 4075 -2210 4100
rect -2190 4075 -2170 4100
rect -2150 4075 -2130 4100
rect -2110 4075 -2090 4100
rect -2065 4075 -2045 4100
rect -2220 4065 -2045 4075
rect 455 4065 470 4110
rect -5610 3970 -5595 4015
rect -3095 4005 -2920 4015
rect -3095 3980 -3075 4005
rect -3050 3980 -3030 4005
rect -3010 3980 -2990 4005
rect -2970 3980 -2950 4005
rect -2930 3980 -2920 4005
rect -3095 3970 -2920 3980
rect -2220 4005 -2045 4015
rect -2220 3980 -2210 4005
rect -2190 3980 -2170 4005
rect -2150 3980 -2130 4005
rect -2110 3980 -2090 4005
rect -2065 3980 -2045 4005
rect -2220 3970 -2045 3980
rect 455 3970 470 4015
rect -5610 3875 -5595 3920
rect -3095 3910 -2920 3920
rect -3095 3885 -3075 3910
rect -3050 3885 -3030 3910
rect -3010 3885 -2990 3910
rect -2970 3885 -2950 3910
rect -2930 3885 -2920 3910
rect -3095 3875 -2920 3885
rect -2220 3910 -2045 3920
rect -2220 3885 -2210 3910
rect -2190 3885 -2170 3910
rect -2150 3885 -2130 3910
rect -2110 3885 -2090 3910
rect -2065 3885 -2045 3910
rect -2220 3875 -2045 3885
rect 455 3875 470 3920
rect -5610 3780 -5595 3825
rect -3095 3815 -2920 3825
rect -3095 3790 -3075 3815
rect -3050 3790 -3030 3815
rect -3010 3790 -2990 3815
rect -2970 3790 -2950 3815
rect -2930 3790 -2920 3815
rect -3095 3780 -2920 3790
rect -2220 3815 -2045 3825
rect -2220 3790 -2210 3815
rect -2190 3790 -2170 3815
rect -2150 3790 -2130 3815
rect -2110 3790 -2090 3815
rect -2065 3790 -2045 3815
rect -2220 3780 -2045 3790
rect 455 3780 470 3825
rect -5610 3685 -5595 3730
rect -3095 3720 -2920 3730
rect -3095 3695 -3075 3720
rect -3050 3695 -3030 3720
rect -3010 3695 -2990 3720
rect -2970 3695 -2950 3720
rect -2930 3695 -2920 3720
rect -3095 3685 -2920 3695
rect -2220 3720 -2045 3730
rect -2220 3695 -2210 3720
rect -2190 3695 -2170 3720
rect -2150 3695 -2130 3720
rect -2110 3695 -2090 3720
rect -2065 3695 -2045 3720
rect -2220 3685 -2045 3695
rect 455 3685 470 3730
rect -5610 3590 -5595 3635
rect -3095 3625 -2920 3635
rect -3095 3600 -3075 3625
rect -3050 3600 -3030 3625
rect -3010 3600 -2990 3625
rect -2970 3600 -2950 3625
rect -2930 3600 -2920 3625
rect -3095 3590 -2920 3600
rect -2220 3625 -2045 3635
rect -2220 3600 -2210 3625
rect -2190 3600 -2170 3625
rect -2150 3600 -2130 3625
rect -2110 3600 -2090 3625
rect -2065 3600 -2045 3625
rect -2220 3590 -2045 3600
rect 455 3590 470 3635
<< polycont >>
rect -3145 8415 -3120 8435
rect -3100 8415 -3080 8435
rect -3060 8415 -3040 8435
rect -3020 8415 -3000 8435
rect -3145 8335 -3120 8355
rect -3100 8335 -3080 8355
rect -3060 8335 -3040 8355
rect -3020 8335 -3000 8355
rect -3145 8250 -3120 8270
rect -3100 8250 -3080 8270
rect -3060 8250 -3040 8270
rect -3020 8250 -3000 8270
rect -3145 8170 -3120 8190
rect -3100 8170 -3080 8190
rect -3060 8170 -3040 8190
rect -3020 8170 -3000 8190
rect -3145 8090 -3120 8110
rect -3100 8090 -3080 8110
rect -3060 8090 -3040 8110
rect -3020 8090 -3000 8110
rect -3145 8005 -3120 8025
rect -3100 8005 -3080 8025
rect -3060 8005 -3040 8025
rect -3020 8005 -3000 8025
rect -3145 7925 -3120 7945
rect -3100 7925 -3080 7945
rect -3060 7925 -3040 7945
rect -3020 7925 -3000 7945
rect -3145 7840 -3120 7860
rect -3100 7840 -3080 7860
rect -3060 7840 -3040 7860
rect -3020 7840 -3000 7860
rect -3145 7760 -3120 7780
rect -3100 7760 -3080 7780
rect -3060 7760 -3040 7780
rect -3020 7760 -3000 7780
rect -3145 7680 -3120 7700
rect -3100 7680 -3080 7700
rect -3060 7680 -3040 7700
rect -3020 7680 -3000 7700
rect -3145 7595 -3120 7615
rect -3100 7595 -3080 7615
rect -3060 7595 -3040 7615
rect -3020 7595 -3000 7615
rect -3145 7515 -3120 7535
rect -3100 7515 -3080 7535
rect -3060 7515 -3040 7535
rect -3020 7515 -3000 7535
rect -3145 7430 -3120 7450
rect -3100 7430 -3080 7450
rect -3060 7430 -3040 7450
rect -3020 7430 -3000 7450
rect -3145 7350 -3120 7370
rect -3100 7350 -3080 7370
rect -3060 7350 -3040 7370
rect -3020 7350 -3000 7370
rect -3145 7270 -3120 7290
rect -3100 7270 -3080 7290
rect -3060 7270 -3040 7290
rect -3020 7270 -3000 7290
rect -3145 7185 -3120 7205
rect -3100 7185 -3080 7205
rect -3060 7185 -3040 7205
rect -3020 7185 -3000 7205
rect -3145 7105 -3120 7125
rect -3100 7105 -3080 7125
rect -3060 7105 -3040 7125
rect -3020 7105 -3000 7125
rect -3145 7020 -3120 7040
rect -3100 7020 -3080 7040
rect -3060 7020 -3040 7040
rect -3020 7020 -3000 7040
rect -3145 6940 -3120 6960
rect -3100 6940 -3080 6960
rect -3060 6940 -3040 6960
rect -3020 6940 -3000 6960
rect -3145 6860 -3120 6880
rect -3100 6860 -3080 6880
rect -3060 6860 -3040 6880
rect -3020 6860 -3000 6880
rect -3145 6775 -3120 6795
rect -3100 6775 -3080 6795
rect -3060 6775 -3040 6795
rect -3020 6775 -3000 6795
rect -3145 6695 -3120 6715
rect -3100 6695 -3080 6715
rect -3060 6695 -3040 6715
rect -3020 6695 -3000 6715
rect -3145 6615 -3120 6635
rect -3100 6615 -3080 6635
rect -3060 6615 -3040 6635
rect -3020 6615 -3000 6635
rect -3145 6530 -3120 6550
rect -3100 6530 -3080 6550
rect -3060 6530 -3040 6550
rect -3020 6530 -3000 6550
rect -3145 6450 -3120 6470
rect -3100 6450 -3080 6470
rect -3060 6450 -3040 6470
rect -3020 6450 -3000 6470
rect -3145 6370 -3120 6390
rect -3100 6370 -3080 6390
rect -3060 6370 -3040 6390
rect -3020 6370 -3000 6390
rect -2140 8415 -2120 8435
rect -2100 8415 -2080 8435
rect -2060 8415 -2040 8435
rect -2020 8415 -1995 8435
rect -2140 8335 -2120 8355
rect -2100 8335 -2080 8355
rect -2060 8335 -2040 8355
rect -2020 8335 -1995 8355
rect -2140 8250 -2120 8270
rect -2100 8250 -2080 8270
rect -2060 8250 -2040 8270
rect -2020 8250 -1995 8270
rect -2140 8170 -2120 8190
rect -2100 8170 -2080 8190
rect -2060 8170 -2040 8190
rect -2020 8170 -1995 8190
rect -2140 8090 -2120 8110
rect -2100 8090 -2080 8110
rect -2060 8090 -2040 8110
rect -2020 8090 -1995 8110
rect -2140 8005 -2120 8025
rect -2100 8005 -2080 8025
rect -2060 8005 -2040 8025
rect -2020 8005 -1995 8025
rect -2140 7925 -2120 7945
rect -2100 7925 -2080 7945
rect -2060 7925 -2040 7945
rect -2020 7925 -1995 7945
rect -2140 7840 -2120 7860
rect -2100 7840 -2080 7860
rect -2060 7840 -2040 7860
rect -2020 7840 -1995 7860
rect -2140 7760 -2120 7780
rect -2100 7760 -2080 7780
rect -2060 7760 -2040 7780
rect -2020 7760 -1995 7780
rect -2140 7680 -2120 7700
rect -2100 7680 -2080 7700
rect -2060 7680 -2040 7700
rect -2020 7680 -1995 7700
rect -2140 7595 -2120 7615
rect -2100 7595 -2080 7615
rect -2060 7595 -2040 7615
rect -2020 7595 -1995 7615
rect -2140 7515 -2120 7535
rect -2100 7515 -2080 7535
rect -2060 7515 -2040 7535
rect -2020 7515 -1995 7535
rect -2140 7430 -2120 7450
rect -2100 7430 -2080 7450
rect -2060 7430 -2040 7450
rect -2020 7430 -1995 7450
rect -2140 7350 -2120 7370
rect -2100 7350 -2080 7370
rect -2060 7350 -2040 7370
rect -2020 7350 -1995 7370
rect -2140 7270 -2120 7290
rect -2100 7270 -2080 7290
rect -2060 7270 -2040 7290
rect -2020 7270 -1995 7290
rect -2140 7185 -2120 7205
rect -2100 7185 -2080 7205
rect -2060 7185 -2040 7205
rect -2020 7185 -1995 7205
rect -2140 7105 -2120 7125
rect -2100 7105 -2080 7125
rect -2060 7105 -2040 7125
rect -2020 7105 -1995 7125
rect -2140 7020 -2120 7040
rect -2100 7020 -2080 7040
rect -2060 7020 -2040 7040
rect -2020 7020 -1995 7040
rect -2140 6940 -2120 6960
rect -2100 6940 -2080 6960
rect -2060 6940 -2040 6960
rect -2020 6940 -1995 6960
rect -2140 6860 -2120 6880
rect -2100 6860 -2080 6880
rect -2060 6860 -2040 6880
rect -2020 6860 -1995 6880
rect -2140 6775 -2120 6795
rect -2100 6775 -2080 6795
rect -2060 6775 -2040 6795
rect -2020 6775 -1995 6795
rect -2140 6695 -2120 6715
rect -2100 6695 -2080 6715
rect -2060 6695 -2040 6715
rect -2020 6695 -1995 6715
rect -2140 6615 -2120 6635
rect -2100 6615 -2080 6635
rect -2060 6615 -2040 6635
rect -2020 6615 -1995 6635
rect -2140 6530 -2120 6550
rect -2100 6530 -2080 6550
rect -2060 6530 -2040 6550
rect -2020 6530 -1995 6550
rect -2140 6450 -2120 6470
rect -2100 6450 -2080 6470
rect -2060 6450 -2040 6470
rect -2020 6450 -1995 6470
rect -2140 6370 -2120 6390
rect -2100 6370 -2080 6390
rect -2060 6370 -2040 6390
rect -2020 6370 -1995 6390
rect -3075 5975 -3050 6000
rect -3030 5975 -3010 6000
rect -2990 5975 -2970 6000
rect -2950 5975 -2930 6000
rect -2210 5975 -2190 6000
rect -2170 5975 -2150 6000
rect -2130 5975 -2110 6000
rect -2090 5975 -2065 6000
rect -3075 5880 -3050 5905
rect -3030 5880 -3010 5905
rect -2990 5880 -2970 5905
rect -2950 5880 -2930 5905
rect -2210 5880 -2190 5905
rect -2170 5880 -2150 5905
rect -2130 5880 -2110 5905
rect -2090 5880 -2065 5905
rect -3075 5785 -3050 5810
rect -3030 5785 -3010 5810
rect -2990 5785 -2970 5810
rect -2950 5785 -2930 5810
rect -2210 5785 -2190 5810
rect -2170 5785 -2150 5810
rect -2130 5785 -2110 5810
rect -2090 5785 -2065 5810
rect -3075 5690 -3050 5715
rect -3030 5690 -3010 5715
rect -2990 5690 -2970 5715
rect -2950 5690 -2930 5715
rect -2210 5690 -2190 5715
rect -2170 5690 -2150 5715
rect -2130 5690 -2110 5715
rect -2090 5690 -2065 5715
rect -3075 5595 -3050 5620
rect -3030 5595 -3010 5620
rect -2990 5595 -2970 5620
rect -2950 5595 -2930 5620
rect -2210 5595 -2190 5620
rect -2170 5595 -2150 5620
rect -2130 5595 -2110 5620
rect -2090 5595 -2065 5620
rect -3075 5500 -3050 5525
rect -3030 5500 -3010 5525
rect -2990 5500 -2970 5525
rect -2950 5500 -2930 5525
rect -2210 5500 -2190 5525
rect -2170 5500 -2150 5525
rect -2130 5500 -2110 5525
rect -2090 5500 -2065 5525
rect -3075 5405 -3050 5430
rect -3030 5405 -3010 5430
rect -2990 5405 -2970 5430
rect -2950 5405 -2930 5430
rect -2210 5405 -2190 5430
rect -2170 5405 -2150 5430
rect -2130 5405 -2110 5430
rect -2090 5405 -2065 5430
rect -3075 5310 -3050 5335
rect -3030 5310 -3010 5335
rect -2990 5310 -2970 5335
rect -2950 5310 -2930 5335
rect -2210 5310 -2190 5335
rect -2170 5310 -2150 5335
rect -2130 5310 -2110 5335
rect -2090 5310 -2065 5335
rect -3075 5215 -3050 5240
rect -3030 5215 -3010 5240
rect -2990 5215 -2970 5240
rect -2950 5215 -2930 5240
rect -2210 5215 -2190 5240
rect -2170 5215 -2150 5240
rect -2130 5215 -2110 5240
rect -2090 5215 -2065 5240
rect -3075 5120 -3050 5145
rect -3030 5120 -3010 5145
rect -2990 5120 -2970 5145
rect -2950 5120 -2930 5145
rect -2210 5120 -2190 5145
rect -2170 5120 -2150 5145
rect -2130 5120 -2110 5145
rect -2090 5120 -2065 5145
rect -3075 5025 -3050 5050
rect -3030 5025 -3010 5050
rect -2990 5025 -2970 5050
rect -2950 5025 -2930 5050
rect -2210 5025 -2190 5050
rect -2170 5025 -2150 5050
rect -2130 5025 -2110 5050
rect -2090 5025 -2065 5050
rect -3075 4930 -3050 4955
rect -3030 4930 -3010 4955
rect -2990 4930 -2970 4955
rect -2950 4930 -2930 4955
rect -2210 4930 -2190 4955
rect -2170 4930 -2150 4955
rect -2130 4930 -2110 4955
rect -2090 4930 -2065 4955
rect -3075 4835 -3050 4860
rect -3030 4835 -3010 4860
rect -2990 4835 -2970 4860
rect -2950 4835 -2930 4860
rect -2210 4835 -2190 4860
rect -2170 4835 -2150 4860
rect -2130 4835 -2110 4860
rect -2090 4835 -2065 4860
rect -3075 4740 -3050 4765
rect -3030 4740 -3010 4765
rect -2990 4740 -2970 4765
rect -2950 4740 -2930 4765
rect -2210 4740 -2190 4765
rect -2170 4740 -2150 4765
rect -2130 4740 -2110 4765
rect -2090 4740 -2065 4765
rect -3075 4645 -3050 4670
rect -3030 4645 -3010 4670
rect -2990 4645 -2970 4670
rect -2950 4645 -2930 4670
rect -2210 4645 -2190 4670
rect -2170 4645 -2150 4670
rect -2130 4645 -2110 4670
rect -2090 4645 -2065 4670
rect -3075 4550 -3050 4575
rect -3030 4550 -3010 4575
rect -2990 4550 -2970 4575
rect -2950 4550 -2930 4575
rect -2210 4550 -2190 4575
rect -2170 4550 -2150 4575
rect -2130 4550 -2110 4575
rect -2090 4550 -2065 4575
rect -3075 4455 -3050 4480
rect -3030 4455 -3010 4480
rect -2990 4455 -2970 4480
rect -2950 4455 -2930 4480
rect -2210 4455 -2190 4480
rect -2170 4455 -2150 4480
rect -2130 4455 -2110 4480
rect -2090 4455 -2065 4480
rect -3075 4360 -3050 4385
rect -3030 4360 -3010 4385
rect -2990 4360 -2970 4385
rect -2950 4360 -2930 4385
rect -2210 4360 -2190 4385
rect -2170 4360 -2150 4385
rect -2130 4360 -2110 4385
rect -2090 4360 -2065 4385
rect -3075 4265 -3050 4290
rect -3030 4265 -3010 4290
rect -2990 4265 -2970 4290
rect -2950 4265 -2930 4290
rect -2210 4265 -2190 4290
rect -2170 4265 -2150 4290
rect -2130 4265 -2110 4290
rect -2090 4265 -2065 4290
rect -3075 4170 -3050 4195
rect -3030 4170 -3010 4195
rect -2990 4170 -2970 4195
rect -2950 4170 -2930 4195
rect -2210 4170 -2190 4195
rect -2170 4170 -2150 4195
rect -2130 4170 -2110 4195
rect -2090 4170 -2065 4195
rect -3075 4075 -3050 4100
rect -3030 4075 -3010 4100
rect -2990 4075 -2970 4100
rect -2950 4075 -2930 4100
rect -2210 4075 -2190 4100
rect -2170 4075 -2150 4100
rect -2130 4075 -2110 4100
rect -2090 4075 -2065 4100
rect -3075 3980 -3050 4005
rect -3030 3980 -3010 4005
rect -2990 3980 -2970 4005
rect -2950 3980 -2930 4005
rect -2210 3980 -2190 4005
rect -2170 3980 -2150 4005
rect -2130 3980 -2110 4005
rect -2090 3980 -2065 4005
rect -3075 3885 -3050 3910
rect -3030 3885 -3010 3910
rect -2990 3885 -2970 3910
rect -2950 3885 -2930 3910
rect -2210 3885 -2190 3910
rect -2170 3885 -2150 3910
rect -2130 3885 -2110 3910
rect -2090 3885 -2065 3910
rect -3075 3790 -3050 3815
rect -3030 3790 -3010 3815
rect -2990 3790 -2970 3815
rect -2950 3790 -2930 3815
rect -2210 3790 -2190 3815
rect -2170 3790 -2150 3815
rect -2130 3790 -2110 3815
rect -2090 3790 -2065 3815
rect -3075 3695 -3050 3720
rect -3030 3695 -3010 3720
rect -2990 3695 -2970 3720
rect -2950 3695 -2930 3720
rect -2210 3695 -2190 3720
rect -2170 3695 -2150 3720
rect -2130 3695 -2110 3720
rect -2090 3695 -2065 3720
rect -3075 3600 -3050 3625
rect -3030 3600 -3010 3625
rect -2990 3600 -2970 3625
rect -2950 3600 -2930 3625
rect -2210 3600 -2190 3625
rect -2170 3600 -2150 3625
rect -2130 3600 -2110 3625
rect -2090 3600 -2065 3625
<< locali >>
rect -5775 8605 -2915 8620
rect -5775 8585 -5710 8605
rect -5690 8585 -5670 8605
rect -5650 8585 -5630 8605
rect -5610 8585 -5590 8605
rect -5570 8585 -5550 8605
rect -5530 8585 -5510 8605
rect -5490 8585 -5470 8605
rect -5450 8585 -5430 8605
rect -5410 8585 -5390 8605
rect -5370 8585 -5350 8605
rect -5330 8585 -5310 8605
rect -5290 8585 -5270 8605
rect -5250 8585 -5230 8605
rect -5210 8585 -5190 8605
rect -5170 8585 -5150 8605
rect -5130 8585 -5110 8605
rect -5090 8585 -5070 8605
rect -5050 8585 -5030 8605
rect -5010 8585 -4990 8605
rect -4970 8585 -4950 8605
rect -4930 8585 -4910 8605
rect -4890 8585 -4870 8605
rect -4850 8585 -4830 8605
rect -4810 8585 -4790 8605
rect -4770 8585 -4750 8605
rect -4730 8585 -4710 8605
rect -4690 8585 -4670 8605
rect -4650 8585 -4630 8605
rect -4610 8585 -4590 8605
rect -4570 8585 -4550 8605
rect -4530 8585 -4510 8605
rect -4490 8585 -4470 8605
rect -4450 8585 -4430 8605
rect -4410 8585 -4390 8605
rect -4370 8585 -4350 8605
rect -4330 8585 -4310 8605
rect -4290 8585 -4270 8605
rect -4250 8585 -4230 8605
rect -4210 8585 -4190 8605
rect -4170 8585 -4150 8605
rect -4130 8585 -4110 8605
rect -4090 8585 -4070 8605
rect -4050 8585 -4030 8605
rect -4010 8585 -3990 8605
rect -3970 8585 -3950 8605
rect -3930 8585 -3910 8605
rect -3890 8585 -3870 8605
rect -3850 8585 -3830 8605
rect -3810 8585 -3790 8605
rect -3770 8585 -3750 8605
rect -3730 8585 -3710 8605
rect -3690 8585 -3670 8605
rect -3650 8585 -3630 8605
rect -3610 8585 -3590 8605
rect -3570 8585 -3550 8605
rect -3530 8585 -3510 8605
rect -3490 8585 -3470 8605
rect -3450 8585 -3430 8605
rect -3410 8585 -3390 8605
rect -3370 8585 -3350 8605
rect -3330 8585 -3310 8605
rect -3290 8585 -3270 8605
rect -3250 8585 -3230 8605
rect -3210 8585 -3190 8605
rect -3170 8585 -3150 8605
rect -3130 8585 -3110 8605
rect -3090 8585 -3070 8605
rect -3050 8585 -3030 8605
rect -3010 8585 -2990 8605
rect -2970 8585 -2915 8605
rect -5775 8570 -2915 8585
rect -5775 8550 -5760 8570
rect -5740 8550 -5725 8570
rect -5775 8530 -5725 8550
rect -2965 8550 -2950 8570
rect -2930 8550 -2915 8570
rect -2965 8530 -2915 8550
rect -5775 8510 -5760 8530
rect -5740 8510 -5725 8530
rect -5775 8490 -5725 8510
rect -5775 8470 -5760 8490
rect -5740 8470 -5725 8490
rect -5775 8450 -5725 8470
rect -5775 8430 -5760 8450
rect -5740 8430 -5725 8450
rect -5665 8520 -3165 8530
rect -5665 8500 -5650 8520
rect -5630 8500 -5610 8520
rect -5590 8500 -5570 8520
rect -5550 8500 -5530 8520
rect -5510 8500 -5490 8520
rect -5470 8500 -5450 8520
rect -5430 8500 -5410 8520
rect -5390 8500 -5370 8520
rect -5350 8500 -5330 8520
rect -5310 8500 -5290 8520
rect -5270 8500 -5250 8520
rect -5230 8500 -5210 8520
rect -5190 8500 -5170 8520
rect -5150 8500 -5130 8520
rect -5110 8500 -5090 8520
rect -5070 8500 -5050 8520
rect -5030 8500 -5010 8520
rect -4990 8500 -4970 8520
rect -4950 8500 -4930 8520
rect -4910 8500 -4890 8520
rect -4870 8500 -4850 8520
rect -4830 8500 -4810 8520
rect -4790 8500 -4770 8520
rect -4750 8500 -4730 8520
rect -4710 8500 -4690 8520
rect -4670 8500 -4650 8520
rect -4630 8500 -4610 8520
rect -4590 8500 -4570 8520
rect -4550 8500 -4530 8520
rect -4510 8500 -4490 8520
rect -4470 8500 -4450 8520
rect -4430 8500 -4410 8520
rect -4390 8500 -4370 8520
rect -4350 8500 -4330 8520
rect -4310 8500 -4290 8520
rect -4270 8500 -4250 8520
rect -4230 8500 -4210 8520
rect -4190 8500 -4170 8520
rect -4150 8500 -4130 8520
rect -4110 8500 -4090 8520
rect -4070 8500 -4050 8520
rect -4030 8500 -4010 8520
rect -3990 8500 -3970 8520
rect -3950 8500 -3930 8520
rect -3910 8500 -3890 8520
rect -3870 8500 -3850 8520
rect -3830 8500 -3810 8520
rect -3790 8500 -3770 8520
rect -3750 8500 -3730 8520
rect -3710 8500 -3690 8520
rect -3670 8500 -3650 8520
rect -3630 8500 -3610 8520
rect -3590 8500 -3570 8520
rect -3550 8500 -3530 8520
rect -3510 8500 -3490 8520
rect -3470 8500 -3450 8520
rect -3430 8500 -3410 8520
rect -3390 8500 -3370 8520
rect -3350 8500 -3330 8520
rect -3310 8500 -3290 8520
rect -3270 8500 -3250 8520
rect -3230 8500 -3210 8520
rect -3190 8500 -3165 8520
rect -5665 8477 -3165 8500
rect -5665 8457 -5650 8477
rect -5630 8457 -5610 8477
rect -5590 8457 -5570 8477
rect -5550 8457 -5530 8477
rect -5510 8457 -5490 8477
rect -5470 8457 -5450 8477
rect -5430 8457 -5410 8477
rect -5390 8457 -5370 8477
rect -5350 8457 -5330 8477
rect -5310 8457 -5290 8477
rect -5270 8457 -5250 8477
rect -5230 8457 -5210 8477
rect -5190 8457 -5170 8477
rect -5150 8457 -5130 8477
rect -5110 8457 -5090 8477
rect -5070 8457 -5050 8477
rect -5030 8457 -5010 8477
rect -4990 8457 -4970 8477
rect -4950 8457 -4930 8477
rect -4910 8457 -4890 8477
rect -4870 8457 -4850 8477
rect -4830 8457 -4810 8477
rect -4790 8457 -4770 8477
rect -4750 8457 -4730 8477
rect -4710 8457 -4690 8477
rect -4670 8457 -4650 8477
rect -4630 8457 -4610 8477
rect -4590 8457 -4570 8477
rect -4550 8457 -4530 8477
rect -4510 8457 -4490 8477
rect -4470 8457 -4450 8477
rect -4430 8457 -4410 8477
rect -4390 8457 -4370 8477
rect -4350 8457 -4330 8477
rect -4310 8457 -4290 8477
rect -4270 8457 -4250 8477
rect -4230 8457 -4210 8477
rect -4190 8457 -4170 8477
rect -4150 8457 -4130 8477
rect -4110 8457 -4090 8477
rect -4070 8457 -4050 8477
rect -4030 8457 -4010 8477
rect -3990 8457 -3970 8477
rect -3950 8457 -3930 8477
rect -3910 8457 -3890 8477
rect -3870 8457 -3850 8477
rect -3830 8457 -3810 8477
rect -3790 8457 -3770 8477
rect -3750 8457 -3730 8477
rect -3710 8457 -3690 8477
rect -3670 8457 -3650 8477
rect -3630 8457 -3610 8477
rect -3590 8457 -3570 8477
rect -3550 8457 -3530 8477
rect -3510 8457 -3490 8477
rect -3470 8457 -3450 8477
rect -3430 8457 -3410 8477
rect -3390 8457 -3370 8477
rect -3350 8457 -3330 8477
rect -3310 8457 -3290 8477
rect -3270 8457 -3250 8477
rect -3230 8457 -3210 8477
rect -3190 8457 -3165 8477
rect -5665 8447 -3165 8457
rect -2965 8510 -2950 8530
rect -2930 8510 -2915 8530
rect -2965 8490 -2915 8510
rect -2965 8470 -2950 8490
rect -2930 8470 -2915 8490
rect -2965 8450 -2915 8470
rect -5775 8410 -5725 8430
rect -5775 8390 -5760 8410
rect -5740 8390 -5725 8410
rect -3145 8435 -2990 8445
rect -3120 8415 -3100 8435
rect -3080 8415 -3060 8435
rect -3040 8415 -3020 8435
rect -3000 8415 -2990 8435
rect -3145 8405 -2990 8415
rect -2965 8430 -2950 8450
rect -2930 8430 -2915 8450
rect -2965 8410 -2915 8430
rect -5775 8370 -5725 8390
rect -5775 8350 -5760 8370
rect -5740 8350 -5725 8370
rect -5665 8395 -3165 8405
rect -5665 8375 -5650 8395
rect -5630 8375 -5610 8395
rect -5590 8375 -5570 8395
rect -5550 8375 -5530 8395
rect -5510 8375 -5490 8395
rect -5470 8375 -5450 8395
rect -5430 8375 -5410 8395
rect -5390 8375 -5370 8395
rect -5350 8375 -5330 8395
rect -5310 8375 -5290 8395
rect -5270 8375 -5250 8395
rect -5230 8375 -5210 8395
rect -5190 8375 -5170 8395
rect -5150 8375 -5130 8395
rect -5110 8375 -5090 8395
rect -5070 8375 -5050 8395
rect -5030 8375 -5010 8395
rect -4990 8375 -4970 8395
rect -4950 8375 -4930 8395
rect -4910 8375 -4890 8395
rect -4870 8375 -4850 8395
rect -4830 8375 -4810 8395
rect -4790 8375 -4770 8395
rect -4750 8375 -4730 8395
rect -4710 8375 -4690 8395
rect -4670 8375 -4650 8395
rect -4630 8375 -4610 8395
rect -4590 8375 -4570 8395
rect -4550 8375 -4530 8395
rect -4510 8375 -4490 8395
rect -4470 8375 -4450 8395
rect -4430 8375 -4410 8395
rect -4390 8375 -4370 8395
rect -4350 8375 -4330 8395
rect -4310 8375 -4290 8395
rect -4270 8375 -4250 8395
rect -4230 8375 -4210 8395
rect -4190 8375 -4170 8395
rect -4150 8375 -4130 8395
rect -4110 8375 -4090 8395
rect -4070 8375 -4050 8395
rect -4030 8375 -4010 8395
rect -3990 8375 -3970 8395
rect -3950 8375 -3930 8395
rect -3910 8375 -3890 8395
rect -3870 8375 -3850 8395
rect -3830 8375 -3810 8395
rect -3790 8375 -3770 8395
rect -3750 8375 -3730 8395
rect -3710 8375 -3690 8395
rect -3670 8375 -3650 8395
rect -3630 8375 -3610 8395
rect -3590 8375 -3570 8395
rect -3550 8375 -3530 8395
rect -3510 8375 -3490 8395
rect -3470 8375 -3450 8395
rect -3430 8375 -3410 8395
rect -3390 8375 -3370 8395
rect -3350 8375 -3330 8395
rect -3310 8375 -3290 8395
rect -3270 8375 -3250 8395
rect -3230 8375 -3210 8395
rect -3190 8375 -3165 8395
rect -5665 8365 -3165 8375
rect -2965 8390 -2950 8410
rect -2930 8390 -2915 8410
rect -2965 8370 -2915 8390
rect -5775 8330 -5725 8350
rect -5775 8310 -5760 8330
rect -5740 8310 -5725 8330
rect -3145 8355 -2990 8365
rect -3120 8335 -3100 8355
rect -3080 8335 -3060 8355
rect -3040 8335 -3020 8355
rect -3000 8335 -2990 8355
rect -3145 8325 -2990 8335
rect -2965 8350 -2950 8370
rect -2930 8350 -2915 8370
rect -2965 8330 -2915 8350
rect -5775 8290 -5725 8310
rect -5775 8270 -5760 8290
rect -5740 8270 -5725 8290
rect -5665 8313 -3165 8323
rect -5665 8293 -5650 8313
rect -5630 8293 -5610 8313
rect -5590 8293 -5570 8313
rect -5550 8293 -5530 8313
rect -5510 8293 -5490 8313
rect -5470 8293 -5450 8313
rect -5430 8293 -5410 8313
rect -5390 8293 -5370 8313
rect -5350 8293 -5330 8313
rect -5310 8293 -5290 8313
rect -5270 8293 -5250 8313
rect -5230 8293 -5210 8313
rect -5190 8293 -5170 8313
rect -5150 8293 -5130 8313
rect -5110 8293 -5090 8313
rect -5070 8293 -5050 8313
rect -5030 8293 -5010 8313
rect -4990 8293 -4970 8313
rect -4950 8293 -4930 8313
rect -4910 8293 -4890 8313
rect -4870 8293 -4850 8313
rect -4830 8293 -4810 8313
rect -4790 8293 -4770 8313
rect -4750 8293 -4730 8313
rect -4710 8293 -4690 8313
rect -4670 8293 -4650 8313
rect -4630 8293 -4610 8313
rect -4590 8293 -4570 8313
rect -4550 8293 -4530 8313
rect -4510 8293 -4490 8313
rect -4470 8293 -4450 8313
rect -4430 8293 -4410 8313
rect -4390 8293 -4370 8313
rect -4350 8293 -4330 8313
rect -4310 8293 -4290 8313
rect -4270 8293 -4250 8313
rect -4230 8293 -4210 8313
rect -4190 8293 -4170 8313
rect -4150 8293 -4130 8313
rect -4110 8293 -4090 8313
rect -4070 8293 -4050 8313
rect -4030 8293 -4010 8313
rect -3990 8293 -3970 8313
rect -3950 8293 -3930 8313
rect -3910 8293 -3890 8313
rect -3870 8293 -3850 8313
rect -3830 8293 -3810 8313
rect -3790 8293 -3770 8313
rect -3750 8293 -3730 8313
rect -3710 8293 -3690 8313
rect -3670 8293 -3650 8313
rect -3630 8293 -3610 8313
rect -3590 8293 -3570 8313
rect -3550 8293 -3530 8313
rect -3510 8293 -3490 8313
rect -3470 8293 -3450 8313
rect -3430 8293 -3410 8313
rect -3390 8293 -3370 8313
rect -3350 8293 -3330 8313
rect -3310 8293 -3290 8313
rect -3270 8293 -3250 8313
rect -3230 8293 -3210 8313
rect -3190 8293 -3165 8313
rect -5665 8283 -3165 8293
rect -2965 8310 -2950 8330
rect -2930 8310 -2915 8330
rect -2965 8290 -2915 8310
rect -5775 8250 -5725 8270
rect -5775 8230 -5760 8250
rect -5740 8230 -5725 8250
rect -3145 8270 -2990 8280
rect -3120 8250 -3100 8270
rect -3080 8250 -3060 8270
rect -3040 8250 -3020 8270
rect -3000 8250 -2990 8270
rect -5775 8210 -5725 8230
rect -5775 8190 -5760 8210
rect -5740 8190 -5725 8210
rect -5665 8231 -3165 8241
rect -3145 8240 -2990 8250
rect -2965 8270 -2950 8290
rect -2930 8270 -2915 8290
rect -2965 8250 -2915 8270
rect -5665 8211 -5650 8231
rect -5630 8211 -5610 8231
rect -5590 8211 -5570 8231
rect -5550 8211 -5530 8231
rect -5510 8211 -5490 8231
rect -5470 8211 -5450 8231
rect -5430 8211 -5410 8231
rect -5390 8211 -5370 8231
rect -5350 8211 -5330 8231
rect -5310 8211 -5290 8231
rect -5270 8211 -5250 8231
rect -5230 8211 -5210 8231
rect -5190 8211 -5170 8231
rect -5150 8211 -5130 8231
rect -5110 8211 -5090 8231
rect -5070 8211 -5050 8231
rect -5030 8211 -5010 8231
rect -4990 8211 -4970 8231
rect -4950 8211 -4930 8231
rect -4910 8211 -4890 8231
rect -4870 8211 -4850 8231
rect -4830 8211 -4810 8231
rect -4790 8211 -4770 8231
rect -4750 8211 -4730 8231
rect -4710 8211 -4690 8231
rect -4670 8211 -4650 8231
rect -4630 8211 -4610 8231
rect -4590 8211 -4570 8231
rect -4550 8211 -4530 8231
rect -4510 8211 -4490 8231
rect -4470 8211 -4450 8231
rect -4430 8211 -4410 8231
rect -4390 8211 -4370 8231
rect -4350 8211 -4330 8231
rect -4310 8211 -4290 8231
rect -4270 8211 -4250 8231
rect -4230 8211 -4210 8231
rect -4190 8211 -4170 8231
rect -4150 8211 -4130 8231
rect -4110 8211 -4090 8231
rect -4070 8211 -4050 8231
rect -4030 8211 -4010 8231
rect -3990 8211 -3970 8231
rect -3950 8211 -3930 8231
rect -3910 8211 -3890 8231
rect -3870 8211 -3850 8231
rect -3830 8211 -3810 8231
rect -3790 8211 -3770 8231
rect -3750 8211 -3730 8231
rect -3710 8211 -3690 8231
rect -3670 8211 -3650 8231
rect -3630 8211 -3610 8231
rect -3590 8211 -3570 8231
rect -3550 8211 -3530 8231
rect -3510 8211 -3490 8231
rect -3470 8211 -3450 8231
rect -3430 8211 -3410 8231
rect -3390 8211 -3370 8231
rect -3350 8211 -3330 8231
rect -3310 8211 -3290 8231
rect -3270 8211 -3250 8231
rect -3230 8211 -3210 8231
rect -3190 8211 -3165 8231
rect -5665 8201 -3165 8211
rect -2965 8230 -2950 8250
rect -2930 8230 -2915 8250
rect -2965 8210 -2915 8230
rect -5775 8170 -5725 8190
rect -5775 8150 -5760 8170
rect -5740 8150 -5725 8170
rect -3145 8190 -2990 8200
rect -3120 8170 -3100 8190
rect -3080 8170 -3060 8190
rect -3040 8170 -3020 8190
rect -3000 8170 -2990 8190
rect -3145 8160 -2990 8170
rect -2965 8190 -2950 8210
rect -2930 8190 -2915 8210
rect -2965 8170 -2915 8190
rect -5775 8130 -5725 8150
rect -5775 8110 -5760 8130
rect -5740 8110 -5725 8130
rect -5665 8149 -3165 8159
rect -5665 8129 -5650 8149
rect -5630 8129 -5610 8149
rect -5590 8129 -5570 8149
rect -5550 8129 -5530 8149
rect -5510 8129 -5490 8149
rect -5470 8129 -5450 8149
rect -5430 8129 -5410 8149
rect -5390 8129 -5370 8149
rect -5350 8129 -5330 8149
rect -5310 8129 -5290 8149
rect -5270 8129 -5250 8149
rect -5230 8129 -5210 8149
rect -5190 8129 -5170 8149
rect -5150 8129 -5130 8149
rect -5110 8129 -5090 8149
rect -5070 8129 -5050 8149
rect -5030 8129 -5010 8149
rect -4990 8129 -4970 8149
rect -4950 8129 -4930 8149
rect -4910 8129 -4890 8149
rect -4870 8129 -4850 8149
rect -4830 8129 -4810 8149
rect -4790 8129 -4770 8149
rect -4750 8129 -4730 8149
rect -4710 8129 -4690 8149
rect -4670 8129 -4650 8149
rect -4630 8129 -4610 8149
rect -4590 8129 -4570 8149
rect -4550 8129 -4530 8149
rect -4510 8129 -4490 8149
rect -4470 8129 -4450 8149
rect -4430 8129 -4410 8149
rect -4390 8129 -4370 8149
rect -4350 8129 -4330 8149
rect -4310 8129 -4290 8149
rect -4270 8129 -4250 8149
rect -4230 8129 -4210 8149
rect -4190 8129 -4170 8149
rect -4150 8129 -4130 8149
rect -4110 8129 -4090 8149
rect -4070 8129 -4050 8149
rect -4030 8129 -4010 8149
rect -3990 8129 -3970 8149
rect -3950 8129 -3930 8149
rect -3910 8129 -3890 8149
rect -3870 8129 -3850 8149
rect -3830 8129 -3810 8149
rect -3790 8129 -3770 8149
rect -3750 8129 -3730 8149
rect -3710 8129 -3690 8149
rect -3670 8129 -3650 8149
rect -3630 8129 -3610 8149
rect -3590 8129 -3570 8149
rect -3550 8129 -3530 8149
rect -3510 8129 -3490 8149
rect -3470 8129 -3450 8149
rect -3430 8129 -3410 8149
rect -3390 8129 -3370 8149
rect -3350 8129 -3330 8149
rect -3310 8129 -3290 8149
rect -3270 8129 -3250 8149
rect -3230 8129 -3210 8149
rect -3190 8129 -3165 8149
rect -5665 8119 -3165 8129
rect -2965 8150 -2950 8170
rect -2930 8150 -2915 8170
rect -2965 8130 -2915 8150
rect -5775 8090 -5725 8110
rect -5775 8070 -5760 8090
rect -5740 8070 -5725 8090
rect -3145 8110 -2990 8120
rect -3120 8090 -3100 8110
rect -3080 8090 -3060 8110
rect -3040 8090 -3020 8110
rect -3000 8090 -2990 8110
rect -3145 8080 -2990 8090
rect -2965 8110 -2950 8130
rect -2930 8110 -2915 8130
rect -2965 8090 -2915 8110
rect -5775 8050 -5725 8070
rect -5775 8030 -5760 8050
rect -5740 8030 -5725 8050
rect -5665 8067 -3165 8077
rect -5665 8047 -5650 8067
rect -5630 8047 -5610 8067
rect -5590 8047 -5570 8067
rect -5550 8047 -5530 8067
rect -5510 8047 -5490 8067
rect -5470 8047 -5450 8067
rect -5430 8047 -5410 8067
rect -5390 8047 -5370 8067
rect -5350 8047 -5330 8067
rect -5310 8047 -5290 8067
rect -5270 8047 -5250 8067
rect -5230 8047 -5210 8067
rect -5190 8047 -5170 8067
rect -5150 8047 -5130 8067
rect -5110 8047 -5090 8067
rect -5070 8047 -5050 8067
rect -5030 8047 -5010 8067
rect -4990 8047 -4970 8067
rect -4950 8047 -4930 8067
rect -4910 8047 -4890 8067
rect -4870 8047 -4850 8067
rect -4830 8047 -4810 8067
rect -4790 8047 -4770 8067
rect -4750 8047 -4730 8067
rect -4710 8047 -4690 8067
rect -4670 8047 -4650 8067
rect -4630 8047 -4610 8067
rect -4590 8047 -4570 8067
rect -4550 8047 -4530 8067
rect -4510 8047 -4490 8067
rect -4470 8047 -4450 8067
rect -4430 8047 -4410 8067
rect -4390 8047 -4370 8067
rect -4350 8047 -4330 8067
rect -4310 8047 -4290 8067
rect -4270 8047 -4250 8067
rect -4230 8047 -4210 8067
rect -4190 8047 -4170 8067
rect -4150 8047 -4130 8067
rect -4110 8047 -4090 8067
rect -4070 8047 -4050 8067
rect -4030 8047 -4010 8067
rect -3990 8047 -3970 8067
rect -3950 8047 -3930 8067
rect -3910 8047 -3890 8067
rect -3870 8047 -3850 8067
rect -3830 8047 -3810 8067
rect -3790 8047 -3770 8067
rect -3750 8047 -3730 8067
rect -3710 8047 -3690 8067
rect -3670 8047 -3650 8067
rect -3630 8047 -3610 8067
rect -3590 8047 -3570 8067
rect -3550 8047 -3530 8067
rect -3510 8047 -3490 8067
rect -3470 8047 -3450 8067
rect -3430 8047 -3410 8067
rect -3390 8047 -3370 8067
rect -3350 8047 -3330 8067
rect -3310 8047 -3290 8067
rect -3270 8047 -3250 8067
rect -3230 8047 -3210 8067
rect -3190 8047 -3165 8067
rect -5665 8037 -3165 8047
rect -2965 8070 -2950 8090
rect -2930 8070 -2915 8090
rect -2965 8050 -2915 8070
rect -5775 8010 -5725 8030
rect -5775 7990 -5760 8010
rect -5740 7990 -5725 8010
rect -3145 8025 -2990 8035
rect -3120 8005 -3100 8025
rect -3080 8005 -3060 8025
rect -3040 8005 -3020 8025
rect -3000 8005 -2990 8025
rect -3145 7995 -2990 8005
rect -2965 8030 -2950 8050
rect -2930 8030 -2915 8050
rect -2965 8010 -2915 8030
rect -5775 7970 -5725 7990
rect -5775 7950 -5760 7970
rect -5740 7950 -5725 7970
rect -5665 7985 -3165 7995
rect -5665 7965 -5650 7985
rect -5630 7965 -5610 7985
rect -5590 7965 -5570 7985
rect -5550 7965 -5530 7985
rect -5510 7965 -5490 7985
rect -5470 7965 -5450 7985
rect -5430 7965 -5410 7985
rect -5390 7965 -5370 7985
rect -5350 7965 -5330 7985
rect -5310 7965 -5290 7985
rect -5270 7965 -5250 7985
rect -5230 7965 -5210 7985
rect -5190 7965 -5170 7985
rect -5150 7965 -5130 7985
rect -5110 7965 -5090 7985
rect -5070 7965 -5050 7985
rect -5030 7965 -5010 7985
rect -4990 7965 -4970 7985
rect -4950 7965 -4930 7985
rect -4910 7965 -4890 7985
rect -4870 7965 -4850 7985
rect -4830 7965 -4810 7985
rect -4790 7965 -4770 7985
rect -4750 7965 -4730 7985
rect -4710 7965 -4690 7985
rect -4670 7965 -4650 7985
rect -4630 7965 -4610 7985
rect -4590 7965 -4570 7985
rect -4550 7965 -4530 7985
rect -4510 7965 -4490 7985
rect -4470 7965 -4450 7985
rect -4430 7965 -4410 7985
rect -4390 7965 -4370 7985
rect -4350 7965 -4330 7985
rect -4310 7965 -4290 7985
rect -4270 7965 -4250 7985
rect -4230 7965 -4210 7985
rect -4190 7965 -4170 7985
rect -4150 7965 -4130 7985
rect -4110 7965 -4090 7985
rect -4070 7965 -4050 7985
rect -4030 7965 -4010 7985
rect -3990 7965 -3970 7985
rect -3950 7965 -3930 7985
rect -3910 7965 -3890 7985
rect -3870 7965 -3850 7985
rect -3830 7965 -3810 7985
rect -3790 7965 -3770 7985
rect -3750 7965 -3730 7985
rect -3710 7965 -3690 7985
rect -3670 7965 -3650 7985
rect -3630 7965 -3610 7985
rect -3590 7965 -3570 7985
rect -3550 7965 -3530 7985
rect -3510 7965 -3490 7985
rect -3470 7965 -3450 7985
rect -3430 7965 -3410 7985
rect -3390 7965 -3370 7985
rect -3350 7965 -3330 7985
rect -3310 7965 -3290 7985
rect -3270 7965 -3250 7985
rect -3230 7965 -3210 7985
rect -3190 7965 -3165 7985
rect -5665 7955 -3165 7965
rect -2965 7990 -2950 8010
rect -2930 7990 -2915 8010
rect -2965 7970 -2915 7990
rect -5775 7930 -5725 7950
rect -5775 7910 -5760 7930
rect -5740 7910 -5725 7930
rect -3145 7945 -2990 7955
rect -3120 7925 -3100 7945
rect -3080 7925 -3060 7945
rect -3040 7925 -3020 7945
rect -3000 7925 -2990 7945
rect -3145 7915 -2990 7925
rect -2965 7950 -2950 7970
rect -2930 7950 -2915 7970
rect -2965 7930 -2915 7950
rect -5775 7890 -5725 7910
rect -5775 7870 -5760 7890
rect -5740 7870 -5725 7890
rect -5665 7903 -3165 7913
rect -5665 7883 -5650 7903
rect -5630 7883 -5610 7903
rect -5590 7883 -5570 7903
rect -5550 7883 -5530 7903
rect -5510 7883 -5490 7903
rect -5470 7883 -5450 7903
rect -5430 7883 -5410 7903
rect -5390 7883 -5370 7903
rect -5350 7883 -5330 7903
rect -5310 7883 -5290 7903
rect -5270 7883 -5250 7903
rect -5230 7883 -5210 7903
rect -5190 7883 -5170 7903
rect -5150 7883 -5130 7903
rect -5110 7883 -5090 7903
rect -5070 7883 -5050 7903
rect -5030 7883 -5010 7903
rect -4990 7883 -4970 7903
rect -4950 7883 -4930 7903
rect -4910 7883 -4890 7903
rect -4870 7883 -4850 7903
rect -4830 7883 -4810 7903
rect -4790 7883 -4770 7903
rect -4750 7883 -4730 7903
rect -4710 7883 -4690 7903
rect -4670 7883 -4650 7903
rect -4630 7883 -4610 7903
rect -4590 7883 -4570 7903
rect -4550 7883 -4530 7903
rect -4510 7883 -4490 7903
rect -4470 7883 -4450 7903
rect -4430 7883 -4410 7903
rect -4390 7883 -4370 7903
rect -4350 7883 -4330 7903
rect -4310 7883 -4290 7903
rect -4270 7883 -4250 7903
rect -4230 7883 -4210 7903
rect -4190 7883 -4170 7903
rect -4150 7883 -4130 7903
rect -4110 7883 -4090 7903
rect -4070 7883 -4050 7903
rect -4030 7883 -4010 7903
rect -3990 7883 -3970 7903
rect -3950 7883 -3930 7903
rect -3910 7883 -3890 7903
rect -3870 7883 -3850 7903
rect -3830 7883 -3810 7903
rect -3790 7883 -3770 7903
rect -3750 7883 -3730 7903
rect -3710 7883 -3690 7903
rect -3670 7883 -3650 7903
rect -3630 7883 -3610 7903
rect -3590 7883 -3570 7903
rect -3550 7883 -3530 7903
rect -3510 7883 -3490 7903
rect -3470 7883 -3450 7903
rect -3430 7883 -3410 7903
rect -3390 7883 -3370 7903
rect -3350 7883 -3330 7903
rect -3310 7883 -3290 7903
rect -3270 7883 -3250 7903
rect -3230 7883 -3210 7903
rect -3190 7883 -3165 7903
rect -5665 7873 -3165 7883
rect -2965 7910 -2950 7930
rect -2930 7910 -2915 7930
rect -2965 7890 -2915 7910
rect -2965 7870 -2950 7890
rect -2930 7870 -2915 7890
rect -5775 7850 -5725 7870
rect -5775 7830 -5760 7850
rect -5740 7830 -5725 7850
rect -3145 7860 -2990 7870
rect -3120 7840 -3100 7860
rect -3080 7840 -3060 7860
rect -3040 7840 -3020 7860
rect -3000 7840 -2990 7860
rect -5775 7810 -5725 7830
rect -5775 7790 -5760 7810
rect -5740 7790 -5725 7810
rect -5665 7821 -3165 7831
rect -3145 7830 -2990 7840
rect -2965 7850 -2915 7870
rect -2965 7830 -2950 7850
rect -2930 7830 -2915 7850
rect -5665 7801 -5650 7821
rect -5630 7801 -5610 7821
rect -5590 7801 -5570 7821
rect -5550 7801 -5530 7821
rect -5510 7801 -5490 7821
rect -5470 7801 -5450 7821
rect -5430 7801 -5410 7821
rect -5390 7801 -5370 7821
rect -5350 7801 -5330 7821
rect -5310 7801 -5290 7821
rect -5270 7801 -5250 7821
rect -5230 7801 -5210 7821
rect -5190 7801 -5170 7821
rect -5150 7801 -5130 7821
rect -5110 7801 -5090 7821
rect -5070 7801 -5050 7821
rect -5030 7801 -5010 7821
rect -4990 7801 -4970 7821
rect -4950 7801 -4930 7821
rect -4910 7801 -4890 7821
rect -4870 7801 -4850 7821
rect -4830 7801 -4810 7821
rect -4790 7801 -4770 7821
rect -4750 7801 -4730 7821
rect -4710 7801 -4690 7821
rect -4670 7801 -4650 7821
rect -4630 7801 -4610 7821
rect -4590 7801 -4570 7821
rect -4550 7801 -4530 7821
rect -4510 7801 -4490 7821
rect -4470 7801 -4450 7821
rect -4430 7801 -4410 7821
rect -4390 7801 -4370 7821
rect -4350 7801 -4330 7821
rect -4310 7801 -4290 7821
rect -4270 7801 -4250 7821
rect -4230 7801 -4210 7821
rect -4190 7801 -4170 7821
rect -4150 7801 -4130 7821
rect -4110 7801 -4090 7821
rect -4070 7801 -4050 7821
rect -4030 7801 -4010 7821
rect -3990 7801 -3970 7821
rect -3950 7801 -3930 7821
rect -3910 7801 -3890 7821
rect -3870 7801 -3850 7821
rect -3830 7801 -3810 7821
rect -3790 7801 -3770 7821
rect -3750 7801 -3730 7821
rect -3710 7801 -3690 7821
rect -3670 7801 -3650 7821
rect -3630 7801 -3610 7821
rect -3590 7801 -3570 7821
rect -3550 7801 -3530 7821
rect -3510 7801 -3490 7821
rect -3470 7801 -3450 7821
rect -3430 7801 -3410 7821
rect -3390 7801 -3370 7821
rect -3350 7801 -3330 7821
rect -3310 7801 -3290 7821
rect -3270 7801 -3250 7821
rect -3230 7801 -3210 7821
rect -3190 7801 -3165 7821
rect -5665 7791 -3165 7801
rect -2965 7810 -2915 7830
rect -2965 7790 -2950 7810
rect -2930 7790 -2915 7810
rect -5775 7770 -5725 7790
rect -5775 7750 -5760 7770
rect -5740 7750 -5725 7770
rect -3145 7780 -2990 7790
rect -3120 7760 -3100 7780
rect -3080 7760 -3060 7780
rect -3040 7760 -3020 7780
rect -3000 7760 -2990 7780
rect -3145 7750 -2990 7760
rect -2965 7770 -2915 7790
rect -2965 7750 -2950 7770
rect -2930 7750 -2915 7770
rect -5775 7730 -5725 7750
rect -5775 7710 -5760 7730
rect -5740 7710 -5725 7730
rect -5775 7690 -5725 7710
rect -5665 7739 -3165 7749
rect -5665 7719 -5650 7739
rect -5630 7719 -5610 7739
rect -5590 7719 -5570 7739
rect -5550 7719 -5530 7739
rect -5510 7719 -5490 7739
rect -5470 7719 -5450 7739
rect -5430 7719 -5410 7739
rect -5390 7719 -5370 7739
rect -5350 7719 -5330 7739
rect -5310 7719 -5290 7739
rect -5270 7719 -5250 7739
rect -5230 7719 -5210 7739
rect -5190 7719 -5170 7739
rect -5150 7719 -5130 7739
rect -5110 7719 -5090 7739
rect -5070 7719 -5050 7739
rect -5030 7719 -5010 7739
rect -4990 7719 -4970 7739
rect -4950 7719 -4930 7739
rect -4910 7719 -4890 7739
rect -4870 7719 -4850 7739
rect -4830 7719 -4810 7739
rect -4790 7719 -4770 7739
rect -4750 7719 -4730 7739
rect -4710 7719 -4690 7739
rect -4670 7719 -4650 7739
rect -4630 7719 -4610 7739
rect -4590 7719 -4570 7739
rect -4550 7719 -4530 7739
rect -4510 7719 -4490 7739
rect -4470 7719 -4450 7739
rect -4430 7719 -4410 7739
rect -4390 7719 -4370 7739
rect -4350 7719 -4330 7739
rect -4310 7719 -4290 7739
rect -4270 7719 -4250 7739
rect -4230 7719 -4210 7739
rect -4190 7719 -4170 7739
rect -4150 7719 -4130 7739
rect -4110 7719 -4090 7739
rect -4070 7719 -4050 7739
rect -4030 7719 -4010 7739
rect -3990 7719 -3970 7739
rect -3950 7719 -3930 7739
rect -3910 7719 -3890 7739
rect -3870 7719 -3850 7739
rect -3830 7719 -3810 7739
rect -3790 7719 -3770 7739
rect -3750 7719 -3730 7739
rect -3710 7719 -3690 7739
rect -3670 7719 -3650 7739
rect -3630 7719 -3610 7739
rect -3590 7719 -3570 7739
rect -3550 7719 -3530 7739
rect -3510 7719 -3490 7739
rect -3470 7719 -3450 7739
rect -3430 7719 -3410 7739
rect -3390 7719 -3370 7739
rect -3350 7719 -3330 7739
rect -3310 7719 -3290 7739
rect -3270 7719 -3250 7739
rect -3230 7719 -3210 7739
rect -3190 7719 -3165 7739
rect -5665 7709 -3165 7719
rect -2965 7730 -2915 7750
rect -2965 7710 -2950 7730
rect -2930 7710 -2915 7730
rect -5775 7670 -5760 7690
rect -5740 7670 -5725 7690
rect -3145 7700 -2990 7710
rect -3120 7680 -3100 7700
rect -3080 7680 -3060 7700
rect -3040 7680 -3020 7700
rect -3000 7680 -2990 7700
rect -3145 7670 -2990 7680
rect -2965 7690 -2915 7710
rect -2965 7670 -2950 7690
rect -2930 7670 -2915 7690
rect -5775 7650 -5725 7670
rect -5775 7630 -5760 7650
rect -5740 7630 -5725 7650
rect -5775 7610 -5725 7630
rect -5665 7657 -3165 7667
rect -5665 7637 -5650 7657
rect -5630 7637 -5610 7657
rect -5590 7637 -5570 7657
rect -5550 7637 -5530 7657
rect -5510 7637 -5490 7657
rect -5470 7637 -5450 7657
rect -5430 7637 -5410 7657
rect -5390 7637 -5370 7657
rect -5350 7637 -5330 7657
rect -5310 7637 -5290 7657
rect -5270 7637 -5250 7657
rect -5230 7637 -5210 7657
rect -5190 7637 -5170 7657
rect -5150 7637 -5130 7657
rect -5110 7637 -5090 7657
rect -5070 7637 -5050 7657
rect -5030 7637 -5010 7657
rect -4990 7637 -4970 7657
rect -4950 7637 -4930 7657
rect -4910 7637 -4890 7657
rect -4870 7637 -4850 7657
rect -4830 7637 -4810 7657
rect -4790 7637 -4770 7657
rect -4750 7637 -4730 7657
rect -4710 7637 -4690 7657
rect -4670 7637 -4650 7657
rect -4630 7637 -4610 7657
rect -4590 7637 -4570 7657
rect -4550 7637 -4530 7657
rect -4510 7637 -4490 7657
rect -4470 7637 -4450 7657
rect -4430 7637 -4410 7657
rect -4390 7637 -4370 7657
rect -4350 7637 -4330 7657
rect -4310 7637 -4290 7657
rect -4270 7637 -4250 7657
rect -4230 7637 -4210 7657
rect -4190 7637 -4170 7657
rect -4150 7637 -4130 7657
rect -4110 7637 -4090 7657
rect -4070 7637 -4050 7657
rect -4030 7637 -4010 7657
rect -3990 7637 -3970 7657
rect -3950 7637 -3930 7657
rect -3910 7637 -3890 7657
rect -3870 7637 -3850 7657
rect -3830 7637 -3810 7657
rect -3790 7637 -3770 7657
rect -3750 7637 -3730 7657
rect -3710 7637 -3690 7657
rect -3670 7637 -3650 7657
rect -3630 7637 -3610 7657
rect -3590 7637 -3570 7657
rect -3550 7637 -3530 7657
rect -3510 7637 -3490 7657
rect -3470 7637 -3450 7657
rect -3430 7637 -3410 7657
rect -3390 7637 -3370 7657
rect -3350 7637 -3330 7657
rect -3310 7637 -3290 7657
rect -3270 7637 -3250 7657
rect -3230 7637 -3210 7657
rect -3190 7637 -3165 7657
rect -5665 7627 -3165 7637
rect -2965 7650 -2915 7670
rect -2965 7630 -2950 7650
rect -2930 7630 -2915 7650
rect -5775 7590 -5760 7610
rect -5740 7590 -5725 7610
rect -5775 7570 -5725 7590
rect -3145 7615 -2990 7625
rect -3120 7595 -3100 7615
rect -3080 7595 -3060 7615
rect -3040 7595 -3020 7615
rect -3000 7595 -2990 7615
rect -3145 7585 -2990 7595
rect -2965 7610 -2915 7630
rect -2965 7590 -2950 7610
rect -2930 7590 -2915 7610
rect -5775 7550 -5760 7570
rect -5740 7550 -5725 7570
rect -5775 7530 -5725 7550
rect -5665 7575 -3165 7585
rect -5665 7555 -5650 7575
rect -5630 7555 -5610 7575
rect -5590 7555 -5570 7575
rect -5550 7555 -5530 7575
rect -5510 7555 -5490 7575
rect -5470 7555 -5450 7575
rect -5430 7555 -5410 7575
rect -5390 7555 -5370 7575
rect -5350 7555 -5330 7575
rect -5310 7555 -5290 7575
rect -5270 7555 -5250 7575
rect -5230 7555 -5210 7575
rect -5190 7555 -5170 7575
rect -5150 7555 -5130 7575
rect -5110 7555 -5090 7575
rect -5070 7555 -5050 7575
rect -5030 7555 -5010 7575
rect -4990 7555 -4970 7575
rect -4950 7555 -4930 7575
rect -4910 7555 -4890 7575
rect -4870 7555 -4850 7575
rect -4830 7555 -4810 7575
rect -4790 7555 -4770 7575
rect -4750 7555 -4730 7575
rect -4710 7555 -4690 7575
rect -4670 7555 -4650 7575
rect -4630 7555 -4610 7575
rect -4590 7555 -4570 7575
rect -4550 7555 -4530 7575
rect -4510 7555 -4490 7575
rect -4470 7555 -4450 7575
rect -4430 7555 -4410 7575
rect -4390 7555 -4370 7575
rect -4350 7555 -4330 7575
rect -4310 7555 -4290 7575
rect -4270 7555 -4250 7575
rect -4230 7555 -4210 7575
rect -4190 7555 -4170 7575
rect -4150 7555 -4130 7575
rect -4110 7555 -4090 7575
rect -4070 7555 -4050 7575
rect -4030 7555 -4010 7575
rect -3990 7555 -3970 7575
rect -3950 7555 -3930 7575
rect -3910 7555 -3890 7575
rect -3870 7555 -3850 7575
rect -3830 7555 -3810 7575
rect -3790 7555 -3770 7575
rect -3750 7555 -3730 7575
rect -3710 7555 -3690 7575
rect -3670 7555 -3650 7575
rect -3630 7555 -3610 7575
rect -3590 7555 -3570 7575
rect -3550 7555 -3530 7575
rect -3510 7555 -3490 7575
rect -3470 7555 -3450 7575
rect -3430 7555 -3410 7575
rect -3390 7555 -3370 7575
rect -3350 7555 -3330 7575
rect -3310 7555 -3290 7575
rect -3270 7555 -3250 7575
rect -3230 7555 -3210 7575
rect -3190 7555 -3165 7575
rect -5665 7545 -3165 7555
rect -2965 7570 -2915 7590
rect -2965 7550 -2950 7570
rect -2930 7550 -2915 7570
rect -5775 7510 -5760 7530
rect -5740 7510 -5725 7530
rect -5775 7490 -5725 7510
rect -3145 7535 -2990 7545
rect -3120 7515 -3100 7535
rect -3080 7515 -3060 7535
rect -3040 7515 -3020 7535
rect -3000 7515 -2990 7535
rect -3145 7505 -2990 7515
rect -2965 7530 -2915 7550
rect -2965 7510 -2950 7530
rect -2930 7510 -2915 7530
rect -5775 7470 -5760 7490
rect -5740 7470 -5725 7490
rect -5775 7450 -5725 7470
rect -5665 7493 -3165 7503
rect -5665 7473 -5650 7493
rect -5630 7473 -5610 7493
rect -5590 7473 -5570 7493
rect -5550 7473 -5530 7493
rect -5510 7473 -5490 7493
rect -5470 7473 -5450 7493
rect -5430 7473 -5410 7493
rect -5390 7473 -5370 7493
rect -5350 7473 -5330 7493
rect -5310 7473 -5290 7493
rect -5270 7473 -5250 7493
rect -5230 7473 -5210 7493
rect -5190 7473 -5170 7493
rect -5150 7473 -5130 7493
rect -5110 7473 -5090 7493
rect -5070 7473 -5050 7493
rect -5030 7473 -5010 7493
rect -4990 7473 -4970 7493
rect -4950 7473 -4930 7493
rect -4910 7473 -4890 7493
rect -4870 7473 -4850 7493
rect -4830 7473 -4810 7493
rect -4790 7473 -4770 7493
rect -4750 7473 -4730 7493
rect -4710 7473 -4690 7493
rect -4670 7473 -4650 7493
rect -4630 7473 -4610 7493
rect -4590 7473 -4570 7493
rect -4550 7473 -4530 7493
rect -4510 7473 -4490 7493
rect -4470 7473 -4450 7493
rect -4430 7473 -4410 7493
rect -4390 7473 -4370 7493
rect -4350 7473 -4330 7493
rect -4310 7473 -4290 7493
rect -4270 7473 -4250 7493
rect -4230 7473 -4210 7493
rect -4190 7473 -4170 7493
rect -4150 7473 -4130 7493
rect -4110 7473 -4090 7493
rect -4070 7473 -4050 7493
rect -4030 7473 -4010 7493
rect -3990 7473 -3970 7493
rect -3950 7473 -3930 7493
rect -3910 7473 -3890 7493
rect -3870 7473 -3850 7493
rect -3830 7473 -3810 7493
rect -3790 7473 -3770 7493
rect -3750 7473 -3730 7493
rect -3710 7473 -3690 7493
rect -3670 7473 -3650 7493
rect -3630 7473 -3610 7493
rect -3590 7473 -3570 7493
rect -3550 7473 -3530 7493
rect -3510 7473 -3490 7493
rect -3470 7473 -3450 7493
rect -3430 7473 -3410 7493
rect -3390 7473 -3370 7493
rect -3350 7473 -3330 7493
rect -3310 7473 -3290 7493
rect -3270 7473 -3250 7493
rect -3230 7473 -3210 7493
rect -3190 7473 -3165 7493
rect -5665 7463 -3165 7473
rect -2965 7490 -2915 7510
rect -2965 7470 -2950 7490
rect -2930 7470 -2915 7490
rect -5775 7430 -5760 7450
rect -5740 7430 -5725 7450
rect -5775 7410 -5725 7430
rect -3145 7450 -2990 7460
rect -3120 7430 -3100 7450
rect -3080 7430 -3060 7450
rect -3040 7430 -3020 7450
rect -3000 7430 -2990 7450
rect -5775 7390 -5760 7410
rect -5740 7390 -5725 7410
rect -5775 7370 -5725 7390
rect -5665 7411 -3165 7421
rect -3145 7420 -2990 7430
rect -2965 7450 -2915 7470
rect -2965 7430 -2950 7450
rect -2930 7430 -2915 7450
rect -5665 7391 -5650 7411
rect -5630 7391 -5610 7411
rect -5590 7391 -5570 7411
rect -5550 7391 -5530 7411
rect -5510 7391 -5490 7411
rect -5470 7391 -5450 7411
rect -5430 7391 -5410 7411
rect -5390 7391 -5370 7411
rect -5350 7391 -5330 7411
rect -5310 7391 -5290 7411
rect -5270 7391 -5250 7411
rect -5230 7391 -5210 7411
rect -5190 7391 -5170 7411
rect -5150 7391 -5130 7411
rect -5110 7391 -5090 7411
rect -5070 7391 -5050 7411
rect -5030 7391 -5010 7411
rect -4990 7391 -4970 7411
rect -4950 7391 -4930 7411
rect -4910 7391 -4890 7411
rect -4870 7391 -4850 7411
rect -4830 7391 -4810 7411
rect -4790 7391 -4770 7411
rect -4750 7391 -4730 7411
rect -4710 7391 -4690 7411
rect -4670 7391 -4650 7411
rect -4630 7391 -4610 7411
rect -4590 7391 -4570 7411
rect -4550 7391 -4530 7411
rect -4510 7391 -4490 7411
rect -4470 7391 -4450 7411
rect -4430 7391 -4410 7411
rect -4390 7391 -4370 7411
rect -4350 7391 -4330 7411
rect -4310 7391 -4290 7411
rect -4270 7391 -4250 7411
rect -4230 7391 -4210 7411
rect -4190 7391 -4170 7411
rect -4150 7391 -4130 7411
rect -4110 7391 -4090 7411
rect -4070 7391 -4050 7411
rect -4030 7391 -4010 7411
rect -3990 7391 -3970 7411
rect -3950 7391 -3930 7411
rect -3910 7391 -3890 7411
rect -3870 7391 -3850 7411
rect -3830 7391 -3810 7411
rect -3790 7391 -3770 7411
rect -3750 7391 -3730 7411
rect -3710 7391 -3690 7411
rect -3670 7391 -3650 7411
rect -3630 7391 -3610 7411
rect -3590 7391 -3570 7411
rect -3550 7391 -3530 7411
rect -3510 7391 -3490 7411
rect -3470 7391 -3450 7411
rect -3430 7391 -3410 7411
rect -3390 7391 -3370 7411
rect -3350 7391 -3330 7411
rect -3310 7391 -3290 7411
rect -3270 7391 -3250 7411
rect -3230 7391 -3210 7411
rect -3190 7391 -3165 7411
rect -5665 7381 -3165 7391
rect -2965 7410 -2915 7430
rect -2965 7390 -2950 7410
rect -2930 7390 -2915 7410
rect -5775 7350 -5760 7370
rect -5740 7350 -5725 7370
rect -5775 7330 -5725 7350
rect -3145 7370 -2990 7380
rect -3120 7350 -3100 7370
rect -3080 7350 -3060 7370
rect -3040 7350 -3020 7370
rect -3000 7350 -2990 7370
rect -3145 7340 -2990 7350
rect -2965 7370 -2915 7390
rect -2965 7350 -2950 7370
rect -2930 7350 -2915 7370
rect -5775 7310 -5760 7330
rect -5740 7310 -5725 7330
rect -5775 7290 -5725 7310
rect -5665 7329 -3165 7339
rect -5665 7309 -5650 7329
rect -5630 7309 -5610 7329
rect -5590 7309 -5570 7329
rect -5550 7309 -5530 7329
rect -5510 7309 -5490 7329
rect -5470 7309 -5450 7329
rect -5430 7309 -5410 7329
rect -5390 7309 -5370 7329
rect -5350 7309 -5330 7329
rect -5310 7309 -5290 7329
rect -5270 7309 -5250 7329
rect -5230 7309 -5210 7329
rect -5190 7309 -5170 7329
rect -5150 7309 -5130 7329
rect -5110 7309 -5090 7329
rect -5070 7309 -5050 7329
rect -5030 7309 -5010 7329
rect -4990 7309 -4970 7329
rect -4950 7309 -4930 7329
rect -4910 7309 -4890 7329
rect -4870 7309 -4850 7329
rect -4830 7309 -4810 7329
rect -4790 7309 -4770 7329
rect -4750 7309 -4730 7329
rect -4710 7309 -4690 7329
rect -4670 7309 -4650 7329
rect -4630 7309 -4610 7329
rect -4590 7309 -4570 7329
rect -4550 7309 -4530 7329
rect -4510 7309 -4490 7329
rect -4470 7309 -4450 7329
rect -4430 7309 -4410 7329
rect -4390 7309 -4370 7329
rect -4350 7309 -4330 7329
rect -4310 7309 -4290 7329
rect -4270 7309 -4250 7329
rect -4230 7309 -4210 7329
rect -4190 7309 -4170 7329
rect -4150 7309 -4130 7329
rect -4110 7309 -4090 7329
rect -4070 7309 -4050 7329
rect -4030 7309 -4010 7329
rect -3990 7309 -3970 7329
rect -3950 7309 -3930 7329
rect -3910 7309 -3890 7329
rect -3870 7309 -3850 7329
rect -3830 7309 -3810 7329
rect -3790 7309 -3770 7329
rect -3750 7309 -3730 7329
rect -3710 7309 -3690 7329
rect -3670 7309 -3650 7329
rect -3630 7309 -3610 7329
rect -3590 7309 -3570 7329
rect -3550 7309 -3530 7329
rect -3510 7309 -3490 7329
rect -3470 7309 -3450 7329
rect -3430 7309 -3410 7329
rect -3390 7309 -3370 7329
rect -3350 7309 -3330 7329
rect -3310 7309 -3290 7329
rect -3270 7309 -3250 7329
rect -3230 7309 -3210 7329
rect -3190 7309 -3165 7329
rect -5665 7299 -3165 7309
rect -2965 7330 -2915 7350
rect -2965 7310 -2950 7330
rect -2930 7310 -2915 7330
rect -5775 7270 -5760 7290
rect -5740 7270 -5725 7290
rect -5775 7250 -5725 7270
rect -3145 7290 -2990 7300
rect -3120 7270 -3100 7290
rect -3080 7270 -3060 7290
rect -3040 7270 -3020 7290
rect -3000 7270 -2990 7290
rect -3145 7260 -2990 7270
rect -2965 7290 -2915 7310
rect -2965 7270 -2950 7290
rect -2930 7270 -2915 7290
rect -5775 7230 -5760 7250
rect -5740 7230 -5725 7250
rect -5775 7210 -5725 7230
rect -5665 7247 -3165 7257
rect -5665 7227 -5650 7247
rect -5630 7227 -5610 7247
rect -5590 7227 -5570 7247
rect -5550 7227 -5530 7247
rect -5510 7227 -5490 7247
rect -5470 7227 -5450 7247
rect -5430 7227 -5410 7247
rect -5390 7227 -5370 7247
rect -5350 7227 -5330 7247
rect -5310 7227 -5290 7247
rect -5270 7227 -5250 7247
rect -5230 7227 -5210 7247
rect -5190 7227 -5170 7247
rect -5150 7227 -5130 7247
rect -5110 7227 -5090 7247
rect -5070 7227 -5050 7247
rect -5030 7227 -5010 7247
rect -4990 7227 -4970 7247
rect -4950 7227 -4930 7247
rect -4910 7227 -4890 7247
rect -4870 7227 -4850 7247
rect -4830 7227 -4810 7247
rect -4790 7227 -4770 7247
rect -4750 7227 -4730 7247
rect -4710 7227 -4690 7247
rect -4670 7227 -4650 7247
rect -4630 7227 -4610 7247
rect -4590 7227 -4570 7247
rect -4550 7227 -4530 7247
rect -4510 7227 -4490 7247
rect -4470 7227 -4450 7247
rect -4430 7227 -4410 7247
rect -4390 7227 -4370 7247
rect -4350 7227 -4330 7247
rect -4310 7227 -4290 7247
rect -4270 7227 -4250 7247
rect -4230 7227 -4210 7247
rect -4190 7227 -4170 7247
rect -4150 7227 -4130 7247
rect -4110 7227 -4090 7247
rect -4070 7227 -4050 7247
rect -4030 7227 -4010 7247
rect -3990 7227 -3970 7247
rect -3950 7227 -3930 7247
rect -3910 7227 -3890 7247
rect -3870 7227 -3850 7247
rect -3830 7227 -3810 7247
rect -3790 7227 -3770 7247
rect -3750 7227 -3730 7247
rect -3710 7227 -3690 7247
rect -3670 7227 -3650 7247
rect -3630 7227 -3610 7247
rect -3590 7227 -3570 7247
rect -3550 7227 -3530 7247
rect -3510 7227 -3490 7247
rect -3470 7227 -3450 7247
rect -3430 7227 -3410 7247
rect -3390 7227 -3370 7247
rect -3350 7227 -3330 7247
rect -3310 7227 -3290 7247
rect -3270 7227 -3250 7247
rect -3230 7227 -3210 7247
rect -3190 7227 -3165 7247
rect -5665 7217 -3165 7227
rect -2965 7250 -2915 7270
rect -2965 7230 -2950 7250
rect -2930 7230 -2915 7250
rect -5775 7190 -5760 7210
rect -5740 7190 -5725 7210
rect -5775 7170 -5725 7190
rect -3145 7205 -2990 7215
rect -3120 7185 -3100 7205
rect -3080 7185 -3060 7205
rect -3040 7185 -3020 7205
rect -3000 7185 -2990 7205
rect -3145 7175 -2990 7185
rect -2965 7210 -2915 7230
rect -2965 7190 -2950 7210
rect -2930 7190 -2915 7210
rect -5775 7150 -5760 7170
rect -5740 7150 -5725 7170
rect -5775 7130 -5725 7150
rect -5665 7165 -3165 7175
rect -5665 7145 -5650 7165
rect -5630 7145 -5610 7165
rect -5590 7145 -5570 7165
rect -5550 7145 -5530 7165
rect -5510 7145 -5490 7165
rect -5470 7145 -5450 7165
rect -5430 7145 -5410 7165
rect -5390 7145 -5370 7165
rect -5350 7145 -5330 7165
rect -5310 7145 -5290 7165
rect -5270 7145 -5250 7165
rect -5230 7145 -5210 7165
rect -5190 7145 -5170 7165
rect -5150 7145 -5130 7165
rect -5110 7145 -5090 7165
rect -5070 7145 -5050 7165
rect -5030 7145 -5010 7165
rect -4990 7145 -4970 7165
rect -4950 7145 -4930 7165
rect -4910 7145 -4890 7165
rect -4870 7145 -4850 7165
rect -4830 7145 -4810 7165
rect -4790 7145 -4770 7165
rect -4750 7145 -4730 7165
rect -4710 7145 -4690 7165
rect -4670 7145 -4650 7165
rect -4630 7145 -4610 7165
rect -4590 7145 -4570 7165
rect -4550 7145 -4530 7165
rect -4510 7145 -4490 7165
rect -4470 7145 -4450 7165
rect -4430 7145 -4410 7165
rect -4390 7145 -4370 7165
rect -4350 7145 -4330 7165
rect -4310 7145 -4290 7165
rect -4270 7145 -4250 7165
rect -4230 7145 -4210 7165
rect -4190 7145 -4170 7165
rect -4150 7145 -4130 7165
rect -4110 7145 -4090 7165
rect -4070 7145 -4050 7165
rect -4030 7145 -4010 7165
rect -3990 7145 -3970 7165
rect -3950 7145 -3930 7165
rect -3910 7145 -3890 7165
rect -3870 7145 -3850 7165
rect -3830 7145 -3810 7165
rect -3790 7145 -3770 7165
rect -3750 7145 -3730 7165
rect -3710 7145 -3690 7165
rect -3670 7145 -3650 7165
rect -3630 7145 -3610 7165
rect -3590 7145 -3570 7165
rect -3550 7145 -3530 7165
rect -3510 7145 -3490 7165
rect -3470 7145 -3450 7165
rect -3430 7145 -3410 7165
rect -3390 7145 -3370 7165
rect -3350 7145 -3330 7165
rect -3310 7145 -3290 7165
rect -3270 7145 -3250 7165
rect -3230 7145 -3210 7165
rect -3190 7145 -3165 7165
rect -5665 7135 -3165 7145
rect -2965 7170 -2915 7190
rect -2965 7150 -2950 7170
rect -2930 7150 -2915 7170
rect -5775 7110 -5760 7130
rect -5740 7110 -5725 7130
rect -5775 7090 -5725 7110
rect -3145 7125 -2990 7135
rect -3120 7105 -3100 7125
rect -3080 7105 -3060 7125
rect -3040 7105 -3020 7125
rect -3000 7105 -2990 7125
rect -3145 7095 -2990 7105
rect -2965 7130 -2915 7150
rect -2965 7110 -2950 7130
rect -2930 7110 -2915 7130
rect -5775 7070 -5760 7090
rect -5740 7070 -5725 7090
rect -5775 7050 -5725 7070
rect -5665 7083 -3165 7093
rect -5665 7063 -5650 7083
rect -5630 7063 -5610 7083
rect -5590 7063 -5570 7083
rect -5550 7063 -5530 7083
rect -5510 7063 -5490 7083
rect -5470 7063 -5450 7083
rect -5430 7063 -5410 7083
rect -5390 7063 -5370 7083
rect -5350 7063 -5330 7083
rect -5310 7063 -5290 7083
rect -5270 7063 -5250 7083
rect -5230 7063 -5210 7083
rect -5190 7063 -5170 7083
rect -5150 7063 -5130 7083
rect -5110 7063 -5090 7083
rect -5070 7063 -5050 7083
rect -5030 7063 -5010 7083
rect -4990 7063 -4970 7083
rect -4950 7063 -4930 7083
rect -4910 7063 -4890 7083
rect -4870 7063 -4850 7083
rect -4830 7063 -4810 7083
rect -4790 7063 -4770 7083
rect -4750 7063 -4730 7083
rect -4710 7063 -4690 7083
rect -4670 7063 -4650 7083
rect -4630 7063 -4610 7083
rect -4590 7063 -4570 7083
rect -4550 7063 -4530 7083
rect -4510 7063 -4490 7083
rect -4470 7063 -4450 7083
rect -4430 7063 -4410 7083
rect -4390 7063 -4370 7083
rect -4350 7063 -4330 7083
rect -4310 7063 -4290 7083
rect -4270 7063 -4250 7083
rect -4230 7063 -4210 7083
rect -4190 7063 -4170 7083
rect -4150 7063 -4130 7083
rect -4110 7063 -4090 7083
rect -4070 7063 -4050 7083
rect -4030 7063 -4010 7083
rect -3990 7063 -3970 7083
rect -3950 7063 -3930 7083
rect -3910 7063 -3890 7083
rect -3870 7063 -3850 7083
rect -3830 7063 -3810 7083
rect -3790 7063 -3770 7083
rect -3750 7063 -3730 7083
rect -3710 7063 -3690 7083
rect -3670 7063 -3650 7083
rect -3630 7063 -3610 7083
rect -3590 7063 -3570 7083
rect -3550 7063 -3530 7083
rect -3510 7063 -3490 7083
rect -3470 7063 -3450 7083
rect -3430 7063 -3410 7083
rect -3390 7063 -3370 7083
rect -3350 7063 -3330 7083
rect -3310 7063 -3290 7083
rect -3270 7063 -3250 7083
rect -3230 7063 -3210 7083
rect -3190 7063 -3165 7083
rect -5665 7053 -3165 7063
rect -2965 7090 -2915 7110
rect -2965 7070 -2950 7090
rect -2930 7070 -2915 7090
rect -2965 7050 -2915 7070
rect -5775 7030 -5760 7050
rect -5740 7030 -5725 7050
rect -5775 7010 -5725 7030
rect -3145 7040 -2990 7050
rect -3120 7020 -3100 7040
rect -3080 7020 -3060 7040
rect -3040 7020 -3020 7040
rect -3000 7020 -2990 7040
rect -5775 6990 -5760 7010
rect -5740 6990 -5725 7010
rect -5775 6970 -5725 6990
rect -5665 7001 -3165 7011
rect -3145 7010 -2990 7020
rect -2965 7030 -2950 7050
rect -2930 7030 -2915 7050
rect -2965 7010 -2915 7030
rect -5665 6981 -5650 7001
rect -5630 6981 -5610 7001
rect -5590 6981 -5570 7001
rect -5550 6981 -5530 7001
rect -5510 6981 -5490 7001
rect -5470 6981 -5450 7001
rect -5430 6981 -5410 7001
rect -5390 6981 -5370 7001
rect -5350 6981 -5330 7001
rect -5310 6981 -5290 7001
rect -5270 6981 -5250 7001
rect -5230 6981 -5210 7001
rect -5190 6981 -5170 7001
rect -5150 6981 -5130 7001
rect -5110 6981 -5090 7001
rect -5070 6981 -5050 7001
rect -5030 6981 -5010 7001
rect -4990 6981 -4970 7001
rect -4950 6981 -4930 7001
rect -4910 6981 -4890 7001
rect -4870 6981 -4850 7001
rect -4830 6981 -4810 7001
rect -4790 6981 -4770 7001
rect -4750 6981 -4730 7001
rect -4710 6981 -4690 7001
rect -4670 6981 -4650 7001
rect -4630 6981 -4610 7001
rect -4590 6981 -4570 7001
rect -4550 6981 -4530 7001
rect -4510 6981 -4490 7001
rect -4470 6981 -4450 7001
rect -4430 6981 -4410 7001
rect -4390 6981 -4370 7001
rect -4350 6981 -4330 7001
rect -4310 6981 -4290 7001
rect -4270 6981 -4250 7001
rect -4230 6981 -4210 7001
rect -4190 6981 -4170 7001
rect -4150 6981 -4130 7001
rect -4110 6981 -4090 7001
rect -4070 6981 -4050 7001
rect -4030 6981 -4010 7001
rect -3990 6981 -3970 7001
rect -3950 6981 -3930 7001
rect -3910 6981 -3890 7001
rect -3870 6981 -3850 7001
rect -3830 6981 -3810 7001
rect -3790 6981 -3770 7001
rect -3750 6981 -3730 7001
rect -3710 6981 -3690 7001
rect -3670 6981 -3650 7001
rect -3630 6981 -3610 7001
rect -3590 6981 -3570 7001
rect -3550 6981 -3530 7001
rect -3510 6981 -3490 7001
rect -3470 6981 -3450 7001
rect -3430 6981 -3410 7001
rect -3390 6981 -3370 7001
rect -3350 6981 -3330 7001
rect -3310 6981 -3290 7001
rect -3270 6981 -3250 7001
rect -3230 6981 -3210 7001
rect -3190 6981 -3165 7001
rect -5665 6971 -3165 6981
rect -2965 6990 -2950 7010
rect -2930 6990 -2915 7010
rect -2965 6970 -2915 6990
rect -5775 6950 -5760 6970
rect -5740 6950 -5725 6970
rect -5775 6930 -5725 6950
rect -3145 6960 -2990 6970
rect -3120 6940 -3100 6960
rect -3080 6940 -3060 6960
rect -3040 6940 -3020 6960
rect -3000 6940 -2990 6960
rect -3145 6930 -2990 6940
rect -2965 6950 -2950 6970
rect -2930 6950 -2915 6970
rect -2965 6930 -2915 6950
rect -5775 6910 -5760 6930
rect -5740 6910 -5725 6930
rect -5775 6890 -5725 6910
rect -5775 6870 -5760 6890
rect -5740 6870 -5725 6890
rect -5665 6919 -3165 6929
rect -5665 6899 -5650 6919
rect -5630 6899 -5610 6919
rect -5590 6899 -5570 6919
rect -5550 6899 -5530 6919
rect -5510 6899 -5490 6919
rect -5470 6899 -5450 6919
rect -5430 6899 -5410 6919
rect -5390 6899 -5370 6919
rect -5350 6899 -5330 6919
rect -5310 6899 -5290 6919
rect -5270 6899 -5250 6919
rect -5230 6899 -5210 6919
rect -5190 6899 -5170 6919
rect -5150 6899 -5130 6919
rect -5110 6899 -5090 6919
rect -5070 6899 -5050 6919
rect -5030 6899 -5010 6919
rect -4990 6899 -4970 6919
rect -4950 6899 -4930 6919
rect -4910 6899 -4890 6919
rect -4870 6899 -4850 6919
rect -4830 6899 -4810 6919
rect -4790 6899 -4770 6919
rect -4750 6899 -4730 6919
rect -4710 6899 -4690 6919
rect -4670 6899 -4650 6919
rect -4630 6899 -4610 6919
rect -4590 6899 -4570 6919
rect -4550 6899 -4530 6919
rect -4510 6899 -4490 6919
rect -4470 6899 -4450 6919
rect -4430 6899 -4410 6919
rect -4390 6899 -4370 6919
rect -4350 6899 -4330 6919
rect -4310 6899 -4290 6919
rect -4270 6899 -4250 6919
rect -4230 6899 -4210 6919
rect -4190 6899 -4170 6919
rect -4150 6899 -4130 6919
rect -4110 6899 -4090 6919
rect -4070 6899 -4050 6919
rect -4030 6899 -4010 6919
rect -3990 6899 -3970 6919
rect -3950 6899 -3930 6919
rect -3910 6899 -3890 6919
rect -3870 6899 -3850 6919
rect -3830 6899 -3810 6919
rect -3790 6899 -3770 6919
rect -3750 6899 -3730 6919
rect -3710 6899 -3690 6919
rect -3670 6899 -3650 6919
rect -3630 6899 -3610 6919
rect -3590 6899 -3570 6919
rect -3550 6899 -3530 6919
rect -3510 6899 -3490 6919
rect -3470 6899 -3450 6919
rect -3430 6899 -3410 6919
rect -3390 6899 -3370 6919
rect -3350 6899 -3330 6919
rect -3310 6899 -3290 6919
rect -3270 6899 -3250 6919
rect -3230 6899 -3210 6919
rect -3190 6899 -3165 6919
rect -5665 6889 -3165 6899
rect -2965 6910 -2950 6930
rect -2930 6910 -2915 6930
rect -2965 6890 -2915 6910
rect -5775 6850 -5725 6870
rect -3145 6880 -2990 6890
rect -3120 6860 -3100 6880
rect -3080 6860 -3060 6880
rect -3040 6860 -3020 6880
rect -3000 6860 -2990 6880
rect -3145 6850 -2990 6860
rect -2965 6870 -2950 6890
rect -2930 6870 -2915 6890
rect -2965 6850 -2915 6870
rect -5775 6830 -5760 6850
rect -5740 6830 -5725 6850
rect -5775 6810 -5725 6830
rect -5775 6790 -5760 6810
rect -5740 6790 -5725 6810
rect -5665 6837 -3165 6847
rect -5665 6817 -5650 6837
rect -5630 6817 -5610 6837
rect -5590 6817 -5570 6837
rect -5550 6817 -5530 6837
rect -5510 6817 -5490 6837
rect -5470 6817 -5450 6837
rect -5430 6817 -5410 6837
rect -5390 6817 -5370 6837
rect -5350 6817 -5330 6837
rect -5310 6817 -5290 6837
rect -5270 6817 -5250 6837
rect -5230 6817 -5210 6837
rect -5190 6817 -5170 6837
rect -5150 6817 -5130 6837
rect -5110 6817 -5090 6837
rect -5070 6817 -5050 6837
rect -5030 6817 -5010 6837
rect -4990 6817 -4970 6837
rect -4950 6817 -4930 6837
rect -4910 6817 -4890 6837
rect -4870 6817 -4850 6837
rect -4830 6817 -4810 6837
rect -4790 6817 -4770 6837
rect -4750 6817 -4730 6837
rect -4710 6817 -4690 6837
rect -4670 6817 -4650 6837
rect -4630 6817 -4610 6837
rect -4590 6817 -4570 6837
rect -4550 6817 -4530 6837
rect -4510 6817 -4490 6837
rect -4470 6817 -4450 6837
rect -4430 6817 -4410 6837
rect -4390 6817 -4370 6837
rect -4350 6817 -4330 6837
rect -4310 6817 -4290 6837
rect -4270 6817 -4250 6837
rect -4230 6817 -4210 6837
rect -4190 6817 -4170 6837
rect -4150 6817 -4130 6837
rect -4110 6817 -4090 6837
rect -4070 6817 -4050 6837
rect -4030 6817 -4010 6837
rect -3990 6817 -3970 6837
rect -3950 6817 -3930 6837
rect -3910 6817 -3890 6837
rect -3870 6817 -3850 6837
rect -3830 6817 -3810 6837
rect -3790 6817 -3770 6837
rect -3750 6817 -3730 6837
rect -3710 6817 -3690 6837
rect -3670 6817 -3650 6837
rect -3630 6817 -3610 6837
rect -3590 6817 -3570 6837
rect -3550 6817 -3530 6837
rect -3510 6817 -3490 6837
rect -3470 6817 -3450 6837
rect -3430 6817 -3410 6837
rect -3390 6817 -3370 6837
rect -3350 6817 -3330 6837
rect -3310 6817 -3290 6837
rect -3270 6817 -3250 6837
rect -3230 6817 -3210 6837
rect -3190 6817 -3165 6837
rect -5665 6807 -3165 6817
rect -2965 6830 -2950 6850
rect -2930 6830 -2915 6850
rect -2965 6810 -2915 6830
rect -5775 6770 -5725 6790
rect -5775 6750 -5760 6770
rect -5740 6750 -5725 6770
rect -3145 6795 -2990 6805
rect -3120 6775 -3100 6795
rect -3080 6775 -3060 6795
rect -3040 6775 -3020 6795
rect -3000 6775 -2990 6795
rect -3145 6765 -2990 6775
rect -2965 6790 -2950 6810
rect -2930 6790 -2915 6810
rect -2965 6770 -2915 6790
rect -5775 6730 -5725 6750
rect -5775 6710 -5760 6730
rect -5740 6710 -5725 6730
rect -5665 6755 -3165 6765
rect -5665 6735 -5650 6755
rect -5630 6735 -5610 6755
rect -5590 6735 -5570 6755
rect -5550 6735 -5530 6755
rect -5510 6735 -5490 6755
rect -5470 6735 -5450 6755
rect -5430 6735 -5410 6755
rect -5390 6735 -5370 6755
rect -5350 6735 -5330 6755
rect -5310 6735 -5290 6755
rect -5270 6735 -5250 6755
rect -5230 6735 -5210 6755
rect -5190 6735 -5170 6755
rect -5150 6735 -5130 6755
rect -5110 6735 -5090 6755
rect -5070 6735 -5050 6755
rect -5030 6735 -5010 6755
rect -4990 6735 -4970 6755
rect -4950 6735 -4930 6755
rect -4910 6735 -4890 6755
rect -4870 6735 -4850 6755
rect -4830 6735 -4810 6755
rect -4790 6735 -4770 6755
rect -4750 6735 -4730 6755
rect -4710 6735 -4690 6755
rect -4670 6735 -4650 6755
rect -4630 6735 -4610 6755
rect -4590 6735 -4570 6755
rect -4550 6735 -4530 6755
rect -4510 6735 -4490 6755
rect -4470 6735 -4450 6755
rect -4430 6735 -4410 6755
rect -4390 6735 -4370 6755
rect -4350 6735 -4330 6755
rect -4310 6735 -4290 6755
rect -4270 6735 -4250 6755
rect -4230 6735 -4210 6755
rect -4190 6735 -4170 6755
rect -4150 6735 -4130 6755
rect -4110 6735 -4090 6755
rect -4070 6735 -4050 6755
rect -4030 6735 -4010 6755
rect -3990 6735 -3970 6755
rect -3950 6735 -3930 6755
rect -3910 6735 -3890 6755
rect -3870 6735 -3850 6755
rect -3830 6735 -3810 6755
rect -3790 6735 -3770 6755
rect -3750 6735 -3730 6755
rect -3710 6735 -3690 6755
rect -3670 6735 -3650 6755
rect -3630 6735 -3610 6755
rect -3590 6735 -3570 6755
rect -3550 6735 -3530 6755
rect -3510 6735 -3490 6755
rect -3470 6735 -3450 6755
rect -3430 6735 -3410 6755
rect -3390 6735 -3370 6755
rect -3350 6735 -3330 6755
rect -3310 6735 -3290 6755
rect -3270 6735 -3250 6755
rect -3230 6735 -3210 6755
rect -3190 6735 -3165 6755
rect -5665 6725 -3165 6735
rect -2965 6750 -2950 6770
rect -2930 6750 -2915 6770
rect -2965 6730 -2915 6750
rect -5775 6690 -5725 6710
rect -5775 6670 -5760 6690
rect -5740 6670 -5725 6690
rect -3145 6715 -2990 6725
rect -3120 6695 -3100 6715
rect -3080 6695 -3060 6715
rect -3040 6695 -3020 6715
rect -3000 6695 -2990 6715
rect -3145 6685 -2990 6695
rect -2965 6710 -2950 6730
rect -2930 6710 -2915 6730
rect -2965 6690 -2915 6710
rect -5775 6650 -5725 6670
rect -5775 6630 -5760 6650
rect -5740 6630 -5725 6650
rect -5665 6673 -3165 6683
rect -5665 6653 -5650 6673
rect -5630 6653 -5610 6673
rect -5590 6653 -5570 6673
rect -5550 6653 -5530 6673
rect -5510 6653 -5490 6673
rect -5470 6653 -5450 6673
rect -5430 6653 -5410 6673
rect -5390 6653 -5370 6673
rect -5350 6653 -5330 6673
rect -5310 6653 -5290 6673
rect -5270 6653 -5250 6673
rect -5230 6653 -5210 6673
rect -5190 6653 -5170 6673
rect -5150 6653 -5130 6673
rect -5110 6653 -5090 6673
rect -5070 6653 -5050 6673
rect -5030 6653 -5010 6673
rect -4990 6653 -4970 6673
rect -4950 6653 -4930 6673
rect -4910 6653 -4890 6673
rect -4870 6653 -4850 6673
rect -4830 6653 -4810 6673
rect -4790 6653 -4770 6673
rect -4750 6653 -4730 6673
rect -4710 6653 -4690 6673
rect -4670 6653 -4650 6673
rect -4630 6653 -4610 6673
rect -4590 6653 -4570 6673
rect -4550 6653 -4530 6673
rect -4510 6653 -4490 6673
rect -4470 6653 -4450 6673
rect -4430 6653 -4410 6673
rect -4390 6653 -4370 6673
rect -4350 6653 -4330 6673
rect -4310 6653 -4290 6673
rect -4270 6653 -4250 6673
rect -4230 6653 -4210 6673
rect -4190 6653 -4170 6673
rect -4150 6653 -4130 6673
rect -4110 6653 -4090 6673
rect -4070 6653 -4050 6673
rect -4030 6653 -4010 6673
rect -3990 6653 -3970 6673
rect -3950 6653 -3930 6673
rect -3910 6653 -3890 6673
rect -3870 6653 -3850 6673
rect -3830 6653 -3810 6673
rect -3790 6653 -3770 6673
rect -3750 6653 -3730 6673
rect -3710 6653 -3690 6673
rect -3670 6653 -3650 6673
rect -3630 6653 -3610 6673
rect -3590 6653 -3570 6673
rect -3550 6653 -3530 6673
rect -3510 6653 -3490 6673
rect -3470 6653 -3450 6673
rect -3430 6653 -3410 6673
rect -3390 6653 -3370 6673
rect -3350 6653 -3330 6673
rect -3310 6653 -3290 6673
rect -3270 6653 -3250 6673
rect -3230 6653 -3210 6673
rect -3190 6653 -3165 6673
rect -5665 6643 -3165 6653
rect -2965 6670 -2950 6690
rect -2930 6670 -2915 6690
rect -2965 6650 -2915 6670
rect -5775 6610 -5725 6630
rect -5775 6590 -5760 6610
rect -5740 6590 -5725 6610
rect -3145 6635 -2990 6645
rect -3120 6615 -3100 6635
rect -3080 6615 -3060 6635
rect -3040 6615 -3020 6635
rect -3000 6615 -2990 6635
rect -3145 6605 -2990 6615
rect -2965 6630 -2950 6650
rect -2930 6630 -2915 6650
rect -2965 6610 -2915 6630
rect -5775 6570 -5725 6590
rect -5775 6550 -5760 6570
rect -5740 6550 -5725 6570
rect -5665 6591 -3165 6601
rect -5665 6571 -5650 6591
rect -5630 6571 -5610 6591
rect -5590 6571 -5570 6591
rect -5550 6571 -5530 6591
rect -5510 6571 -5490 6591
rect -5470 6571 -5450 6591
rect -5430 6571 -5410 6591
rect -5390 6571 -5370 6591
rect -5350 6571 -5330 6591
rect -5310 6571 -5290 6591
rect -5270 6571 -5250 6591
rect -5230 6571 -5210 6591
rect -5190 6571 -5170 6591
rect -5150 6571 -5130 6591
rect -5110 6571 -5090 6591
rect -5070 6571 -5050 6591
rect -5030 6571 -5010 6591
rect -4990 6571 -4970 6591
rect -4950 6571 -4930 6591
rect -4910 6571 -4890 6591
rect -4870 6571 -4850 6591
rect -4830 6571 -4810 6591
rect -4790 6571 -4770 6591
rect -4750 6571 -4730 6591
rect -4710 6571 -4690 6591
rect -4670 6571 -4650 6591
rect -4630 6571 -4610 6591
rect -4590 6571 -4570 6591
rect -4550 6571 -4530 6591
rect -4510 6571 -4490 6591
rect -4470 6571 -4450 6591
rect -4430 6571 -4410 6591
rect -4390 6571 -4370 6591
rect -4350 6571 -4330 6591
rect -4310 6571 -4290 6591
rect -4270 6571 -4250 6591
rect -4230 6571 -4210 6591
rect -4190 6571 -4170 6591
rect -4150 6571 -4130 6591
rect -4110 6571 -4090 6591
rect -4070 6571 -4050 6591
rect -4030 6571 -4010 6591
rect -3990 6571 -3970 6591
rect -3950 6571 -3930 6591
rect -3910 6571 -3890 6591
rect -3870 6571 -3850 6591
rect -3830 6571 -3810 6591
rect -3790 6571 -3770 6591
rect -3750 6571 -3730 6591
rect -3710 6571 -3690 6591
rect -3670 6571 -3650 6591
rect -3630 6571 -3610 6591
rect -3590 6571 -3570 6591
rect -3550 6571 -3530 6591
rect -3510 6571 -3490 6591
rect -3470 6571 -3450 6591
rect -3430 6571 -3410 6591
rect -3390 6571 -3370 6591
rect -3350 6571 -3330 6591
rect -3310 6571 -3290 6591
rect -3270 6571 -3250 6591
rect -3230 6571 -3210 6591
rect -3190 6571 -3165 6591
rect -5665 6561 -3165 6571
rect -2965 6590 -2950 6610
rect -2930 6590 -2915 6610
rect -2965 6570 -2915 6590
rect -5775 6530 -5725 6550
rect -5775 6510 -5760 6530
rect -5740 6510 -5725 6530
rect -3145 6550 -2990 6560
rect -3120 6530 -3100 6550
rect -3080 6530 -3060 6550
rect -3040 6530 -3020 6550
rect -3000 6530 -2990 6550
rect -3145 6520 -2990 6530
rect -2965 6550 -2950 6570
rect -2930 6550 -2915 6570
rect -2965 6530 -2915 6550
rect -5775 6490 -5725 6510
rect -5775 6470 -5760 6490
rect -5740 6470 -5725 6490
rect -5665 6509 -3165 6519
rect -5665 6489 -5650 6509
rect -5630 6489 -5610 6509
rect -5590 6489 -5570 6509
rect -5550 6489 -5530 6509
rect -5510 6489 -5490 6509
rect -5470 6489 -5450 6509
rect -5430 6489 -5410 6509
rect -5390 6489 -5370 6509
rect -5350 6489 -5330 6509
rect -5310 6489 -5290 6509
rect -5270 6489 -5250 6509
rect -5230 6489 -5210 6509
rect -5190 6489 -5170 6509
rect -5150 6489 -5130 6509
rect -5110 6489 -5090 6509
rect -5070 6489 -5050 6509
rect -5030 6489 -5010 6509
rect -4990 6489 -4970 6509
rect -4950 6489 -4930 6509
rect -4910 6489 -4890 6509
rect -4870 6489 -4850 6509
rect -4830 6489 -4810 6509
rect -4790 6489 -4770 6509
rect -4750 6489 -4730 6509
rect -4710 6489 -4690 6509
rect -4670 6489 -4650 6509
rect -4630 6489 -4610 6509
rect -4590 6489 -4570 6509
rect -4550 6489 -4530 6509
rect -4510 6489 -4490 6509
rect -4470 6489 -4450 6509
rect -4430 6489 -4410 6509
rect -4390 6489 -4370 6509
rect -4350 6489 -4330 6509
rect -4310 6489 -4290 6509
rect -4270 6489 -4250 6509
rect -4230 6489 -4210 6509
rect -4190 6489 -4170 6509
rect -4150 6489 -4130 6509
rect -4110 6489 -4090 6509
rect -4070 6489 -4050 6509
rect -4030 6489 -4010 6509
rect -3990 6489 -3970 6509
rect -3950 6489 -3930 6509
rect -3910 6489 -3890 6509
rect -3870 6489 -3850 6509
rect -3830 6489 -3810 6509
rect -3790 6489 -3770 6509
rect -3750 6489 -3730 6509
rect -3710 6489 -3690 6509
rect -3670 6489 -3650 6509
rect -3630 6489 -3610 6509
rect -3590 6489 -3570 6509
rect -3550 6489 -3530 6509
rect -3510 6489 -3490 6509
rect -3470 6489 -3450 6509
rect -3430 6489 -3410 6509
rect -3390 6489 -3370 6509
rect -3350 6489 -3330 6509
rect -3310 6489 -3290 6509
rect -3270 6489 -3250 6509
rect -3230 6489 -3210 6509
rect -3190 6489 -3165 6509
rect -5665 6479 -3165 6489
rect -2965 6510 -2950 6530
rect -2930 6510 -2915 6530
rect -2965 6490 -2915 6510
rect -5775 6450 -5725 6470
rect -5775 6430 -5760 6450
rect -5740 6430 -5725 6450
rect -3145 6470 -2990 6480
rect -3120 6450 -3100 6470
rect -3080 6450 -3060 6470
rect -3040 6450 -3020 6470
rect -3000 6450 -2990 6470
rect -3145 6440 -2990 6450
rect -2965 6470 -2950 6490
rect -2930 6470 -2915 6490
rect -2965 6450 -2915 6470
rect -5775 6410 -5725 6430
rect -5775 6390 -5760 6410
rect -5740 6390 -5725 6410
rect -5665 6427 -3165 6437
rect -5665 6407 -5650 6427
rect -5630 6407 -5610 6427
rect -5590 6407 -5570 6427
rect -5550 6407 -5530 6427
rect -5510 6407 -5490 6427
rect -5470 6407 -5450 6427
rect -5430 6407 -5410 6427
rect -5390 6407 -5370 6427
rect -5350 6407 -5330 6427
rect -5310 6407 -5290 6427
rect -5270 6407 -5250 6427
rect -5230 6407 -5210 6427
rect -5190 6407 -5170 6427
rect -5150 6407 -5130 6427
rect -5110 6407 -5090 6427
rect -5070 6407 -5050 6427
rect -5030 6407 -5010 6427
rect -4990 6407 -4970 6427
rect -4950 6407 -4930 6427
rect -4910 6407 -4890 6427
rect -4870 6407 -4850 6427
rect -4830 6407 -4810 6427
rect -4790 6407 -4770 6427
rect -4750 6407 -4730 6427
rect -4710 6407 -4690 6427
rect -4670 6407 -4650 6427
rect -4630 6407 -4610 6427
rect -4590 6407 -4570 6427
rect -4550 6407 -4530 6427
rect -4510 6407 -4490 6427
rect -4470 6407 -4450 6427
rect -4430 6407 -4410 6427
rect -4390 6407 -4370 6427
rect -4350 6407 -4330 6427
rect -4310 6407 -4290 6427
rect -4270 6407 -4250 6427
rect -4230 6407 -4210 6427
rect -4190 6407 -4170 6427
rect -4150 6407 -4130 6427
rect -4110 6407 -4090 6427
rect -4070 6407 -4050 6427
rect -4030 6407 -4010 6427
rect -3990 6407 -3970 6427
rect -3950 6407 -3930 6427
rect -3910 6407 -3890 6427
rect -3870 6407 -3850 6427
rect -3830 6407 -3810 6427
rect -3790 6407 -3770 6427
rect -3750 6407 -3730 6427
rect -3710 6407 -3690 6427
rect -3670 6407 -3650 6427
rect -3630 6407 -3610 6427
rect -3590 6407 -3570 6427
rect -3550 6407 -3530 6427
rect -3510 6407 -3490 6427
rect -3470 6407 -3450 6427
rect -3430 6407 -3410 6427
rect -3390 6407 -3370 6427
rect -3350 6407 -3330 6427
rect -3310 6407 -3290 6427
rect -3270 6407 -3250 6427
rect -3230 6407 -3210 6427
rect -3190 6407 -3165 6427
rect -5665 6397 -3165 6407
rect -2965 6430 -2950 6450
rect -2930 6430 -2915 6450
rect -2965 6410 -2915 6430
rect -5775 6370 -5725 6390
rect -5775 6350 -5760 6370
rect -5740 6350 -5725 6370
rect -3145 6390 -2990 6400
rect -3120 6370 -3100 6390
rect -3080 6370 -3060 6390
rect -3040 6370 -3020 6390
rect -3000 6370 -2990 6390
rect -3145 6360 -2990 6370
rect -2965 6390 -2950 6410
rect -2930 6390 -2915 6410
rect -2965 6370 -2915 6390
rect -5775 6330 -5725 6350
rect -5775 6310 -5760 6330
rect -5740 6310 -5725 6330
rect -5775 6290 -5725 6310
rect -5775 6270 -5760 6290
rect -5740 6270 -5725 6290
rect -5665 6345 -3165 6355
rect -5665 6325 -5650 6345
rect -5630 6325 -5610 6345
rect -5590 6325 -5570 6345
rect -5550 6325 -5530 6345
rect -5510 6325 -5490 6345
rect -5470 6325 -5450 6345
rect -5430 6325 -5410 6345
rect -5390 6325 -5370 6345
rect -5350 6325 -5330 6345
rect -5310 6325 -5290 6345
rect -5270 6325 -5250 6345
rect -5230 6325 -5210 6345
rect -5190 6325 -5170 6345
rect -5150 6325 -5130 6345
rect -5110 6325 -5090 6345
rect -5070 6325 -5050 6345
rect -5030 6325 -5010 6345
rect -4990 6325 -4970 6345
rect -4950 6325 -4930 6345
rect -4910 6325 -4890 6345
rect -4870 6325 -4850 6345
rect -4830 6325 -4810 6345
rect -4790 6325 -4770 6345
rect -4750 6325 -4730 6345
rect -4710 6325 -4690 6345
rect -4670 6325 -4650 6345
rect -4630 6325 -4610 6345
rect -4590 6325 -4570 6345
rect -4550 6325 -4530 6345
rect -4510 6325 -4490 6345
rect -4470 6325 -4450 6345
rect -4430 6325 -4410 6345
rect -4390 6325 -4370 6345
rect -4350 6325 -4330 6345
rect -4310 6325 -4290 6345
rect -4270 6325 -4250 6345
rect -4230 6325 -4210 6345
rect -4190 6325 -4170 6345
rect -4150 6325 -4130 6345
rect -4110 6325 -4090 6345
rect -4070 6325 -4050 6345
rect -4030 6325 -4010 6345
rect -3990 6325 -3970 6345
rect -3950 6325 -3930 6345
rect -3910 6325 -3890 6345
rect -3870 6325 -3850 6345
rect -3830 6325 -3810 6345
rect -3790 6325 -3770 6345
rect -3750 6325 -3730 6345
rect -3710 6325 -3690 6345
rect -3670 6325 -3650 6345
rect -3630 6325 -3610 6345
rect -3590 6325 -3570 6345
rect -3550 6325 -3530 6345
rect -3510 6325 -3490 6345
rect -3470 6325 -3450 6345
rect -3430 6325 -3410 6345
rect -3390 6325 -3370 6345
rect -3350 6325 -3330 6345
rect -3310 6325 -3290 6345
rect -3270 6325 -3250 6345
rect -3230 6325 -3210 6345
rect -3190 6325 -3165 6345
rect -5665 6305 -3165 6325
rect -5665 6285 -5650 6305
rect -5630 6285 -5610 6305
rect -5590 6285 -5570 6305
rect -5550 6285 -5530 6305
rect -5510 6285 -5490 6305
rect -5470 6285 -5450 6305
rect -5430 6285 -5410 6305
rect -5390 6285 -5370 6305
rect -5350 6285 -5330 6305
rect -5310 6285 -5290 6305
rect -5270 6285 -5250 6305
rect -5230 6285 -5210 6305
rect -5190 6285 -5170 6305
rect -5150 6285 -5130 6305
rect -5110 6285 -5090 6305
rect -5070 6285 -5050 6305
rect -5030 6285 -5010 6305
rect -4990 6285 -4970 6305
rect -4950 6285 -4930 6305
rect -4910 6285 -4890 6305
rect -4870 6285 -4850 6305
rect -4830 6285 -4810 6305
rect -4790 6285 -4770 6305
rect -4750 6285 -4730 6305
rect -4710 6285 -4690 6305
rect -4670 6285 -4650 6305
rect -4630 6285 -4610 6305
rect -4590 6285 -4570 6305
rect -4550 6285 -4530 6305
rect -4510 6285 -4490 6305
rect -4470 6285 -4450 6305
rect -4430 6285 -4410 6305
rect -4390 6285 -4370 6305
rect -4350 6285 -4330 6305
rect -4310 6285 -4290 6305
rect -4270 6285 -4250 6305
rect -4230 6285 -4210 6305
rect -4190 6285 -4170 6305
rect -4150 6285 -4130 6305
rect -4110 6285 -4090 6305
rect -4070 6285 -4050 6305
rect -4030 6285 -4010 6305
rect -3990 6285 -3970 6305
rect -3950 6285 -3930 6305
rect -3910 6285 -3890 6305
rect -3870 6285 -3850 6305
rect -3830 6285 -3810 6305
rect -3790 6285 -3770 6305
rect -3750 6285 -3730 6305
rect -3710 6285 -3690 6305
rect -3670 6285 -3650 6305
rect -3630 6285 -3610 6305
rect -3590 6285 -3570 6305
rect -3550 6285 -3530 6305
rect -3510 6285 -3490 6305
rect -3470 6285 -3450 6305
rect -3430 6285 -3410 6305
rect -3390 6285 -3370 6305
rect -3350 6285 -3330 6305
rect -3310 6285 -3290 6305
rect -3270 6285 -3250 6305
rect -3230 6285 -3210 6305
rect -3190 6285 -3165 6305
rect -5665 6275 -3165 6285
rect -2965 6350 -2950 6370
rect -2930 6350 -2915 6370
rect -2965 6330 -2915 6350
rect -2965 6310 -2950 6330
rect -2930 6310 -2915 6330
rect -2965 6290 -2915 6310
rect -5775 6250 -5725 6270
rect -5775 6230 -5760 6250
rect -5740 6235 -5725 6250
rect -2965 6270 -2950 6290
rect -2930 6270 -2915 6290
rect -2965 6250 -2915 6270
rect -2965 6235 -2950 6250
rect -5740 6230 -2950 6235
rect -2930 6230 -2915 6250
rect -5775 6220 -2915 6230
rect -5775 6200 -5710 6220
rect -5690 6200 -5670 6220
rect -5650 6200 -5630 6220
rect -5610 6200 -5590 6220
rect -5570 6200 -5550 6220
rect -5530 6200 -5510 6220
rect -5490 6200 -5470 6220
rect -5450 6200 -5430 6220
rect -5410 6200 -5390 6220
rect -5370 6200 -5350 6220
rect -5330 6200 -5310 6220
rect -5290 6200 -5270 6220
rect -5250 6200 -5230 6220
rect -5210 6200 -5190 6220
rect -5170 6200 -5150 6220
rect -5130 6200 -5110 6220
rect -5090 6200 -5070 6220
rect -5050 6200 -5030 6220
rect -5010 6200 -4990 6220
rect -4970 6200 -4950 6220
rect -4930 6200 -4910 6220
rect -4890 6200 -4870 6220
rect -4850 6200 -4830 6220
rect -4810 6200 -4790 6220
rect -4770 6200 -4750 6220
rect -4730 6200 -4710 6220
rect -4690 6200 -4670 6220
rect -4650 6200 -4630 6220
rect -4610 6200 -4590 6220
rect -4570 6200 -4550 6220
rect -4530 6200 -4510 6220
rect -4490 6200 -4470 6220
rect -4450 6200 -4430 6220
rect -4410 6200 -4390 6220
rect -4370 6200 -4350 6220
rect -4330 6200 -4310 6220
rect -4290 6200 -4270 6220
rect -4250 6200 -4230 6220
rect -4210 6200 -4190 6220
rect -4170 6200 -4150 6220
rect -4130 6200 -4110 6220
rect -4090 6200 -4070 6220
rect -4050 6200 -4030 6220
rect -4010 6200 -3990 6220
rect -3970 6200 -3950 6220
rect -3930 6200 -3910 6220
rect -3890 6200 -3870 6220
rect -3850 6200 -3830 6220
rect -3810 6200 -3790 6220
rect -3770 6200 -3750 6220
rect -3730 6200 -3710 6220
rect -3690 6200 -3670 6220
rect -3650 6200 -3630 6220
rect -3610 6200 -3590 6220
rect -3570 6200 -3550 6220
rect -3530 6200 -3510 6220
rect -3490 6200 -3470 6220
rect -3450 6200 -3430 6220
rect -3410 6200 -3390 6220
rect -3370 6200 -3350 6220
rect -3330 6200 -3310 6220
rect -3290 6200 -3270 6220
rect -3250 6200 -3230 6220
rect -3210 6200 -3190 6220
rect -3170 6200 -3150 6220
rect -3130 6200 -3110 6220
rect -3090 6200 -3070 6220
rect -3050 6200 -3030 6220
rect -3010 6200 -2990 6220
rect -2970 6200 -2915 6220
rect -5775 6185 -2915 6200
rect -2225 8605 635 8620
rect -2225 8585 -2170 8605
rect -2150 8585 -2130 8605
rect -2110 8585 -2090 8605
rect -2070 8585 -2050 8605
rect -2030 8585 -2010 8605
rect -1990 8585 -1970 8605
rect -1950 8585 -1930 8605
rect -1910 8585 -1890 8605
rect -1870 8585 -1850 8605
rect -1830 8585 -1810 8605
rect -1790 8585 -1770 8605
rect -1750 8585 -1730 8605
rect -1710 8585 -1690 8605
rect -1670 8585 -1650 8605
rect -1630 8585 -1610 8605
rect -1590 8585 -1570 8605
rect -1550 8585 -1530 8605
rect -1510 8585 -1490 8605
rect -1470 8585 -1450 8605
rect -1430 8585 -1410 8605
rect -1390 8585 -1370 8605
rect -1350 8585 -1330 8605
rect -1310 8585 -1290 8605
rect -1270 8585 -1250 8605
rect -1230 8585 -1210 8605
rect -1190 8585 -1170 8605
rect -1150 8585 -1130 8605
rect -1110 8585 -1090 8605
rect -1070 8585 -1050 8605
rect -1030 8585 -1010 8605
rect -990 8585 -970 8605
rect -950 8585 -930 8605
rect -910 8585 -890 8605
rect -870 8585 -850 8605
rect -830 8585 -810 8605
rect -790 8585 -770 8605
rect -750 8585 -730 8605
rect -710 8585 -690 8605
rect -670 8585 -650 8605
rect -630 8585 -610 8605
rect -590 8585 -570 8605
rect -550 8585 -530 8605
rect -510 8585 -490 8605
rect -470 8585 -450 8605
rect -430 8585 -410 8605
rect -390 8585 -370 8605
rect -350 8585 -330 8605
rect -310 8585 -290 8605
rect -270 8585 -250 8605
rect -230 8585 -210 8605
rect -190 8585 -170 8605
rect -150 8585 -130 8605
rect -110 8585 -90 8605
rect -70 8585 -50 8605
rect -30 8585 -10 8605
rect 10 8585 30 8605
rect 50 8585 70 8605
rect 90 8585 110 8605
rect 130 8585 150 8605
rect 170 8585 190 8605
rect 210 8585 230 8605
rect 250 8585 270 8605
rect 290 8585 310 8605
rect 330 8585 350 8605
rect 370 8585 390 8605
rect 410 8585 430 8605
rect 450 8585 470 8605
rect 490 8585 510 8605
rect 530 8585 550 8605
rect 570 8585 635 8605
rect -2225 8570 635 8585
rect -2225 8550 -2210 8570
rect -2190 8550 -2175 8570
rect -2225 8530 -2175 8550
rect 585 8550 600 8570
rect 620 8550 635 8570
rect 585 8530 635 8550
rect -2225 8510 -2210 8530
rect -2190 8510 -2175 8530
rect -2225 8490 -2175 8510
rect -2225 8470 -2210 8490
rect -2190 8470 -2175 8490
rect -2225 8450 -2175 8470
rect -2225 8430 -2210 8450
rect -2190 8430 -2175 8450
rect -1975 8520 525 8530
rect -1975 8500 -1950 8520
rect -1930 8500 -1910 8520
rect -1890 8500 -1870 8520
rect -1850 8500 -1830 8520
rect -1810 8500 -1790 8520
rect -1770 8500 -1750 8520
rect -1730 8500 -1710 8520
rect -1690 8500 -1670 8520
rect -1650 8500 -1630 8520
rect -1610 8500 -1590 8520
rect -1570 8500 -1550 8520
rect -1530 8500 -1510 8520
rect -1490 8500 -1470 8520
rect -1450 8500 -1430 8520
rect -1410 8500 -1390 8520
rect -1370 8500 -1350 8520
rect -1330 8500 -1310 8520
rect -1290 8500 -1270 8520
rect -1250 8500 -1230 8520
rect -1210 8500 -1190 8520
rect -1170 8500 -1150 8520
rect -1130 8500 -1110 8520
rect -1090 8500 -1070 8520
rect -1050 8500 -1030 8520
rect -1010 8500 -990 8520
rect -970 8500 -950 8520
rect -930 8500 -910 8520
rect -890 8500 -870 8520
rect -850 8500 -830 8520
rect -810 8500 -790 8520
rect -770 8500 -750 8520
rect -730 8500 -710 8520
rect -690 8500 -670 8520
rect -650 8500 -630 8520
rect -610 8500 -590 8520
rect -570 8500 -550 8520
rect -530 8500 -510 8520
rect -490 8500 -470 8520
rect -450 8500 -430 8520
rect -410 8500 -390 8520
rect -370 8500 -350 8520
rect -330 8500 -310 8520
rect -290 8500 -270 8520
rect -250 8500 -230 8520
rect -210 8500 -190 8520
rect -170 8500 -150 8520
rect -130 8500 -110 8520
rect -90 8500 -70 8520
rect -50 8500 -30 8520
rect -10 8500 10 8520
rect 30 8500 50 8520
rect 70 8500 90 8520
rect 110 8500 130 8520
rect 150 8500 170 8520
rect 190 8500 210 8520
rect 230 8500 250 8520
rect 270 8500 290 8520
rect 310 8500 330 8520
rect 350 8500 370 8520
rect 390 8500 410 8520
rect 430 8500 450 8520
rect 470 8500 490 8520
rect 510 8500 525 8520
rect -1975 8477 525 8500
rect -1975 8457 -1950 8477
rect -1930 8457 -1910 8477
rect -1890 8457 -1870 8477
rect -1850 8457 -1830 8477
rect -1810 8457 -1790 8477
rect -1770 8457 -1750 8477
rect -1730 8457 -1710 8477
rect -1690 8457 -1670 8477
rect -1650 8457 -1630 8477
rect -1610 8457 -1590 8477
rect -1570 8457 -1550 8477
rect -1530 8457 -1510 8477
rect -1490 8457 -1470 8477
rect -1450 8457 -1430 8477
rect -1410 8457 -1390 8477
rect -1370 8457 -1350 8477
rect -1330 8457 -1310 8477
rect -1290 8457 -1270 8477
rect -1250 8457 -1230 8477
rect -1210 8457 -1190 8477
rect -1170 8457 -1150 8477
rect -1130 8457 -1110 8477
rect -1090 8457 -1070 8477
rect -1050 8457 -1030 8477
rect -1010 8457 -990 8477
rect -970 8457 -950 8477
rect -930 8457 -910 8477
rect -890 8457 -870 8477
rect -850 8457 -830 8477
rect -810 8457 -790 8477
rect -770 8457 -750 8477
rect -730 8457 -710 8477
rect -690 8457 -670 8477
rect -650 8457 -630 8477
rect -610 8457 -590 8477
rect -570 8457 -550 8477
rect -530 8457 -510 8477
rect -490 8457 -470 8477
rect -450 8457 -430 8477
rect -410 8457 -390 8477
rect -370 8457 -350 8477
rect -330 8457 -310 8477
rect -290 8457 -270 8477
rect -250 8457 -230 8477
rect -210 8457 -190 8477
rect -170 8457 -150 8477
rect -130 8457 -110 8477
rect -90 8457 -70 8477
rect -50 8457 -30 8477
rect -10 8457 10 8477
rect 30 8457 50 8477
rect 70 8457 90 8477
rect 110 8457 130 8477
rect 150 8457 170 8477
rect 190 8457 210 8477
rect 230 8457 250 8477
rect 270 8457 290 8477
rect 310 8457 330 8477
rect 350 8457 370 8477
rect 390 8457 410 8477
rect 430 8457 450 8477
rect 470 8457 490 8477
rect 510 8457 525 8477
rect -1975 8447 525 8457
rect 585 8510 600 8530
rect 620 8510 635 8530
rect 585 8490 635 8510
rect 585 8470 600 8490
rect 620 8470 635 8490
rect 585 8450 635 8470
rect -2225 8410 -2175 8430
rect -2225 8390 -2210 8410
rect -2190 8390 -2175 8410
rect -2150 8435 -1995 8445
rect -2150 8415 -2140 8435
rect -2120 8415 -2100 8435
rect -2080 8415 -2060 8435
rect -2040 8415 -2020 8435
rect -2150 8405 -1995 8415
rect 585 8430 600 8450
rect 620 8430 635 8450
rect 585 8410 635 8430
rect -2225 8370 -2175 8390
rect -2225 8350 -2210 8370
rect -2190 8350 -2175 8370
rect -1975 8395 525 8405
rect -1975 8375 -1950 8395
rect -1930 8375 -1910 8395
rect -1890 8375 -1870 8395
rect -1850 8375 -1830 8395
rect -1810 8375 -1790 8395
rect -1770 8375 -1750 8395
rect -1730 8375 -1710 8395
rect -1690 8375 -1670 8395
rect -1650 8375 -1630 8395
rect -1610 8375 -1590 8395
rect -1570 8375 -1550 8395
rect -1530 8375 -1510 8395
rect -1490 8375 -1470 8395
rect -1450 8375 -1430 8395
rect -1410 8375 -1390 8395
rect -1370 8375 -1350 8395
rect -1330 8375 -1310 8395
rect -1290 8375 -1270 8395
rect -1250 8375 -1230 8395
rect -1210 8375 -1190 8395
rect -1170 8375 -1150 8395
rect -1130 8375 -1110 8395
rect -1090 8375 -1070 8395
rect -1050 8375 -1030 8395
rect -1010 8375 -990 8395
rect -970 8375 -950 8395
rect -930 8375 -910 8395
rect -890 8375 -870 8395
rect -850 8375 -830 8395
rect -810 8375 -790 8395
rect -770 8375 -750 8395
rect -730 8375 -710 8395
rect -690 8375 -670 8395
rect -650 8375 -630 8395
rect -610 8375 -590 8395
rect -570 8375 -550 8395
rect -530 8375 -510 8395
rect -490 8375 -470 8395
rect -450 8375 -430 8395
rect -410 8375 -390 8395
rect -370 8375 -350 8395
rect -330 8375 -310 8395
rect -290 8375 -270 8395
rect -250 8375 -230 8395
rect -210 8375 -190 8395
rect -170 8375 -150 8395
rect -130 8375 -110 8395
rect -90 8375 -70 8395
rect -50 8375 -30 8395
rect -10 8375 10 8395
rect 30 8375 50 8395
rect 70 8375 90 8395
rect 110 8375 130 8395
rect 150 8375 170 8395
rect 190 8375 210 8395
rect 230 8375 250 8395
rect 270 8375 290 8395
rect 310 8375 330 8395
rect 350 8375 370 8395
rect 390 8375 410 8395
rect 430 8375 450 8395
rect 470 8375 490 8395
rect 510 8375 525 8395
rect -1975 8365 525 8375
rect 585 8390 600 8410
rect 620 8390 635 8410
rect 585 8370 635 8390
rect -2225 8330 -2175 8350
rect -2225 8310 -2210 8330
rect -2190 8310 -2175 8330
rect -2150 8355 -1995 8365
rect -2150 8335 -2140 8355
rect -2120 8335 -2100 8355
rect -2080 8335 -2060 8355
rect -2040 8335 -2020 8355
rect -2150 8325 -1995 8335
rect 585 8350 600 8370
rect 620 8350 635 8370
rect 585 8330 635 8350
rect -2225 8290 -2175 8310
rect -2225 8270 -2210 8290
rect -2190 8270 -2175 8290
rect -1975 8313 525 8323
rect -1975 8293 -1950 8313
rect -1930 8293 -1910 8313
rect -1890 8293 -1870 8313
rect -1850 8293 -1830 8313
rect -1810 8293 -1790 8313
rect -1770 8293 -1750 8313
rect -1730 8293 -1710 8313
rect -1690 8293 -1670 8313
rect -1650 8293 -1630 8313
rect -1610 8293 -1590 8313
rect -1570 8293 -1550 8313
rect -1530 8293 -1510 8313
rect -1490 8293 -1470 8313
rect -1450 8293 -1430 8313
rect -1410 8293 -1390 8313
rect -1370 8293 -1350 8313
rect -1330 8293 -1310 8313
rect -1290 8293 -1270 8313
rect -1250 8293 -1230 8313
rect -1210 8293 -1190 8313
rect -1170 8293 -1150 8313
rect -1130 8293 -1110 8313
rect -1090 8293 -1070 8313
rect -1050 8293 -1030 8313
rect -1010 8293 -990 8313
rect -970 8293 -950 8313
rect -930 8293 -910 8313
rect -890 8293 -870 8313
rect -850 8293 -830 8313
rect -810 8293 -790 8313
rect -770 8293 -750 8313
rect -730 8293 -710 8313
rect -690 8293 -670 8313
rect -650 8293 -630 8313
rect -610 8293 -590 8313
rect -570 8293 -550 8313
rect -530 8293 -510 8313
rect -490 8293 -470 8313
rect -450 8293 -430 8313
rect -410 8293 -390 8313
rect -370 8293 -350 8313
rect -330 8293 -310 8313
rect -290 8293 -270 8313
rect -250 8293 -230 8313
rect -210 8293 -190 8313
rect -170 8293 -150 8313
rect -130 8293 -110 8313
rect -90 8293 -70 8313
rect -50 8293 -30 8313
rect -10 8293 10 8313
rect 30 8293 50 8313
rect 70 8293 90 8313
rect 110 8293 130 8313
rect 150 8293 170 8313
rect 190 8293 210 8313
rect 230 8293 250 8313
rect 270 8293 290 8313
rect 310 8293 330 8313
rect 350 8293 370 8313
rect 390 8293 410 8313
rect 430 8293 450 8313
rect 470 8293 490 8313
rect 510 8293 525 8313
rect -1975 8283 525 8293
rect 585 8310 600 8330
rect 620 8310 635 8330
rect 585 8290 635 8310
rect -2225 8250 -2175 8270
rect -2225 8230 -2210 8250
rect -2190 8230 -2175 8250
rect -2150 8270 -1995 8280
rect -2150 8250 -2140 8270
rect -2120 8250 -2100 8270
rect -2080 8250 -2060 8270
rect -2040 8250 -2020 8270
rect -2150 8240 -1995 8250
rect 585 8270 600 8290
rect 620 8270 635 8290
rect 585 8250 635 8270
rect -2225 8210 -2175 8230
rect -2225 8190 -2210 8210
rect -2190 8190 -2175 8210
rect -1975 8231 525 8241
rect -1975 8211 -1950 8231
rect -1930 8211 -1910 8231
rect -1890 8211 -1870 8231
rect -1850 8211 -1830 8231
rect -1810 8211 -1790 8231
rect -1770 8211 -1750 8231
rect -1730 8211 -1710 8231
rect -1690 8211 -1670 8231
rect -1650 8211 -1630 8231
rect -1610 8211 -1590 8231
rect -1570 8211 -1550 8231
rect -1530 8211 -1510 8231
rect -1490 8211 -1470 8231
rect -1450 8211 -1430 8231
rect -1410 8211 -1390 8231
rect -1370 8211 -1350 8231
rect -1330 8211 -1310 8231
rect -1290 8211 -1270 8231
rect -1250 8211 -1230 8231
rect -1210 8211 -1190 8231
rect -1170 8211 -1150 8231
rect -1130 8211 -1110 8231
rect -1090 8211 -1070 8231
rect -1050 8211 -1030 8231
rect -1010 8211 -990 8231
rect -970 8211 -950 8231
rect -930 8211 -910 8231
rect -890 8211 -870 8231
rect -850 8211 -830 8231
rect -810 8211 -790 8231
rect -770 8211 -750 8231
rect -730 8211 -710 8231
rect -690 8211 -670 8231
rect -650 8211 -630 8231
rect -610 8211 -590 8231
rect -570 8211 -550 8231
rect -530 8211 -510 8231
rect -490 8211 -470 8231
rect -450 8211 -430 8231
rect -410 8211 -390 8231
rect -370 8211 -350 8231
rect -330 8211 -310 8231
rect -290 8211 -270 8231
rect -250 8211 -230 8231
rect -210 8211 -190 8231
rect -170 8211 -150 8231
rect -130 8211 -110 8231
rect -90 8211 -70 8231
rect -50 8211 -30 8231
rect -10 8211 10 8231
rect 30 8211 50 8231
rect 70 8211 90 8231
rect 110 8211 130 8231
rect 150 8211 170 8231
rect 190 8211 210 8231
rect 230 8211 250 8231
rect 270 8211 290 8231
rect 310 8211 330 8231
rect 350 8211 370 8231
rect 390 8211 410 8231
rect 430 8211 450 8231
rect 470 8211 490 8231
rect 510 8211 525 8231
rect -1975 8201 525 8211
rect 585 8230 600 8250
rect 620 8230 635 8250
rect 585 8210 635 8230
rect -2225 8170 -2175 8190
rect -2225 8150 -2210 8170
rect -2190 8150 -2175 8170
rect -2150 8190 -1995 8200
rect -2150 8170 -2140 8190
rect -2120 8170 -2100 8190
rect -2080 8170 -2060 8190
rect -2040 8170 -2020 8190
rect -2150 8160 -1995 8170
rect 585 8190 600 8210
rect 620 8190 635 8210
rect 585 8170 635 8190
rect -2225 8130 -2175 8150
rect -2225 8110 -2210 8130
rect -2190 8110 -2175 8130
rect -1975 8149 525 8159
rect -1975 8129 -1950 8149
rect -1930 8129 -1910 8149
rect -1890 8129 -1870 8149
rect -1850 8129 -1830 8149
rect -1810 8129 -1790 8149
rect -1770 8129 -1750 8149
rect -1730 8129 -1710 8149
rect -1690 8129 -1670 8149
rect -1650 8129 -1630 8149
rect -1610 8129 -1590 8149
rect -1570 8129 -1550 8149
rect -1530 8129 -1510 8149
rect -1490 8129 -1470 8149
rect -1450 8129 -1430 8149
rect -1410 8129 -1390 8149
rect -1370 8129 -1350 8149
rect -1330 8129 -1310 8149
rect -1290 8129 -1270 8149
rect -1250 8129 -1230 8149
rect -1210 8129 -1190 8149
rect -1170 8129 -1150 8149
rect -1130 8129 -1110 8149
rect -1090 8129 -1070 8149
rect -1050 8129 -1030 8149
rect -1010 8129 -990 8149
rect -970 8129 -950 8149
rect -930 8129 -910 8149
rect -890 8129 -870 8149
rect -850 8129 -830 8149
rect -810 8129 -790 8149
rect -770 8129 -750 8149
rect -730 8129 -710 8149
rect -690 8129 -670 8149
rect -650 8129 -630 8149
rect -610 8129 -590 8149
rect -570 8129 -550 8149
rect -530 8129 -510 8149
rect -490 8129 -470 8149
rect -450 8129 -430 8149
rect -410 8129 -390 8149
rect -370 8129 -350 8149
rect -330 8129 -310 8149
rect -290 8129 -270 8149
rect -250 8129 -230 8149
rect -210 8129 -190 8149
rect -170 8129 -150 8149
rect -130 8129 -110 8149
rect -90 8129 -70 8149
rect -50 8129 -30 8149
rect -10 8129 10 8149
rect 30 8129 50 8149
rect 70 8129 90 8149
rect 110 8129 130 8149
rect 150 8129 170 8149
rect 190 8129 210 8149
rect 230 8129 250 8149
rect 270 8129 290 8149
rect 310 8129 330 8149
rect 350 8129 370 8149
rect 390 8129 410 8149
rect 430 8129 450 8149
rect 470 8129 490 8149
rect 510 8129 525 8149
rect -2225 8090 -2175 8110
rect -2225 8070 -2210 8090
rect -2190 8070 -2175 8090
rect -2150 8110 -1995 8120
rect -1975 8119 525 8129
rect 585 8150 600 8170
rect 620 8150 635 8170
rect 585 8130 635 8150
rect -2150 8090 -2140 8110
rect -2120 8090 -2100 8110
rect -2080 8090 -2060 8110
rect -2040 8090 -2020 8110
rect -2150 8080 -1995 8090
rect 585 8110 600 8130
rect 620 8110 635 8130
rect 585 8090 635 8110
rect -2225 8050 -2175 8070
rect -2225 8030 -2210 8050
rect -2190 8030 -2175 8050
rect -1975 8067 525 8077
rect -1975 8047 -1950 8067
rect -1930 8047 -1910 8067
rect -1890 8047 -1870 8067
rect -1850 8047 -1830 8067
rect -1810 8047 -1790 8067
rect -1770 8047 -1750 8067
rect -1730 8047 -1710 8067
rect -1690 8047 -1670 8067
rect -1650 8047 -1630 8067
rect -1610 8047 -1590 8067
rect -1570 8047 -1550 8067
rect -1530 8047 -1510 8067
rect -1490 8047 -1470 8067
rect -1450 8047 -1430 8067
rect -1410 8047 -1390 8067
rect -1370 8047 -1350 8067
rect -1330 8047 -1310 8067
rect -1290 8047 -1270 8067
rect -1250 8047 -1230 8067
rect -1210 8047 -1190 8067
rect -1170 8047 -1150 8067
rect -1130 8047 -1110 8067
rect -1090 8047 -1070 8067
rect -1050 8047 -1030 8067
rect -1010 8047 -990 8067
rect -970 8047 -950 8067
rect -930 8047 -910 8067
rect -890 8047 -870 8067
rect -850 8047 -830 8067
rect -810 8047 -790 8067
rect -770 8047 -750 8067
rect -730 8047 -710 8067
rect -690 8047 -670 8067
rect -650 8047 -630 8067
rect -610 8047 -590 8067
rect -570 8047 -550 8067
rect -530 8047 -510 8067
rect -490 8047 -470 8067
rect -450 8047 -430 8067
rect -410 8047 -390 8067
rect -370 8047 -350 8067
rect -330 8047 -310 8067
rect -290 8047 -270 8067
rect -250 8047 -230 8067
rect -210 8047 -190 8067
rect -170 8047 -150 8067
rect -130 8047 -110 8067
rect -90 8047 -70 8067
rect -50 8047 -30 8067
rect -10 8047 10 8067
rect 30 8047 50 8067
rect 70 8047 90 8067
rect 110 8047 130 8067
rect 150 8047 170 8067
rect 190 8047 210 8067
rect 230 8047 250 8067
rect 270 8047 290 8067
rect 310 8047 330 8067
rect 350 8047 370 8067
rect 390 8047 410 8067
rect 430 8047 450 8067
rect 470 8047 490 8067
rect 510 8047 525 8067
rect -1975 8037 525 8047
rect 585 8070 600 8090
rect 620 8070 635 8090
rect 585 8050 635 8070
rect -2225 8010 -2175 8030
rect -2225 7990 -2210 8010
rect -2190 7990 -2175 8010
rect -2150 8025 -1995 8035
rect -2150 8005 -2140 8025
rect -2120 8005 -2100 8025
rect -2080 8005 -2060 8025
rect -2040 8005 -2020 8025
rect -2150 7995 -1995 8005
rect 585 8030 600 8050
rect 620 8030 635 8050
rect 585 8010 635 8030
rect -2225 7970 -2175 7990
rect -2225 7950 -2210 7970
rect -2190 7950 -2175 7970
rect -1975 7985 525 7995
rect -1975 7965 -1950 7985
rect -1930 7965 -1910 7985
rect -1890 7965 -1870 7985
rect -1850 7965 -1830 7985
rect -1810 7965 -1790 7985
rect -1770 7965 -1750 7985
rect -1730 7965 -1710 7985
rect -1690 7965 -1670 7985
rect -1650 7965 -1630 7985
rect -1610 7965 -1590 7985
rect -1570 7965 -1550 7985
rect -1530 7965 -1510 7985
rect -1490 7965 -1470 7985
rect -1450 7965 -1430 7985
rect -1410 7965 -1390 7985
rect -1370 7965 -1350 7985
rect -1330 7965 -1310 7985
rect -1290 7965 -1270 7985
rect -1250 7965 -1230 7985
rect -1210 7965 -1190 7985
rect -1170 7965 -1150 7985
rect -1130 7965 -1110 7985
rect -1090 7965 -1070 7985
rect -1050 7965 -1030 7985
rect -1010 7965 -990 7985
rect -970 7965 -950 7985
rect -930 7965 -910 7985
rect -890 7965 -870 7985
rect -850 7965 -830 7985
rect -810 7965 -790 7985
rect -770 7965 -750 7985
rect -730 7965 -710 7985
rect -690 7965 -670 7985
rect -650 7965 -630 7985
rect -610 7965 -590 7985
rect -570 7965 -550 7985
rect -530 7965 -510 7985
rect -490 7965 -470 7985
rect -450 7965 -430 7985
rect -410 7965 -390 7985
rect -370 7965 -350 7985
rect -330 7965 -310 7985
rect -290 7965 -270 7985
rect -250 7965 -230 7985
rect -210 7965 -190 7985
rect -170 7965 -150 7985
rect -130 7965 -110 7985
rect -90 7965 -70 7985
rect -50 7965 -30 7985
rect -10 7965 10 7985
rect 30 7965 50 7985
rect 70 7965 90 7985
rect 110 7965 130 7985
rect 150 7965 170 7985
rect 190 7965 210 7985
rect 230 7965 250 7985
rect 270 7965 290 7985
rect 310 7965 330 7985
rect 350 7965 370 7985
rect 390 7965 410 7985
rect 430 7965 450 7985
rect 470 7965 490 7985
rect 510 7965 525 7985
rect -1975 7955 525 7965
rect 585 7990 600 8010
rect 620 7990 635 8010
rect 585 7970 635 7990
rect -2225 7930 -2175 7950
rect -2225 7910 -2210 7930
rect -2190 7910 -2175 7930
rect -2150 7945 -1995 7955
rect -2150 7925 -2140 7945
rect -2120 7925 -2100 7945
rect -2080 7925 -2060 7945
rect -2040 7925 -2020 7945
rect -2150 7915 -1995 7925
rect 585 7950 600 7970
rect 620 7950 635 7970
rect 585 7930 635 7950
rect -2225 7890 -2175 7910
rect -2225 7870 -2210 7890
rect -2190 7870 -2175 7890
rect -1975 7903 525 7913
rect -1975 7883 -1950 7903
rect -1930 7883 -1910 7903
rect -1890 7883 -1870 7903
rect -1850 7883 -1830 7903
rect -1810 7883 -1790 7903
rect -1770 7883 -1750 7903
rect -1730 7883 -1710 7903
rect -1690 7883 -1670 7903
rect -1650 7883 -1630 7903
rect -1610 7883 -1590 7903
rect -1570 7883 -1550 7903
rect -1530 7883 -1510 7903
rect -1490 7883 -1470 7903
rect -1450 7883 -1430 7903
rect -1410 7883 -1390 7903
rect -1370 7883 -1350 7903
rect -1330 7883 -1310 7903
rect -1290 7883 -1270 7903
rect -1250 7883 -1230 7903
rect -1210 7883 -1190 7903
rect -1170 7883 -1150 7903
rect -1130 7883 -1110 7903
rect -1090 7883 -1070 7903
rect -1050 7883 -1030 7903
rect -1010 7883 -990 7903
rect -970 7883 -950 7903
rect -930 7883 -910 7903
rect -890 7883 -870 7903
rect -850 7883 -830 7903
rect -810 7883 -790 7903
rect -770 7883 -750 7903
rect -730 7883 -710 7903
rect -690 7883 -670 7903
rect -650 7883 -630 7903
rect -610 7883 -590 7903
rect -570 7883 -550 7903
rect -530 7883 -510 7903
rect -490 7883 -470 7903
rect -450 7883 -430 7903
rect -410 7883 -390 7903
rect -370 7883 -350 7903
rect -330 7883 -310 7903
rect -290 7883 -270 7903
rect -250 7883 -230 7903
rect -210 7883 -190 7903
rect -170 7883 -150 7903
rect -130 7883 -110 7903
rect -90 7883 -70 7903
rect -50 7883 -30 7903
rect -10 7883 10 7903
rect 30 7883 50 7903
rect 70 7883 90 7903
rect 110 7883 130 7903
rect 150 7883 170 7903
rect 190 7883 210 7903
rect 230 7883 250 7903
rect 270 7883 290 7903
rect 310 7883 330 7903
rect 350 7883 370 7903
rect 390 7883 410 7903
rect 430 7883 450 7903
rect 470 7883 490 7903
rect 510 7883 525 7903
rect -1975 7873 525 7883
rect 585 7910 600 7930
rect 620 7910 635 7930
rect 585 7890 635 7910
rect 585 7870 600 7890
rect 620 7870 635 7890
rect -2225 7850 -2175 7870
rect -2225 7830 -2210 7850
rect -2190 7830 -2175 7850
rect -2150 7860 -1995 7870
rect -2150 7840 -2140 7860
rect -2120 7840 -2100 7860
rect -2080 7840 -2060 7860
rect -2040 7840 -2020 7860
rect -2150 7830 -1995 7840
rect 585 7850 635 7870
rect -2225 7810 -2175 7830
rect -2225 7790 -2210 7810
rect -2190 7790 -2175 7810
rect -1975 7821 525 7831
rect -1975 7801 -1950 7821
rect -1930 7801 -1910 7821
rect -1890 7801 -1870 7821
rect -1850 7801 -1830 7821
rect -1810 7801 -1790 7821
rect -1770 7801 -1750 7821
rect -1730 7801 -1710 7821
rect -1690 7801 -1670 7821
rect -1650 7801 -1630 7821
rect -1610 7801 -1590 7821
rect -1570 7801 -1550 7821
rect -1530 7801 -1510 7821
rect -1490 7801 -1470 7821
rect -1450 7801 -1430 7821
rect -1410 7801 -1390 7821
rect -1370 7801 -1350 7821
rect -1330 7801 -1310 7821
rect -1290 7801 -1270 7821
rect -1250 7801 -1230 7821
rect -1210 7801 -1190 7821
rect -1170 7801 -1150 7821
rect -1130 7801 -1110 7821
rect -1090 7801 -1070 7821
rect -1050 7801 -1030 7821
rect -1010 7801 -990 7821
rect -970 7801 -950 7821
rect -930 7801 -910 7821
rect -890 7801 -870 7821
rect -850 7801 -830 7821
rect -810 7801 -790 7821
rect -770 7801 -750 7821
rect -730 7801 -710 7821
rect -690 7801 -670 7821
rect -650 7801 -630 7821
rect -610 7801 -590 7821
rect -570 7801 -550 7821
rect -530 7801 -510 7821
rect -490 7801 -470 7821
rect -450 7801 -430 7821
rect -410 7801 -390 7821
rect -370 7801 -350 7821
rect -330 7801 -310 7821
rect -290 7801 -270 7821
rect -250 7801 -230 7821
rect -210 7801 -190 7821
rect -170 7801 -150 7821
rect -130 7801 -110 7821
rect -90 7801 -70 7821
rect -50 7801 -30 7821
rect -10 7801 10 7821
rect 30 7801 50 7821
rect 70 7801 90 7821
rect 110 7801 130 7821
rect 150 7801 170 7821
rect 190 7801 210 7821
rect 230 7801 250 7821
rect 270 7801 290 7821
rect 310 7801 330 7821
rect 350 7801 370 7821
rect 390 7801 410 7821
rect 430 7801 450 7821
rect 470 7801 490 7821
rect 510 7801 525 7821
rect -1975 7791 525 7801
rect 585 7830 600 7850
rect 620 7830 635 7850
rect 585 7810 635 7830
rect 585 7790 600 7810
rect 620 7790 635 7810
rect -2225 7770 -2175 7790
rect -2225 7750 -2210 7770
rect -2190 7750 -2175 7770
rect -2150 7780 -1995 7790
rect -2150 7760 -2140 7780
rect -2120 7760 -2100 7780
rect -2080 7760 -2060 7780
rect -2040 7760 -2020 7780
rect -2150 7750 -1995 7760
rect 585 7770 635 7790
rect 585 7750 600 7770
rect 620 7750 635 7770
rect -2225 7730 -2175 7750
rect -2225 7710 -2210 7730
rect -2190 7710 -2175 7730
rect -1975 7739 525 7749
rect -1975 7719 -1950 7739
rect -1930 7719 -1910 7739
rect -1890 7719 -1870 7739
rect -1850 7719 -1830 7739
rect -1810 7719 -1790 7739
rect -1770 7719 -1750 7739
rect -1730 7719 -1710 7739
rect -1690 7719 -1670 7739
rect -1650 7719 -1630 7739
rect -1610 7719 -1590 7739
rect -1570 7719 -1550 7739
rect -1530 7719 -1510 7739
rect -1490 7719 -1470 7739
rect -1450 7719 -1430 7739
rect -1410 7719 -1390 7739
rect -1370 7719 -1350 7739
rect -1330 7719 -1310 7739
rect -1290 7719 -1270 7739
rect -1250 7719 -1230 7739
rect -1210 7719 -1190 7739
rect -1170 7719 -1150 7739
rect -1130 7719 -1110 7739
rect -1090 7719 -1070 7739
rect -1050 7719 -1030 7739
rect -1010 7719 -990 7739
rect -970 7719 -950 7739
rect -930 7719 -910 7739
rect -890 7719 -870 7739
rect -850 7719 -830 7739
rect -810 7719 -790 7739
rect -770 7719 -750 7739
rect -730 7719 -710 7739
rect -690 7719 -670 7739
rect -650 7719 -630 7739
rect -610 7719 -590 7739
rect -570 7719 -550 7739
rect -530 7719 -510 7739
rect -490 7719 -470 7739
rect -450 7719 -430 7739
rect -410 7719 -390 7739
rect -370 7719 -350 7739
rect -330 7719 -310 7739
rect -290 7719 -270 7739
rect -250 7719 -230 7739
rect -210 7719 -190 7739
rect -170 7719 -150 7739
rect -130 7719 -110 7739
rect -90 7719 -70 7739
rect -50 7719 -30 7739
rect -10 7719 10 7739
rect 30 7719 50 7739
rect 70 7719 90 7739
rect 110 7719 130 7739
rect 150 7719 170 7739
rect 190 7719 210 7739
rect 230 7719 250 7739
rect 270 7719 290 7739
rect 310 7719 330 7739
rect 350 7719 370 7739
rect 390 7719 410 7739
rect 430 7719 450 7739
rect 470 7719 490 7739
rect 510 7719 525 7739
rect -2225 7690 -2175 7710
rect -2225 7670 -2210 7690
rect -2190 7670 -2175 7690
rect -2150 7700 -1995 7710
rect -1975 7709 525 7719
rect 585 7730 635 7750
rect 585 7710 600 7730
rect 620 7710 635 7730
rect -2150 7680 -2140 7700
rect -2120 7680 -2100 7700
rect -2080 7680 -2060 7700
rect -2040 7680 -2020 7700
rect -2150 7670 -1995 7680
rect 585 7690 635 7710
rect 585 7670 600 7690
rect 620 7670 635 7690
rect -2225 7650 -2175 7670
rect -2225 7630 -2210 7650
rect -2190 7630 -2175 7650
rect -2225 7610 -2175 7630
rect -1975 7657 525 7667
rect -1975 7637 -1950 7657
rect -1930 7637 -1910 7657
rect -1890 7637 -1870 7657
rect -1850 7637 -1830 7657
rect -1810 7637 -1790 7657
rect -1770 7637 -1750 7657
rect -1730 7637 -1710 7657
rect -1690 7637 -1670 7657
rect -1650 7637 -1630 7657
rect -1610 7637 -1590 7657
rect -1570 7637 -1550 7657
rect -1530 7637 -1510 7657
rect -1490 7637 -1470 7657
rect -1450 7637 -1430 7657
rect -1410 7637 -1390 7657
rect -1370 7637 -1350 7657
rect -1330 7637 -1310 7657
rect -1290 7637 -1270 7657
rect -1250 7637 -1230 7657
rect -1210 7637 -1190 7657
rect -1170 7637 -1150 7657
rect -1130 7637 -1110 7657
rect -1090 7637 -1070 7657
rect -1050 7637 -1030 7657
rect -1010 7637 -990 7657
rect -970 7637 -950 7657
rect -930 7637 -910 7657
rect -890 7637 -870 7657
rect -850 7637 -830 7657
rect -810 7637 -790 7657
rect -770 7637 -750 7657
rect -730 7637 -710 7657
rect -690 7637 -670 7657
rect -650 7637 -630 7657
rect -610 7637 -590 7657
rect -570 7637 -550 7657
rect -530 7637 -510 7657
rect -490 7637 -470 7657
rect -450 7637 -430 7657
rect -410 7637 -390 7657
rect -370 7637 -350 7657
rect -330 7637 -310 7657
rect -290 7637 -270 7657
rect -250 7637 -230 7657
rect -210 7637 -190 7657
rect -170 7637 -150 7657
rect -130 7637 -110 7657
rect -90 7637 -70 7657
rect -50 7637 -30 7657
rect -10 7637 10 7657
rect 30 7637 50 7657
rect 70 7637 90 7657
rect 110 7637 130 7657
rect 150 7637 170 7657
rect 190 7637 210 7657
rect 230 7637 250 7657
rect 270 7637 290 7657
rect 310 7637 330 7657
rect 350 7637 370 7657
rect 390 7637 410 7657
rect 430 7637 450 7657
rect 470 7637 490 7657
rect 510 7637 525 7657
rect -1975 7627 525 7637
rect 585 7650 635 7670
rect 585 7630 600 7650
rect 620 7630 635 7650
rect -2225 7590 -2210 7610
rect -2190 7590 -2175 7610
rect -2225 7570 -2175 7590
rect -2150 7615 -1995 7625
rect -2150 7595 -2140 7615
rect -2120 7595 -2100 7615
rect -2080 7595 -2060 7615
rect -2040 7595 -2020 7615
rect -2150 7585 -1995 7595
rect 585 7610 635 7630
rect 585 7590 600 7610
rect 620 7590 635 7610
rect -2225 7550 -2210 7570
rect -2190 7550 -2175 7570
rect -2225 7530 -2175 7550
rect -1975 7575 525 7585
rect -1975 7555 -1950 7575
rect -1930 7555 -1910 7575
rect -1890 7555 -1870 7575
rect -1850 7555 -1830 7575
rect -1810 7555 -1790 7575
rect -1770 7555 -1750 7575
rect -1730 7555 -1710 7575
rect -1690 7555 -1670 7575
rect -1650 7555 -1630 7575
rect -1610 7555 -1590 7575
rect -1570 7555 -1550 7575
rect -1530 7555 -1510 7575
rect -1490 7555 -1470 7575
rect -1450 7555 -1430 7575
rect -1410 7555 -1390 7575
rect -1370 7555 -1350 7575
rect -1330 7555 -1310 7575
rect -1290 7555 -1270 7575
rect -1250 7555 -1230 7575
rect -1210 7555 -1190 7575
rect -1170 7555 -1150 7575
rect -1130 7555 -1110 7575
rect -1090 7555 -1070 7575
rect -1050 7555 -1030 7575
rect -1010 7555 -990 7575
rect -970 7555 -950 7575
rect -930 7555 -910 7575
rect -890 7555 -870 7575
rect -850 7555 -830 7575
rect -810 7555 -790 7575
rect -770 7555 -750 7575
rect -730 7555 -710 7575
rect -690 7555 -670 7575
rect -650 7555 -630 7575
rect -610 7555 -590 7575
rect -570 7555 -550 7575
rect -530 7555 -510 7575
rect -490 7555 -470 7575
rect -450 7555 -430 7575
rect -410 7555 -390 7575
rect -370 7555 -350 7575
rect -330 7555 -310 7575
rect -290 7555 -270 7575
rect -250 7555 -230 7575
rect -210 7555 -190 7575
rect -170 7555 -150 7575
rect -130 7555 -110 7575
rect -90 7555 -70 7575
rect -50 7555 -30 7575
rect -10 7555 10 7575
rect 30 7555 50 7575
rect 70 7555 90 7575
rect 110 7555 130 7575
rect 150 7555 170 7575
rect 190 7555 210 7575
rect 230 7555 250 7575
rect 270 7555 290 7575
rect 310 7555 330 7575
rect 350 7555 370 7575
rect 390 7555 410 7575
rect 430 7555 450 7575
rect 470 7555 490 7575
rect 510 7555 525 7575
rect -1975 7545 525 7555
rect 585 7570 635 7590
rect 585 7550 600 7570
rect 620 7550 635 7570
rect -2225 7510 -2210 7530
rect -2190 7510 -2175 7530
rect -2225 7490 -2175 7510
rect -2150 7535 -1995 7545
rect -2150 7515 -2140 7535
rect -2120 7515 -2100 7535
rect -2080 7515 -2060 7535
rect -2040 7515 -2020 7535
rect -2150 7505 -1995 7515
rect 585 7530 635 7550
rect 585 7510 600 7530
rect 620 7510 635 7530
rect -2225 7470 -2210 7490
rect -2190 7470 -2175 7490
rect -2225 7450 -2175 7470
rect -1975 7493 525 7503
rect -1975 7473 -1950 7493
rect -1930 7473 -1910 7493
rect -1890 7473 -1870 7493
rect -1850 7473 -1830 7493
rect -1810 7473 -1790 7493
rect -1770 7473 -1750 7493
rect -1730 7473 -1710 7493
rect -1690 7473 -1670 7493
rect -1650 7473 -1630 7493
rect -1610 7473 -1590 7493
rect -1570 7473 -1550 7493
rect -1530 7473 -1510 7493
rect -1490 7473 -1470 7493
rect -1450 7473 -1430 7493
rect -1410 7473 -1390 7493
rect -1370 7473 -1350 7493
rect -1330 7473 -1310 7493
rect -1290 7473 -1270 7493
rect -1250 7473 -1230 7493
rect -1210 7473 -1190 7493
rect -1170 7473 -1150 7493
rect -1130 7473 -1110 7493
rect -1090 7473 -1070 7493
rect -1050 7473 -1030 7493
rect -1010 7473 -990 7493
rect -970 7473 -950 7493
rect -930 7473 -910 7493
rect -890 7473 -870 7493
rect -850 7473 -830 7493
rect -810 7473 -790 7493
rect -770 7473 -750 7493
rect -730 7473 -710 7493
rect -690 7473 -670 7493
rect -650 7473 -630 7493
rect -610 7473 -590 7493
rect -570 7473 -550 7493
rect -530 7473 -510 7493
rect -490 7473 -470 7493
rect -450 7473 -430 7493
rect -410 7473 -390 7493
rect -370 7473 -350 7493
rect -330 7473 -310 7493
rect -290 7473 -270 7493
rect -250 7473 -230 7493
rect -210 7473 -190 7493
rect -170 7473 -150 7493
rect -130 7473 -110 7493
rect -90 7473 -70 7493
rect -50 7473 -30 7493
rect -10 7473 10 7493
rect 30 7473 50 7493
rect 70 7473 90 7493
rect 110 7473 130 7493
rect 150 7473 170 7493
rect 190 7473 210 7493
rect 230 7473 250 7493
rect 270 7473 290 7493
rect 310 7473 330 7493
rect 350 7473 370 7493
rect 390 7473 410 7493
rect 430 7473 450 7493
rect 470 7473 490 7493
rect 510 7473 525 7493
rect -1975 7463 525 7473
rect 585 7490 635 7510
rect 585 7470 600 7490
rect 620 7470 635 7490
rect -2225 7430 -2210 7450
rect -2190 7430 -2175 7450
rect -2225 7410 -2175 7430
rect -2150 7450 -1995 7460
rect -2150 7430 -2140 7450
rect -2120 7430 -2100 7450
rect -2080 7430 -2060 7450
rect -2040 7430 -2020 7450
rect -2150 7420 -1995 7430
rect 585 7450 635 7470
rect 585 7430 600 7450
rect 620 7430 635 7450
rect -2225 7390 -2210 7410
rect -2190 7390 -2175 7410
rect -2225 7370 -2175 7390
rect -1975 7411 525 7421
rect -1975 7391 -1950 7411
rect -1930 7391 -1910 7411
rect -1890 7391 -1870 7411
rect -1850 7391 -1830 7411
rect -1810 7391 -1790 7411
rect -1770 7391 -1750 7411
rect -1730 7391 -1710 7411
rect -1690 7391 -1670 7411
rect -1650 7391 -1630 7411
rect -1610 7391 -1590 7411
rect -1570 7391 -1550 7411
rect -1530 7391 -1510 7411
rect -1490 7391 -1470 7411
rect -1450 7391 -1430 7411
rect -1410 7391 -1390 7411
rect -1370 7391 -1350 7411
rect -1330 7391 -1310 7411
rect -1290 7391 -1270 7411
rect -1250 7391 -1230 7411
rect -1210 7391 -1190 7411
rect -1170 7391 -1150 7411
rect -1130 7391 -1110 7411
rect -1090 7391 -1070 7411
rect -1050 7391 -1030 7411
rect -1010 7391 -990 7411
rect -970 7391 -950 7411
rect -930 7391 -910 7411
rect -890 7391 -870 7411
rect -850 7391 -830 7411
rect -810 7391 -790 7411
rect -770 7391 -750 7411
rect -730 7391 -710 7411
rect -690 7391 -670 7411
rect -650 7391 -630 7411
rect -610 7391 -590 7411
rect -570 7391 -550 7411
rect -530 7391 -510 7411
rect -490 7391 -470 7411
rect -450 7391 -430 7411
rect -410 7391 -390 7411
rect -370 7391 -350 7411
rect -330 7391 -310 7411
rect -290 7391 -270 7411
rect -250 7391 -230 7411
rect -210 7391 -190 7411
rect -170 7391 -150 7411
rect -130 7391 -110 7411
rect -90 7391 -70 7411
rect -50 7391 -30 7411
rect -10 7391 10 7411
rect 30 7391 50 7411
rect 70 7391 90 7411
rect 110 7391 130 7411
rect 150 7391 170 7411
rect 190 7391 210 7411
rect 230 7391 250 7411
rect 270 7391 290 7411
rect 310 7391 330 7411
rect 350 7391 370 7411
rect 390 7391 410 7411
rect 430 7391 450 7411
rect 470 7391 490 7411
rect 510 7391 525 7411
rect -1975 7381 525 7391
rect 585 7410 635 7430
rect 585 7390 600 7410
rect 620 7390 635 7410
rect -2225 7350 -2210 7370
rect -2190 7350 -2175 7370
rect -2225 7330 -2175 7350
rect -2150 7370 -1995 7380
rect -2150 7350 -2140 7370
rect -2120 7350 -2100 7370
rect -2080 7350 -2060 7370
rect -2040 7350 -2020 7370
rect -2150 7340 -1995 7350
rect 585 7370 635 7390
rect 585 7350 600 7370
rect 620 7350 635 7370
rect -2225 7310 -2210 7330
rect -2190 7310 -2175 7330
rect -2225 7290 -2175 7310
rect -1975 7329 525 7339
rect -1975 7309 -1950 7329
rect -1930 7309 -1910 7329
rect -1890 7309 -1870 7329
rect -1850 7309 -1830 7329
rect -1810 7309 -1790 7329
rect -1770 7309 -1750 7329
rect -1730 7309 -1710 7329
rect -1690 7309 -1670 7329
rect -1650 7309 -1630 7329
rect -1610 7309 -1590 7329
rect -1570 7309 -1550 7329
rect -1530 7309 -1510 7329
rect -1490 7309 -1470 7329
rect -1450 7309 -1430 7329
rect -1410 7309 -1390 7329
rect -1370 7309 -1350 7329
rect -1330 7309 -1310 7329
rect -1290 7309 -1270 7329
rect -1250 7309 -1230 7329
rect -1210 7309 -1190 7329
rect -1170 7309 -1150 7329
rect -1130 7309 -1110 7329
rect -1090 7309 -1070 7329
rect -1050 7309 -1030 7329
rect -1010 7309 -990 7329
rect -970 7309 -950 7329
rect -930 7309 -910 7329
rect -890 7309 -870 7329
rect -850 7309 -830 7329
rect -810 7309 -790 7329
rect -770 7309 -750 7329
rect -730 7309 -710 7329
rect -690 7309 -670 7329
rect -650 7309 -630 7329
rect -610 7309 -590 7329
rect -570 7309 -550 7329
rect -530 7309 -510 7329
rect -490 7309 -470 7329
rect -450 7309 -430 7329
rect -410 7309 -390 7329
rect -370 7309 -350 7329
rect -330 7309 -310 7329
rect -290 7309 -270 7329
rect -250 7309 -230 7329
rect -210 7309 -190 7329
rect -170 7309 -150 7329
rect -130 7309 -110 7329
rect -90 7309 -70 7329
rect -50 7309 -30 7329
rect -10 7309 10 7329
rect 30 7309 50 7329
rect 70 7309 90 7329
rect 110 7309 130 7329
rect 150 7309 170 7329
rect 190 7309 210 7329
rect 230 7309 250 7329
rect 270 7309 290 7329
rect 310 7309 330 7329
rect 350 7309 370 7329
rect 390 7309 410 7329
rect 430 7309 450 7329
rect 470 7309 490 7329
rect 510 7309 525 7329
rect -2225 7270 -2210 7290
rect -2190 7270 -2175 7290
rect -2225 7250 -2175 7270
rect -2150 7290 -1995 7300
rect -1975 7299 525 7309
rect 585 7330 635 7350
rect 585 7310 600 7330
rect 620 7310 635 7330
rect -2150 7270 -2140 7290
rect -2120 7270 -2100 7290
rect -2080 7270 -2060 7290
rect -2040 7270 -2020 7290
rect -2150 7260 -1995 7270
rect 585 7290 635 7310
rect 585 7270 600 7290
rect 620 7270 635 7290
rect -2225 7230 -2210 7250
rect -2190 7230 -2175 7250
rect -2225 7210 -2175 7230
rect -1975 7247 525 7257
rect -1975 7227 -1950 7247
rect -1930 7227 -1910 7247
rect -1890 7227 -1870 7247
rect -1850 7227 -1830 7247
rect -1810 7227 -1790 7247
rect -1770 7227 -1750 7247
rect -1730 7227 -1710 7247
rect -1690 7227 -1670 7247
rect -1650 7227 -1630 7247
rect -1610 7227 -1590 7247
rect -1570 7227 -1550 7247
rect -1530 7227 -1510 7247
rect -1490 7227 -1470 7247
rect -1450 7227 -1430 7247
rect -1410 7227 -1390 7247
rect -1370 7227 -1350 7247
rect -1330 7227 -1310 7247
rect -1290 7227 -1270 7247
rect -1250 7227 -1230 7247
rect -1210 7227 -1190 7247
rect -1170 7227 -1150 7247
rect -1130 7227 -1110 7247
rect -1090 7227 -1070 7247
rect -1050 7227 -1030 7247
rect -1010 7227 -990 7247
rect -970 7227 -950 7247
rect -930 7227 -910 7247
rect -890 7227 -870 7247
rect -850 7227 -830 7247
rect -810 7227 -790 7247
rect -770 7227 -750 7247
rect -730 7227 -710 7247
rect -690 7227 -670 7247
rect -650 7227 -630 7247
rect -610 7227 -590 7247
rect -570 7227 -550 7247
rect -530 7227 -510 7247
rect -490 7227 -470 7247
rect -450 7227 -430 7247
rect -410 7227 -390 7247
rect -370 7227 -350 7247
rect -330 7227 -310 7247
rect -290 7227 -270 7247
rect -250 7227 -230 7247
rect -210 7227 -190 7247
rect -170 7227 -150 7247
rect -130 7227 -110 7247
rect -90 7227 -70 7247
rect -50 7227 -30 7247
rect -10 7227 10 7247
rect 30 7227 50 7247
rect 70 7227 90 7247
rect 110 7227 130 7247
rect 150 7227 170 7247
rect 190 7227 210 7247
rect 230 7227 250 7247
rect 270 7227 290 7247
rect 310 7227 330 7247
rect 350 7227 370 7247
rect 390 7227 410 7247
rect 430 7227 450 7247
rect 470 7227 490 7247
rect 510 7227 525 7247
rect -1975 7217 525 7227
rect 585 7250 635 7270
rect 585 7230 600 7250
rect 620 7230 635 7250
rect -2225 7190 -2210 7210
rect -2190 7190 -2175 7210
rect -2225 7170 -2175 7190
rect -2150 7205 -1995 7215
rect -2150 7185 -2140 7205
rect -2120 7185 -2100 7205
rect -2080 7185 -2060 7205
rect -2040 7185 -2020 7205
rect -2150 7175 -1995 7185
rect 585 7210 635 7230
rect 585 7190 600 7210
rect 620 7190 635 7210
rect -2225 7150 -2210 7170
rect -2190 7150 -2175 7170
rect -2225 7130 -2175 7150
rect -1975 7165 525 7175
rect -1975 7145 -1950 7165
rect -1930 7145 -1910 7165
rect -1890 7145 -1870 7165
rect -1850 7145 -1830 7165
rect -1810 7145 -1790 7165
rect -1770 7145 -1750 7165
rect -1730 7145 -1710 7165
rect -1690 7145 -1670 7165
rect -1650 7145 -1630 7165
rect -1610 7145 -1590 7165
rect -1570 7145 -1550 7165
rect -1530 7145 -1510 7165
rect -1490 7145 -1470 7165
rect -1450 7145 -1430 7165
rect -1410 7145 -1390 7165
rect -1370 7145 -1350 7165
rect -1330 7145 -1310 7165
rect -1290 7145 -1270 7165
rect -1250 7145 -1230 7165
rect -1210 7145 -1190 7165
rect -1170 7145 -1150 7165
rect -1130 7145 -1110 7165
rect -1090 7145 -1070 7165
rect -1050 7145 -1030 7165
rect -1010 7145 -990 7165
rect -970 7145 -950 7165
rect -930 7145 -910 7165
rect -890 7145 -870 7165
rect -850 7145 -830 7165
rect -810 7145 -790 7165
rect -770 7145 -750 7165
rect -730 7145 -710 7165
rect -690 7145 -670 7165
rect -650 7145 -630 7165
rect -610 7145 -590 7165
rect -570 7145 -550 7165
rect -530 7145 -510 7165
rect -490 7145 -470 7165
rect -450 7145 -430 7165
rect -410 7145 -390 7165
rect -370 7145 -350 7165
rect -330 7145 -310 7165
rect -290 7145 -270 7165
rect -250 7145 -230 7165
rect -210 7145 -190 7165
rect -170 7145 -150 7165
rect -130 7145 -110 7165
rect -90 7145 -70 7165
rect -50 7145 -30 7165
rect -10 7145 10 7165
rect 30 7145 50 7165
rect 70 7145 90 7165
rect 110 7145 130 7165
rect 150 7145 170 7165
rect 190 7145 210 7165
rect 230 7145 250 7165
rect 270 7145 290 7165
rect 310 7145 330 7165
rect 350 7145 370 7165
rect 390 7145 410 7165
rect 430 7145 450 7165
rect 470 7145 490 7165
rect 510 7145 525 7165
rect -1975 7135 525 7145
rect 585 7170 635 7190
rect 585 7150 600 7170
rect 620 7150 635 7170
rect -2225 7110 -2210 7130
rect -2190 7110 -2175 7130
rect -2225 7090 -2175 7110
rect -2150 7125 -1995 7135
rect -2150 7105 -2140 7125
rect -2120 7105 -2100 7125
rect -2080 7105 -2060 7125
rect -2040 7105 -2020 7125
rect -2150 7095 -1995 7105
rect 585 7130 635 7150
rect 585 7110 600 7130
rect 620 7110 635 7130
rect -2225 7070 -2210 7090
rect -2190 7070 -2175 7090
rect -2225 7050 -2175 7070
rect -1975 7083 525 7093
rect -1975 7063 -1950 7083
rect -1930 7063 -1910 7083
rect -1890 7063 -1870 7083
rect -1850 7063 -1830 7083
rect -1810 7063 -1790 7083
rect -1770 7063 -1750 7083
rect -1730 7063 -1710 7083
rect -1690 7063 -1670 7083
rect -1650 7063 -1630 7083
rect -1610 7063 -1590 7083
rect -1570 7063 -1550 7083
rect -1530 7063 -1510 7083
rect -1490 7063 -1470 7083
rect -1450 7063 -1430 7083
rect -1410 7063 -1390 7083
rect -1370 7063 -1350 7083
rect -1330 7063 -1310 7083
rect -1290 7063 -1270 7083
rect -1250 7063 -1230 7083
rect -1210 7063 -1190 7083
rect -1170 7063 -1150 7083
rect -1130 7063 -1110 7083
rect -1090 7063 -1070 7083
rect -1050 7063 -1030 7083
rect -1010 7063 -990 7083
rect -970 7063 -950 7083
rect -930 7063 -910 7083
rect -890 7063 -870 7083
rect -850 7063 -830 7083
rect -810 7063 -790 7083
rect -770 7063 -750 7083
rect -730 7063 -710 7083
rect -690 7063 -670 7083
rect -650 7063 -630 7083
rect -610 7063 -590 7083
rect -570 7063 -550 7083
rect -530 7063 -510 7083
rect -490 7063 -470 7083
rect -450 7063 -430 7083
rect -410 7063 -390 7083
rect -370 7063 -350 7083
rect -330 7063 -310 7083
rect -290 7063 -270 7083
rect -250 7063 -230 7083
rect -210 7063 -190 7083
rect -170 7063 -150 7083
rect -130 7063 -110 7083
rect -90 7063 -70 7083
rect -50 7063 -30 7083
rect -10 7063 10 7083
rect 30 7063 50 7083
rect 70 7063 90 7083
rect 110 7063 130 7083
rect 150 7063 170 7083
rect 190 7063 210 7083
rect 230 7063 250 7083
rect 270 7063 290 7083
rect 310 7063 330 7083
rect 350 7063 370 7083
rect 390 7063 410 7083
rect 430 7063 450 7083
rect 470 7063 490 7083
rect 510 7063 525 7083
rect -1975 7053 525 7063
rect 585 7090 635 7110
rect 585 7070 600 7090
rect 620 7070 635 7090
rect 585 7050 635 7070
rect -2225 7030 -2210 7050
rect -2190 7030 -2175 7050
rect -2225 7010 -2175 7030
rect -2150 7040 -1995 7050
rect -2150 7020 -2140 7040
rect -2120 7020 -2100 7040
rect -2080 7020 -2060 7040
rect -2040 7020 -2020 7040
rect -2150 7010 -1995 7020
rect 585 7030 600 7050
rect 620 7030 635 7050
rect -2225 6990 -2210 7010
rect -2190 6990 -2175 7010
rect -2225 6970 -2175 6990
rect -1975 7001 525 7011
rect -1975 6981 -1950 7001
rect -1930 6981 -1910 7001
rect -1890 6981 -1870 7001
rect -1850 6981 -1830 7001
rect -1810 6981 -1790 7001
rect -1770 6981 -1750 7001
rect -1730 6981 -1710 7001
rect -1690 6981 -1670 7001
rect -1650 6981 -1630 7001
rect -1610 6981 -1590 7001
rect -1570 6981 -1550 7001
rect -1530 6981 -1510 7001
rect -1490 6981 -1470 7001
rect -1450 6981 -1430 7001
rect -1410 6981 -1390 7001
rect -1370 6981 -1350 7001
rect -1330 6981 -1310 7001
rect -1290 6981 -1270 7001
rect -1250 6981 -1230 7001
rect -1210 6981 -1190 7001
rect -1170 6981 -1150 7001
rect -1130 6981 -1110 7001
rect -1090 6981 -1070 7001
rect -1050 6981 -1030 7001
rect -1010 6981 -990 7001
rect -970 6981 -950 7001
rect -930 6981 -910 7001
rect -890 6981 -870 7001
rect -850 6981 -830 7001
rect -810 6981 -790 7001
rect -770 6981 -750 7001
rect -730 6981 -710 7001
rect -690 6981 -670 7001
rect -650 6981 -630 7001
rect -610 6981 -590 7001
rect -570 6981 -550 7001
rect -530 6981 -510 7001
rect -490 6981 -470 7001
rect -450 6981 -430 7001
rect -410 6981 -390 7001
rect -370 6981 -350 7001
rect -330 6981 -310 7001
rect -290 6981 -270 7001
rect -250 6981 -230 7001
rect -210 6981 -190 7001
rect -170 6981 -150 7001
rect -130 6981 -110 7001
rect -90 6981 -70 7001
rect -50 6981 -30 7001
rect -10 6981 10 7001
rect 30 6981 50 7001
rect 70 6981 90 7001
rect 110 6981 130 7001
rect 150 6981 170 7001
rect 190 6981 210 7001
rect 230 6981 250 7001
rect 270 6981 290 7001
rect 310 6981 330 7001
rect 350 6981 370 7001
rect 390 6981 410 7001
rect 430 6981 450 7001
rect 470 6981 490 7001
rect 510 6981 525 7001
rect -1975 6971 525 6981
rect 585 7010 635 7030
rect 585 6990 600 7010
rect 620 6990 635 7010
rect 585 6970 635 6990
rect -2225 6950 -2210 6970
rect -2190 6950 -2175 6970
rect -2225 6930 -2175 6950
rect -2150 6960 -1995 6970
rect -2150 6940 -2140 6960
rect -2120 6940 -2100 6960
rect -2080 6940 -2060 6960
rect -2040 6940 -2020 6960
rect -2150 6930 -1995 6940
rect 585 6950 600 6970
rect 620 6950 635 6970
rect 585 6930 635 6950
rect -2225 6910 -2210 6930
rect -2190 6910 -2175 6930
rect -2225 6890 -2175 6910
rect -1975 6919 525 6929
rect -1975 6899 -1950 6919
rect -1930 6899 -1910 6919
rect -1890 6899 -1870 6919
rect -1850 6899 -1830 6919
rect -1810 6899 -1790 6919
rect -1770 6899 -1750 6919
rect -1730 6899 -1710 6919
rect -1690 6899 -1670 6919
rect -1650 6899 -1630 6919
rect -1610 6899 -1590 6919
rect -1570 6899 -1550 6919
rect -1530 6899 -1510 6919
rect -1490 6899 -1470 6919
rect -1450 6899 -1430 6919
rect -1410 6899 -1390 6919
rect -1370 6899 -1350 6919
rect -1330 6899 -1310 6919
rect -1290 6899 -1270 6919
rect -1250 6899 -1230 6919
rect -1210 6899 -1190 6919
rect -1170 6899 -1150 6919
rect -1130 6899 -1110 6919
rect -1090 6899 -1070 6919
rect -1050 6899 -1030 6919
rect -1010 6899 -990 6919
rect -970 6899 -950 6919
rect -930 6899 -910 6919
rect -890 6899 -870 6919
rect -850 6899 -830 6919
rect -810 6899 -790 6919
rect -770 6899 -750 6919
rect -730 6899 -710 6919
rect -690 6899 -670 6919
rect -650 6899 -630 6919
rect -610 6899 -590 6919
rect -570 6899 -550 6919
rect -530 6899 -510 6919
rect -490 6899 -470 6919
rect -450 6899 -430 6919
rect -410 6899 -390 6919
rect -370 6899 -350 6919
rect -330 6899 -310 6919
rect -290 6899 -270 6919
rect -250 6899 -230 6919
rect -210 6899 -190 6919
rect -170 6899 -150 6919
rect -130 6899 -110 6919
rect -90 6899 -70 6919
rect -50 6899 -30 6919
rect -10 6899 10 6919
rect 30 6899 50 6919
rect 70 6899 90 6919
rect 110 6899 130 6919
rect 150 6899 170 6919
rect 190 6899 210 6919
rect 230 6899 250 6919
rect 270 6899 290 6919
rect 310 6899 330 6919
rect 350 6899 370 6919
rect 390 6899 410 6919
rect 430 6899 450 6919
rect 470 6899 490 6919
rect 510 6899 525 6919
rect -2225 6870 -2210 6890
rect -2190 6870 -2175 6890
rect -2225 6850 -2175 6870
rect -2150 6880 -1995 6890
rect -1975 6889 525 6899
rect 585 6910 600 6930
rect 620 6910 635 6930
rect 585 6890 635 6910
rect -2150 6860 -2140 6880
rect -2120 6860 -2100 6880
rect -2080 6860 -2060 6880
rect -2040 6860 -2020 6880
rect -2150 6850 -1995 6860
rect 585 6870 600 6890
rect 620 6870 635 6890
rect 585 6850 635 6870
rect -2225 6830 -2210 6850
rect -2190 6830 -2175 6850
rect -2225 6810 -2175 6830
rect -2225 6790 -2210 6810
rect -2190 6790 -2175 6810
rect -1975 6837 525 6847
rect -1975 6817 -1950 6837
rect -1930 6817 -1910 6837
rect -1890 6817 -1870 6837
rect -1850 6817 -1830 6837
rect -1810 6817 -1790 6837
rect -1770 6817 -1750 6837
rect -1730 6817 -1710 6837
rect -1690 6817 -1670 6837
rect -1650 6817 -1630 6837
rect -1610 6817 -1590 6837
rect -1570 6817 -1550 6837
rect -1530 6817 -1510 6837
rect -1490 6817 -1470 6837
rect -1450 6817 -1430 6837
rect -1410 6817 -1390 6837
rect -1370 6817 -1350 6837
rect -1330 6817 -1310 6837
rect -1290 6817 -1270 6837
rect -1250 6817 -1230 6837
rect -1210 6817 -1190 6837
rect -1170 6817 -1150 6837
rect -1130 6817 -1110 6837
rect -1090 6817 -1070 6837
rect -1050 6817 -1030 6837
rect -1010 6817 -990 6837
rect -970 6817 -950 6837
rect -930 6817 -910 6837
rect -890 6817 -870 6837
rect -850 6817 -830 6837
rect -810 6817 -790 6837
rect -770 6817 -750 6837
rect -730 6817 -710 6837
rect -690 6817 -670 6837
rect -650 6817 -630 6837
rect -610 6817 -590 6837
rect -570 6817 -550 6837
rect -530 6817 -510 6837
rect -490 6817 -470 6837
rect -450 6817 -430 6837
rect -410 6817 -390 6837
rect -370 6817 -350 6837
rect -330 6817 -310 6837
rect -290 6817 -270 6837
rect -250 6817 -230 6837
rect -210 6817 -190 6837
rect -170 6817 -150 6837
rect -130 6817 -110 6837
rect -90 6817 -70 6837
rect -50 6817 -30 6837
rect -10 6817 10 6837
rect 30 6817 50 6837
rect 70 6817 90 6837
rect 110 6817 130 6837
rect 150 6817 170 6837
rect 190 6817 210 6837
rect 230 6817 250 6837
rect 270 6817 290 6837
rect 310 6817 330 6837
rect 350 6817 370 6837
rect 390 6817 410 6837
rect 430 6817 450 6837
rect 470 6817 490 6837
rect 510 6817 525 6837
rect -1975 6807 525 6817
rect 585 6830 600 6850
rect 620 6830 635 6850
rect 585 6810 635 6830
rect -2225 6770 -2175 6790
rect -2225 6750 -2210 6770
rect -2190 6750 -2175 6770
rect -2150 6795 -1995 6805
rect -2150 6775 -2140 6795
rect -2120 6775 -2100 6795
rect -2080 6775 -2060 6795
rect -2040 6775 -2020 6795
rect -2150 6765 -1995 6775
rect 585 6790 600 6810
rect 620 6790 635 6810
rect 585 6770 635 6790
rect -2225 6730 -2175 6750
rect -2225 6710 -2210 6730
rect -2190 6710 -2175 6730
rect -1975 6755 525 6765
rect -1975 6735 -1950 6755
rect -1930 6735 -1910 6755
rect -1890 6735 -1870 6755
rect -1850 6735 -1830 6755
rect -1810 6735 -1790 6755
rect -1770 6735 -1750 6755
rect -1730 6735 -1710 6755
rect -1690 6735 -1670 6755
rect -1650 6735 -1630 6755
rect -1610 6735 -1590 6755
rect -1570 6735 -1550 6755
rect -1530 6735 -1510 6755
rect -1490 6735 -1470 6755
rect -1450 6735 -1430 6755
rect -1410 6735 -1390 6755
rect -1370 6735 -1350 6755
rect -1330 6735 -1310 6755
rect -1290 6735 -1270 6755
rect -1250 6735 -1230 6755
rect -1210 6735 -1190 6755
rect -1170 6735 -1150 6755
rect -1130 6735 -1110 6755
rect -1090 6735 -1070 6755
rect -1050 6735 -1030 6755
rect -1010 6735 -990 6755
rect -970 6735 -950 6755
rect -930 6735 -910 6755
rect -890 6735 -870 6755
rect -850 6735 -830 6755
rect -810 6735 -790 6755
rect -770 6735 -750 6755
rect -730 6735 -710 6755
rect -690 6735 -670 6755
rect -650 6735 -630 6755
rect -610 6735 -590 6755
rect -570 6735 -550 6755
rect -530 6735 -510 6755
rect -490 6735 -470 6755
rect -450 6735 -430 6755
rect -410 6735 -390 6755
rect -370 6735 -350 6755
rect -330 6735 -310 6755
rect -290 6735 -270 6755
rect -250 6735 -230 6755
rect -210 6735 -190 6755
rect -170 6735 -150 6755
rect -130 6735 -110 6755
rect -90 6735 -70 6755
rect -50 6735 -30 6755
rect -10 6735 10 6755
rect 30 6735 50 6755
rect 70 6735 90 6755
rect 110 6735 130 6755
rect 150 6735 170 6755
rect 190 6735 210 6755
rect 230 6735 250 6755
rect 270 6735 290 6755
rect 310 6735 330 6755
rect 350 6735 370 6755
rect 390 6735 410 6755
rect 430 6735 450 6755
rect 470 6735 490 6755
rect 510 6735 525 6755
rect -1975 6725 525 6735
rect 585 6750 600 6770
rect 620 6750 635 6770
rect 585 6730 635 6750
rect -2225 6690 -2175 6710
rect -2225 6670 -2210 6690
rect -2190 6670 -2175 6690
rect -2150 6715 -1995 6725
rect -2150 6695 -2140 6715
rect -2120 6695 -2100 6715
rect -2080 6695 -2060 6715
rect -2040 6695 -2020 6715
rect -2150 6685 -1995 6695
rect 585 6710 600 6730
rect 620 6710 635 6730
rect 585 6690 635 6710
rect -2225 6650 -2175 6670
rect -2225 6630 -2210 6650
rect -2190 6630 -2175 6650
rect -1975 6673 525 6683
rect -1975 6653 -1950 6673
rect -1930 6653 -1910 6673
rect -1890 6653 -1870 6673
rect -1850 6653 -1830 6673
rect -1810 6653 -1790 6673
rect -1770 6653 -1750 6673
rect -1730 6653 -1710 6673
rect -1690 6653 -1670 6673
rect -1650 6653 -1630 6673
rect -1610 6653 -1590 6673
rect -1570 6653 -1550 6673
rect -1530 6653 -1510 6673
rect -1490 6653 -1470 6673
rect -1450 6653 -1430 6673
rect -1410 6653 -1390 6673
rect -1370 6653 -1350 6673
rect -1330 6653 -1310 6673
rect -1290 6653 -1270 6673
rect -1250 6653 -1230 6673
rect -1210 6653 -1190 6673
rect -1170 6653 -1150 6673
rect -1130 6653 -1110 6673
rect -1090 6653 -1070 6673
rect -1050 6653 -1030 6673
rect -1010 6653 -990 6673
rect -970 6653 -950 6673
rect -930 6653 -910 6673
rect -890 6653 -870 6673
rect -850 6653 -830 6673
rect -810 6653 -790 6673
rect -770 6653 -750 6673
rect -730 6653 -710 6673
rect -690 6653 -670 6673
rect -650 6653 -630 6673
rect -610 6653 -590 6673
rect -570 6653 -550 6673
rect -530 6653 -510 6673
rect -490 6653 -470 6673
rect -450 6653 -430 6673
rect -410 6653 -390 6673
rect -370 6653 -350 6673
rect -330 6653 -310 6673
rect -290 6653 -270 6673
rect -250 6653 -230 6673
rect -210 6653 -190 6673
rect -170 6653 -150 6673
rect -130 6653 -110 6673
rect -90 6653 -70 6673
rect -50 6653 -30 6673
rect -10 6653 10 6673
rect 30 6653 50 6673
rect 70 6653 90 6673
rect 110 6653 130 6673
rect 150 6653 170 6673
rect 190 6653 210 6673
rect 230 6653 250 6673
rect 270 6653 290 6673
rect 310 6653 330 6673
rect 350 6653 370 6673
rect 390 6653 410 6673
rect 430 6653 450 6673
rect 470 6653 490 6673
rect 510 6653 525 6673
rect -2225 6610 -2175 6630
rect -2225 6590 -2210 6610
rect -2190 6590 -2175 6610
rect -2150 6635 -1995 6645
rect -1975 6643 525 6653
rect 585 6670 600 6690
rect 620 6670 635 6690
rect 585 6650 635 6670
rect -2150 6615 -2140 6635
rect -2120 6615 -2100 6635
rect -2080 6615 -2060 6635
rect -2040 6615 -2020 6635
rect -2150 6605 -1995 6615
rect 585 6630 600 6650
rect 620 6630 635 6650
rect 585 6610 635 6630
rect -2225 6570 -2175 6590
rect -2225 6550 -2210 6570
rect -2190 6550 -2175 6570
rect -1975 6591 525 6601
rect -1975 6571 -1950 6591
rect -1930 6571 -1910 6591
rect -1890 6571 -1870 6591
rect -1850 6571 -1830 6591
rect -1810 6571 -1790 6591
rect -1770 6571 -1750 6591
rect -1730 6571 -1710 6591
rect -1690 6571 -1670 6591
rect -1650 6571 -1630 6591
rect -1610 6571 -1590 6591
rect -1570 6571 -1550 6591
rect -1530 6571 -1510 6591
rect -1490 6571 -1470 6591
rect -1450 6571 -1430 6591
rect -1410 6571 -1390 6591
rect -1370 6571 -1350 6591
rect -1330 6571 -1310 6591
rect -1290 6571 -1270 6591
rect -1250 6571 -1230 6591
rect -1210 6571 -1190 6591
rect -1170 6571 -1150 6591
rect -1130 6571 -1110 6591
rect -1090 6571 -1070 6591
rect -1050 6571 -1030 6591
rect -1010 6571 -990 6591
rect -970 6571 -950 6591
rect -930 6571 -910 6591
rect -890 6571 -870 6591
rect -850 6571 -830 6591
rect -810 6571 -790 6591
rect -770 6571 -750 6591
rect -730 6571 -710 6591
rect -690 6571 -670 6591
rect -650 6571 -630 6591
rect -610 6571 -590 6591
rect -570 6571 -550 6591
rect -530 6571 -510 6591
rect -490 6571 -470 6591
rect -450 6571 -430 6591
rect -410 6571 -390 6591
rect -370 6571 -350 6591
rect -330 6571 -310 6591
rect -290 6571 -270 6591
rect -250 6571 -230 6591
rect -210 6571 -190 6591
rect -170 6571 -150 6591
rect -130 6571 -110 6591
rect -90 6571 -70 6591
rect -50 6571 -30 6591
rect -10 6571 10 6591
rect 30 6571 50 6591
rect 70 6571 90 6591
rect 110 6571 130 6591
rect 150 6571 170 6591
rect 190 6571 210 6591
rect 230 6571 250 6591
rect 270 6571 290 6591
rect 310 6571 330 6591
rect 350 6571 370 6591
rect 390 6571 410 6591
rect 430 6571 450 6591
rect 470 6571 490 6591
rect 510 6571 525 6591
rect -1975 6561 525 6571
rect 585 6590 600 6610
rect 620 6590 635 6610
rect 585 6570 635 6590
rect -2225 6530 -2175 6550
rect -2225 6510 -2210 6530
rect -2190 6510 -2175 6530
rect -2150 6550 -1995 6560
rect -2150 6530 -2140 6550
rect -2120 6530 -2100 6550
rect -2080 6530 -2060 6550
rect -2040 6530 -2020 6550
rect -2150 6520 -1995 6530
rect 585 6550 600 6570
rect 620 6550 635 6570
rect 585 6530 635 6550
rect -2225 6490 -2175 6510
rect -2225 6470 -2210 6490
rect -2190 6470 -2175 6490
rect -1975 6509 525 6519
rect -1975 6489 -1950 6509
rect -1930 6489 -1910 6509
rect -1890 6489 -1870 6509
rect -1850 6489 -1830 6509
rect -1810 6489 -1790 6509
rect -1770 6489 -1750 6509
rect -1730 6489 -1710 6509
rect -1690 6489 -1670 6509
rect -1650 6489 -1630 6509
rect -1610 6489 -1590 6509
rect -1570 6489 -1550 6509
rect -1530 6489 -1510 6509
rect -1490 6489 -1470 6509
rect -1450 6489 -1430 6509
rect -1410 6489 -1390 6509
rect -1370 6489 -1350 6509
rect -1330 6489 -1310 6509
rect -1290 6489 -1270 6509
rect -1250 6489 -1230 6509
rect -1210 6489 -1190 6509
rect -1170 6489 -1150 6509
rect -1130 6489 -1110 6509
rect -1090 6489 -1070 6509
rect -1050 6489 -1030 6509
rect -1010 6489 -990 6509
rect -970 6489 -950 6509
rect -930 6489 -910 6509
rect -890 6489 -870 6509
rect -850 6489 -830 6509
rect -810 6489 -790 6509
rect -770 6489 -750 6509
rect -730 6489 -710 6509
rect -690 6489 -670 6509
rect -650 6489 -630 6509
rect -610 6489 -590 6509
rect -570 6489 -550 6509
rect -530 6489 -510 6509
rect -490 6489 -470 6509
rect -450 6489 -430 6509
rect -410 6489 -390 6509
rect -370 6489 -350 6509
rect -330 6489 -310 6509
rect -290 6489 -270 6509
rect -250 6489 -230 6509
rect -210 6489 -190 6509
rect -170 6489 -150 6509
rect -130 6489 -110 6509
rect -90 6489 -70 6509
rect -50 6489 -30 6509
rect -10 6489 10 6509
rect 30 6489 50 6509
rect 70 6489 90 6509
rect 110 6489 130 6509
rect 150 6489 170 6509
rect 190 6489 210 6509
rect 230 6489 250 6509
rect 270 6489 290 6509
rect 310 6489 330 6509
rect 350 6489 370 6509
rect 390 6489 410 6509
rect 430 6489 450 6509
rect 470 6489 490 6509
rect 510 6489 525 6509
rect -2225 6450 -2175 6470
rect -2225 6430 -2210 6450
rect -2190 6430 -2175 6450
rect -2150 6470 -1995 6480
rect -1975 6479 525 6489
rect 585 6510 600 6530
rect 620 6510 635 6530
rect 585 6490 635 6510
rect -2150 6450 -2140 6470
rect -2120 6450 -2100 6470
rect -2080 6450 -2060 6470
rect -2040 6450 -2020 6470
rect -2150 6440 -1995 6450
rect 585 6470 600 6490
rect 620 6470 635 6490
rect 585 6450 635 6470
rect -2225 6410 -2175 6430
rect -2225 6390 -2210 6410
rect -2190 6390 -2175 6410
rect -1975 6427 525 6437
rect -1975 6407 -1950 6427
rect -1930 6407 -1910 6427
rect -1890 6407 -1870 6427
rect -1850 6407 -1830 6427
rect -1810 6407 -1790 6427
rect -1770 6407 -1750 6427
rect -1730 6407 -1710 6427
rect -1690 6407 -1670 6427
rect -1650 6407 -1630 6427
rect -1610 6407 -1590 6427
rect -1570 6407 -1550 6427
rect -1530 6407 -1510 6427
rect -1490 6407 -1470 6427
rect -1450 6407 -1430 6427
rect -1410 6407 -1390 6427
rect -1370 6407 -1350 6427
rect -1330 6407 -1310 6427
rect -1290 6407 -1270 6427
rect -1250 6407 -1230 6427
rect -1210 6407 -1190 6427
rect -1170 6407 -1150 6427
rect -1130 6407 -1110 6427
rect -1090 6407 -1070 6427
rect -1050 6407 -1030 6427
rect -1010 6407 -990 6427
rect -970 6407 -950 6427
rect -930 6407 -910 6427
rect -890 6407 -870 6427
rect -850 6407 -830 6427
rect -810 6407 -790 6427
rect -770 6407 -750 6427
rect -730 6407 -710 6427
rect -690 6407 -670 6427
rect -650 6407 -630 6427
rect -610 6407 -590 6427
rect -570 6407 -550 6427
rect -530 6407 -510 6427
rect -490 6407 -470 6427
rect -450 6407 -430 6427
rect -410 6407 -390 6427
rect -370 6407 -350 6427
rect -330 6407 -310 6427
rect -290 6407 -270 6427
rect -250 6407 -230 6427
rect -210 6407 -190 6427
rect -170 6407 -150 6427
rect -130 6407 -110 6427
rect -90 6407 -70 6427
rect -50 6407 -30 6427
rect -10 6407 10 6427
rect 30 6407 50 6427
rect 70 6407 90 6427
rect 110 6407 130 6427
rect 150 6407 170 6427
rect 190 6407 210 6427
rect 230 6407 250 6427
rect 270 6407 290 6427
rect 310 6407 330 6427
rect 350 6407 370 6427
rect 390 6407 410 6427
rect 430 6407 450 6427
rect 470 6407 490 6427
rect 510 6407 525 6427
rect -2225 6370 -2175 6390
rect -2225 6350 -2210 6370
rect -2190 6350 -2175 6370
rect -2150 6390 -1995 6400
rect -1975 6397 525 6407
rect 585 6430 600 6450
rect 620 6430 635 6450
rect 585 6410 635 6430
rect -2150 6370 -2140 6390
rect -2120 6370 -2100 6390
rect -2080 6370 -2060 6390
rect -2040 6370 -2020 6390
rect -2150 6360 -1995 6370
rect 585 6390 600 6410
rect 620 6390 635 6410
rect 585 6370 635 6390
rect -2225 6330 -2175 6350
rect -2225 6310 -2210 6330
rect -2190 6310 -2175 6330
rect -2225 6290 -2175 6310
rect -2225 6270 -2210 6290
rect -2190 6270 -2175 6290
rect -1975 6345 525 6355
rect -1975 6325 -1950 6345
rect -1930 6325 -1910 6345
rect -1890 6325 -1870 6345
rect -1850 6325 -1830 6345
rect -1810 6325 -1790 6345
rect -1770 6325 -1750 6345
rect -1730 6325 -1710 6345
rect -1690 6325 -1670 6345
rect -1650 6325 -1630 6345
rect -1610 6325 -1590 6345
rect -1570 6325 -1550 6345
rect -1530 6325 -1510 6345
rect -1490 6325 -1470 6345
rect -1450 6325 -1430 6345
rect -1410 6325 -1390 6345
rect -1370 6325 -1350 6345
rect -1330 6325 -1310 6345
rect -1290 6325 -1270 6345
rect -1250 6325 -1230 6345
rect -1210 6325 -1190 6345
rect -1170 6325 -1150 6345
rect -1130 6325 -1110 6345
rect -1090 6325 -1070 6345
rect -1050 6325 -1030 6345
rect -1010 6325 -990 6345
rect -970 6325 -950 6345
rect -930 6325 -910 6345
rect -890 6325 -870 6345
rect -850 6325 -830 6345
rect -810 6325 -790 6345
rect -770 6325 -750 6345
rect -730 6325 -710 6345
rect -690 6325 -670 6345
rect -650 6325 -630 6345
rect -610 6325 -590 6345
rect -570 6325 -550 6345
rect -530 6325 -510 6345
rect -490 6325 -470 6345
rect -450 6325 -430 6345
rect -410 6325 -390 6345
rect -370 6325 -350 6345
rect -330 6325 -310 6345
rect -290 6325 -270 6345
rect -250 6325 -230 6345
rect -210 6325 -190 6345
rect -170 6325 -150 6345
rect -130 6325 -110 6345
rect -90 6325 -70 6345
rect -50 6325 -30 6345
rect -10 6325 10 6345
rect 30 6325 50 6345
rect 70 6325 90 6345
rect 110 6325 130 6345
rect 150 6325 170 6345
rect 190 6325 210 6345
rect 230 6325 250 6345
rect 270 6325 290 6345
rect 310 6325 330 6345
rect 350 6325 370 6345
rect 390 6325 410 6345
rect 430 6325 450 6345
rect 470 6325 490 6345
rect 510 6325 525 6345
rect -1975 6305 525 6325
rect -1975 6285 -1950 6305
rect -1930 6285 -1910 6305
rect -1890 6285 -1870 6305
rect -1850 6285 -1830 6305
rect -1810 6285 -1790 6305
rect -1770 6285 -1750 6305
rect -1730 6285 -1710 6305
rect -1690 6285 -1670 6305
rect -1650 6285 -1630 6305
rect -1610 6285 -1590 6305
rect -1570 6285 -1550 6305
rect -1530 6285 -1510 6305
rect -1490 6285 -1470 6305
rect -1450 6285 -1430 6305
rect -1410 6285 -1390 6305
rect -1370 6285 -1350 6305
rect -1330 6285 -1310 6305
rect -1290 6285 -1270 6305
rect -1250 6285 -1230 6305
rect -1210 6285 -1190 6305
rect -1170 6285 -1150 6305
rect -1130 6285 -1110 6305
rect -1090 6285 -1070 6305
rect -1050 6285 -1030 6305
rect -1010 6285 -990 6305
rect -970 6285 -950 6305
rect -930 6285 -910 6305
rect -890 6285 -870 6305
rect -850 6285 -830 6305
rect -810 6285 -790 6305
rect -770 6285 -750 6305
rect -730 6285 -710 6305
rect -690 6285 -670 6305
rect -650 6285 -630 6305
rect -610 6285 -590 6305
rect -570 6285 -550 6305
rect -530 6285 -510 6305
rect -490 6285 -470 6305
rect -450 6285 -430 6305
rect -410 6285 -390 6305
rect -370 6285 -350 6305
rect -330 6285 -310 6305
rect -290 6285 -270 6305
rect -250 6285 -230 6305
rect -210 6285 -190 6305
rect -170 6285 -150 6305
rect -130 6285 -110 6305
rect -90 6285 -70 6305
rect -50 6285 -30 6305
rect -10 6285 10 6305
rect 30 6285 50 6305
rect 70 6285 90 6305
rect 110 6285 130 6305
rect 150 6285 170 6305
rect 190 6285 210 6305
rect 230 6285 250 6305
rect 270 6285 290 6305
rect 310 6285 330 6305
rect 350 6285 370 6305
rect 390 6285 410 6305
rect 430 6285 450 6305
rect 470 6285 490 6305
rect 510 6285 525 6305
rect -1975 6275 525 6285
rect 585 6350 600 6370
rect 620 6350 635 6370
rect 585 6330 635 6350
rect 585 6310 600 6330
rect 620 6310 635 6330
rect 585 6290 635 6310
rect -2225 6250 -2175 6270
rect -2225 6230 -2210 6250
rect -2190 6235 -2175 6250
rect 585 6270 600 6290
rect 620 6270 635 6290
rect 585 6250 635 6270
rect 585 6235 600 6250
rect -2190 6230 600 6235
rect 620 6230 635 6250
rect -2225 6220 635 6230
rect -2225 6200 -2170 6220
rect -2150 6200 -2130 6220
rect -2110 6200 -2090 6220
rect -2070 6200 -2050 6220
rect -2030 6200 -2010 6220
rect -1990 6200 -1970 6220
rect -1950 6200 -1930 6220
rect -1910 6200 -1890 6220
rect -1870 6200 -1850 6220
rect -1830 6200 -1810 6220
rect -1790 6200 -1770 6220
rect -1750 6200 -1730 6220
rect -1710 6200 -1690 6220
rect -1670 6200 -1650 6220
rect -1630 6200 -1610 6220
rect -1590 6200 -1570 6220
rect -1550 6200 -1530 6220
rect -1510 6200 -1490 6220
rect -1470 6200 -1450 6220
rect -1430 6200 -1410 6220
rect -1390 6200 -1370 6220
rect -1350 6200 -1330 6220
rect -1310 6200 -1290 6220
rect -1270 6200 -1250 6220
rect -1230 6200 -1210 6220
rect -1190 6200 -1170 6220
rect -1150 6200 -1130 6220
rect -1110 6200 -1090 6220
rect -1070 6200 -1050 6220
rect -1030 6200 -1010 6220
rect -990 6200 -970 6220
rect -950 6200 -930 6220
rect -910 6200 -890 6220
rect -870 6200 -850 6220
rect -830 6200 -810 6220
rect -790 6200 -770 6220
rect -750 6200 -730 6220
rect -710 6200 -690 6220
rect -670 6200 -650 6220
rect -630 6200 -610 6220
rect -590 6200 -570 6220
rect -550 6200 -530 6220
rect -510 6200 -490 6220
rect -470 6200 -450 6220
rect -430 6200 -410 6220
rect -390 6200 -370 6220
rect -350 6200 -330 6220
rect -310 6200 -290 6220
rect -270 6200 -250 6220
rect -230 6200 -210 6220
rect -190 6200 -170 6220
rect -150 6200 -130 6220
rect -110 6200 -90 6220
rect -70 6200 -50 6220
rect -30 6200 -10 6220
rect 10 6200 30 6220
rect 50 6200 70 6220
rect 90 6200 110 6220
rect 130 6200 150 6220
rect 170 6200 190 6220
rect 210 6200 230 6220
rect 250 6200 270 6220
rect 290 6200 310 6220
rect 330 6200 350 6220
rect 370 6200 390 6220
rect 410 6200 430 6220
rect 450 6200 470 6220
rect 490 6200 510 6220
rect 530 6200 550 6220
rect 570 6200 635 6220
rect -2225 6185 635 6200
rect -5595 6085 -3095 6095
rect -5595 6065 -5580 6085
rect -5550 6065 -5530 6085
rect -5510 6065 -5490 6085
rect -5470 6065 -5450 6085
rect -5430 6065 -5410 6085
rect -5390 6065 -5370 6085
rect -5350 6065 -5330 6085
rect -5310 6065 -5290 6085
rect -5270 6065 -5250 6085
rect -5230 6065 -5210 6085
rect -5190 6065 -5170 6085
rect -5150 6065 -5130 6085
rect -5110 6065 -5090 6085
rect -5070 6065 -5050 6085
rect -5030 6065 -5010 6085
rect -4990 6065 -4970 6085
rect -4950 6065 -4930 6085
rect -4910 6065 -4890 6085
rect -4870 6065 -4850 6085
rect -4830 6065 -4810 6085
rect -4790 6065 -4770 6085
rect -4750 6065 -4730 6085
rect -4710 6065 -4690 6085
rect -4670 6065 -4650 6085
rect -4630 6065 -4610 6085
rect -4590 6065 -4570 6085
rect -4550 6065 -4530 6085
rect -4510 6065 -4490 6085
rect -4470 6065 -4450 6085
rect -4430 6065 -4410 6085
rect -4390 6065 -4370 6085
rect -4350 6065 -4330 6085
rect -4310 6065 -4290 6085
rect -4270 6065 -4250 6085
rect -4230 6065 -4210 6085
rect -4190 6065 -4170 6085
rect -4150 6065 -4130 6085
rect -4110 6065 -4090 6085
rect -4070 6065 -4050 6085
rect -4030 6065 -4010 6085
rect -3990 6065 -3970 6085
rect -3950 6065 -3930 6085
rect -3910 6065 -3890 6085
rect -3870 6065 -3850 6085
rect -3830 6065 -3810 6085
rect -3790 6065 -3770 6085
rect -3750 6065 -3730 6085
rect -3710 6065 -3690 6085
rect -3670 6065 -3650 6085
rect -3630 6065 -3610 6085
rect -3590 6065 -3570 6085
rect -3550 6065 -3530 6085
rect -3510 6065 -3490 6085
rect -3470 6065 -3450 6085
rect -3430 6065 -3410 6085
rect -3390 6065 -3370 6085
rect -3350 6065 -3330 6085
rect -3310 6065 -3290 6085
rect -3270 6065 -3250 6085
rect -3230 6065 -3210 6085
rect -3190 6065 -3170 6085
rect -3150 6065 -3130 6085
rect -3110 6065 -3095 6085
rect -5595 6045 -3095 6065
rect -5595 6025 -5580 6045
rect -5550 6025 -5530 6045
rect -5510 6025 -5490 6045
rect -5470 6025 -5450 6045
rect -5430 6025 -5410 6045
rect -5390 6025 -5370 6045
rect -5350 6025 -5330 6045
rect -5310 6025 -5290 6045
rect -5270 6025 -5250 6045
rect -5230 6025 -5210 6045
rect -5190 6025 -5170 6045
rect -5150 6025 -5130 6045
rect -5110 6025 -5090 6045
rect -5070 6025 -5050 6045
rect -5030 6025 -5010 6045
rect -4990 6025 -4970 6045
rect -4950 6025 -4930 6045
rect -4910 6025 -4890 6045
rect -4870 6025 -4850 6045
rect -4830 6025 -4810 6045
rect -4790 6025 -4770 6045
rect -4750 6025 -4730 6045
rect -4710 6025 -4690 6045
rect -4670 6025 -4650 6045
rect -4630 6025 -4610 6045
rect -4590 6025 -4570 6045
rect -4550 6025 -4530 6045
rect -4510 6025 -4490 6045
rect -4470 6025 -4450 6045
rect -4430 6025 -4410 6045
rect -4390 6025 -4370 6045
rect -4350 6025 -4330 6045
rect -4310 6025 -4290 6045
rect -4270 6025 -4250 6045
rect -4230 6025 -4210 6045
rect -4190 6025 -4170 6045
rect -4150 6025 -4130 6045
rect -4110 6025 -4090 6045
rect -4070 6025 -4050 6045
rect -4030 6025 -4010 6045
rect -3990 6025 -3970 6045
rect -3950 6025 -3930 6045
rect -3910 6025 -3890 6045
rect -3870 6025 -3850 6045
rect -3830 6025 -3810 6045
rect -3790 6025 -3770 6045
rect -3750 6025 -3730 6045
rect -3710 6025 -3690 6045
rect -3670 6025 -3650 6045
rect -3630 6025 -3610 6045
rect -3590 6025 -3570 6045
rect -3550 6025 -3530 6045
rect -3510 6025 -3490 6045
rect -3470 6025 -3450 6045
rect -3430 6025 -3410 6045
rect -3390 6025 -3370 6045
rect -3350 6025 -3330 6045
rect -3310 6025 -3290 6045
rect -3270 6025 -3250 6045
rect -3230 6025 -3210 6045
rect -3190 6025 -3170 6045
rect -3150 6025 -3130 6045
rect -3110 6025 -3095 6045
rect -5595 6015 -3095 6025
rect -2045 6085 455 6095
rect -2045 6065 -2030 6085
rect -2010 6065 -1990 6085
rect -1970 6065 -1950 6085
rect -1930 6065 -1910 6085
rect -1890 6065 -1870 6085
rect -1850 6065 -1830 6085
rect -1810 6065 -1790 6085
rect -1770 6065 -1750 6085
rect -1730 6065 -1710 6085
rect -1690 6065 -1670 6085
rect -1650 6065 -1630 6085
rect -1610 6065 -1590 6085
rect -1570 6065 -1550 6085
rect -1530 6065 -1510 6085
rect -1490 6065 -1470 6085
rect -1450 6065 -1430 6085
rect -1410 6065 -1390 6085
rect -1370 6065 -1350 6085
rect -1330 6065 -1310 6085
rect -1290 6065 -1270 6085
rect -1250 6065 -1230 6085
rect -1210 6065 -1190 6085
rect -1170 6065 -1150 6085
rect -1130 6065 -1110 6085
rect -1090 6065 -1070 6085
rect -1050 6065 -1030 6085
rect -1010 6065 -990 6085
rect -970 6065 -950 6085
rect -930 6065 -910 6085
rect -890 6065 -870 6085
rect -850 6065 -830 6085
rect -810 6065 -790 6085
rect -770 6065 -750 6085
rect -730 6065 -710 6085
rect -690 6065 -670 6085
rect -650 6065 -630 6085
rect -610 6065 -590 6085
rect -570 6065 -550 6085
rect -530 6065 -510 6085
rect -490 6065 -470 6085
rect -450 6065 -430 6085
rect -410 6065 -390 6085
rect -370 6065 -350 6085
rect -330 6065 -310 6085
rect -290 6065 -270 6085
rect -250 6065 -230 6085
rect -210 6065 -190 6085
rect -170 6065 -150 6085
rect -130 6065 -110 6085
rect -90 6065 -70 6085
rect -50 6065 -30 6085
rect -10 6065 10 6085
rect 30 6065 50 6085
rect 70 6065 90 6085
rect 110 6065 130 6085
rect 150 6065 170 6085
rect 190 6065 210 6085
rect 230 6065 250 6085
rect 270 6065 290 6085
rect 310 6065 330 6085
rect 350 6065 370 6085
rect 390 6065 410 6085
rect 440 6065 455 6085
rect -2045 6045 455 6065
rect -2045 6025 -2030 6045
rect -2010 6025 -1990 6045
rect -1970 6025 -1950 6045
rect -1930 6025 -1910 6045
rect -1890 6025 -1870 6045
rect -1850 6025 -1830 6045
rect -1810 6025 -1790 6045
rect -1770 6025 -1750 6045
rect -1730 6025 -1710 6045
rect -1690 6025 -1670 6045
rect -1650 6025 -1630 6045
rect -1610 6025 -1590 6045
rect -1570 6025 -1550 6045
rect -1530 6025 -1510 6045
rect -1490 6025 -1470 6045
rect -1450 6025 -1430 6045
rect -1410 6025 -1390 6045
rect -1370 6025 -1350 6045
rect -1330 6025 -1310 6045
rect -1290 6025 -1270 6045
rect -1250 6025 -1230 6045
rect -1210 6025 -1190 6045
rect -1170 6025 -1150 6045
rect -1130 6025 -1110 6045
rect -1090 6025 -1070 6045
rect -1050 6025 -1030 6045
rect -1010 6025 -990 6045
rect -970 6025 -950 6045
rect -930 6025 -910 6045
rect -890 6025 -870 6045
rect -850 6025 -830 6045
rect -810 6025 -790 6045
rect -770 6025 -750 6045
rect -730 6025 -710 6045
rect -690 6025 -670 6045
rect -650 6025 -630 6045
rect -610 6025 -590 6045
rect -570 6025 -550 6045
rect -530 6025 -510 6045
rect -490 6025 -470 6045
rect -450 6025 -430 6045
rect -410 6025 -390 6045
rect -370 6025 -350 6045
rect -330 6025 -310 6045
rect -290 6025 -270 6045
rect -250 6025 -230 6045
rect -210 6025 -190 6045
rect -170 6025 -150 6045
rect -130 6025 -110 6045
rect -90 6025 -70 6045
rect -50 6025 -30 6045
rect -10 6025 10 6045
rect 30 6025 50 6045
rect 70 6025 90 6045
rect 110 6025 130 6045
rect 150 6025 170 6045
rect 190 6025 210 6045
rect 230 6025 250 6045
rect 270 6025 290 6045
rect 310 6025 330 6045
rect 350 6025 370 6045
rect 390 6025 410 6045
rect 440 6025 455 6045
rect -2045 6015 455 6025
rect -3075 6000 -2920 6010
rect -3050 5975 -3030 6000
rect -3010 5975 -2990 6000
rect -2970 5975 -2950 6000
rect -2930 5975 -2920 6000
rect -3075 5965 -2920 5975
rect -2220 6000 -2065 6010
rect -2220 5975 -2210 6000
rect -2190 5975 -2170 6000
rect -2150 5975 -2130 6000
rect -2110 5975 -2090 6000
rect -2220 5965 -2065 5975
rect -5595 5950 -3095 5960
rect -5595 5930 -5580 5950
rect -5550 5930 -5530 5950
rect -5510 5930 -5490 5950
rect -5470 5930 -5450 5950
rect -5430 5930 -5410 5950
rect -5390 5930 -5370 5950
rect -5350 5930 -5330 5950
rect -5310 5930 -5290 5950
rect -5270 5930 -5250 5950
rect -5230 5930 -5210 5950
rect -5190 5930 -5170 5950
rect -5150 5930 -5130 5950
rect -5110 5930 -5090 5950
rect -5070 5930 -5050 5950
rect -5030 5930 -5010 5950
rect -4990 5930 -4970 5950
rect -4950 5930 -4930 5950
rect -4910 5930 -4890 5950
rect -4870 5930 -4850 5950
rect -4830 5930 -4810 5950
rect -4790 5930 -4770 5950
rect -4750 5930 -4730 5950
rect -4710 5930 -4690 5950
rect -4670 5930 -4650 5950
rect -4630 5930 -4610 5950
rect -4590 5930 -4570 5950
rect -4550 5930 -4530 5950
rect -4510 5930 -4490 5950
rect -4470 5930 -4450 5950
rect -4430 5930 -4410 5950
rect -4390 5930 -4370 5950
rect -4350 5930 -4330 5950
rect -4310 5930 -4290 5950
rect -4270 5930 -4250 5950
rect -4230 5930 -4210 5950
rect -4190 5930 -4170 5950
rect -4150 5930 -4130 5950
rect -4110 5930 -4090 5950
rect -4070 5930 -4050 5950
rect -4030 5930 -4010 5950
rect -3990 5930 -3970 5950
rect -3950 5930 -3930 5950
rect -3910 5930 -3890 5950
rect -3870 5930 -3850 5950
rect -3830 5930 -3810 5950
rect -3790 5930 -3770 5950
rect -3750 5930 -3730 5950
rect -3710 5930 -3690 5950
rect -3670 5930 -3650 5950
rect -3630 5930 -3610 5950
rect -3590 5930 -3570 5950
rect -3550 5930 -3530 5950
rect -3510 5930 -3490 5950
rect -3470 5930 -3450 5950
rect -3430 5930 -3410 5950
rect -3390 5930 -3370 5950
rect -3350 5930 -3330 5950
rect -3310 5930 -3290 5950
rect -3270 5930 -3250 5950
rect -3230 5930 -3210 5950
rect -3190 5930 -3170 5950
rect -3150 5930 -3130 5950
rect -3110 5930 -3095 5950
rect -5595 5920 -3095 5930
rect -2045 5950 455 5960
rect -2045 5930 -2030 5950
rect -2010 5930 -1990 5950
rect -1970 5930 -1950 5950
rect -1930 5930 -1910 5950
rect -1890 5930 -1870 5950
rect -1850 5930 -1830 5950
rect -1810 5930 -1790 5950
rect -1770 5930 -1750 5950
rect -1730 5930 -1710 5950
rect -1690 5930 -1670 5950
rect -1650 5930 -1630 5950
rect -1610 5930 -1590 5950
rect -1570 5930 -1550 5950
rect -1530 5930 -1510 5950
rect -1490 5930 -1470 5950
rect -1450 5930 -1430 5950
rect -1410 5930 -1390 5950
rect -1370 5930 -1350 5950
rect -1330 5930 -1310 5950
rect -1290 5930 -1270 5950
rect -1250 5930 -1230 5950
rect -1210 5930 -1190 5950
rect -1170 5930 -1150 5950
rect -1130 5930 -1110 5950
rect -1090 5930 -1070 5950
rect -1050 5930 -1030 5950
rect -1010 5930 -990 5950
rect -970 5930 -950 5950
rect -930 5930 -910 5950
rect -890 5930 -870 5950
rect -850 5930 -830 5950
rect -810 5930 -790 5950
rect -770 5930 -750 5950
rect -730 5930 -710 5950
rect -690 5930 -670 5950
rect -650 5930 -630 5950
rect -610 5930 -590 5950
rect -570 5930 -550 5950
rect -530 5930 -510 5950
rect -490 5930 -470 5950
rect -450 5930 -430 5950
rect -410 5930 -390 5950
rect -370 5930 -350 5950
rect -330 5930 -310 5950
rect -290 5930 -270 5950
rect -250 5930 -230 5950
rect -210 5930 -190 5950
rect -170 5930 -150 5950
rect -130 5930 -110 5950
rect -90 5930 -70 5950
rect -50 5930 -30 5950
rect -10 5930 10 5950
rect 30 5930 50 5950
rect 70 5930 90 5950
rect 110 5930 130 5950
rect 150 5930 170 5950
rect 190 5930 210 5950
rect 230 5930 250 5950
rect 270 5930 290 5950
rect 310 5930 330 5950
rect 350 5930 370 5950
rect 390 5930 410 5950
rect 440 5930 455 5950
rect -2045 5920 455 5930
rect -3075 5905 -2920 5915
rect -3050 5880 -3030 5905
rect -3010 5880 -2990 5905
rect -2970 5880 -2950 5905
rect -2930 5880 -2920 5905
rect -3075 5870 -2920 5880
rect -2220 5905 -2065 5915
rect -2220 5880 -2210 5905
rect -2190 5880 -2170 5905
rect -2150 5880 -2130 5905
rect -2110 5880 -2090 5905
rect -2220 5870 -2065 5880
rect -5595 5855 -3095 5865
rect -5595 5835 -5580 5855
rect -5550 5835 -5530 5855
rect -5510 5835 -5490 5855
rect -5470 5835 -5450 5855
rect -5430 5835 -5410 5855
rect -5390 5835 -5370 5855
rect -5350 5835 -5330 5855
rect -5310 5835 -5290 5855
rect -5270 5835 -5250 5855
rect -5230 5835 -5210 5855
rect -5190 5835 -5170 5855
rect -5150 5835 -5130 5855
rect -5110 5835 -5090 5855
rect -5070 5835 -5050 5855
rect -5030 5835 -5010 5855
rect -4990 5835 -4970 5855
rect -4950 5835 -4930 5855
rect -4910 5835 -4890 5855
rect -4870 5835 -4850 5855
rect -4830 5835 -4810 5855
rect -4790 5835 -4770 5855
rect -4750 5835 -4730 5855
rect -4710 5835 -4690 5855
rect -4670 5835 -4650 5855
rect -4630 5835 -4610 5855
rect -4590 5835 -4570 5855
rect -4550 5835 -4530 5855
rect -4510 5835 -4490 5855
rect -4470 5835 -4450 5855
rect -4430 5835 -4410 5855
rect -4390 5835 -4370 5855
rect -4350 5835 -4330 5855
rect -4310 5835 -4290 5855
rect -4270 5835 -4250 5855
rect -4230 5835 -4210 5855
rect -4190 5835 -4170 5855
rect -4150 5835 -4130 5855
rect -4110 5835 -4090 5855
rect -4070 5835 -4050 5855
rect -4030 5835 -4010 5855
rect -3990 5835 -3970 5855
rect -3950 5835 -3930 5855
rect -3910 5835 -3890 5855
rect -3870 5835 -3850 5855
rect -3830 5835 -3810 5855
rect -3790 5835 -3770 5855
rect -3750 5835 -3730 5855
rect -3710 5835 -3690 5855
rect -3670 5835 -3650 5855
rect -3630 5835 -3610 5855
rect -3590 5835 -3570 5855
rect -3550 5835 -3530 5855
rect -3510 5835 -3490 5855
rect -3470 5835 -3450 5855
rect -3430 5835 -3410 5855
rect -3390 5835 -3370 5855
rect -3350 5835 -3330 5855
rect -3310 5835 -3290 5855
rect -3270 5835 -3250 5855
rect -3230 5835 -3210 5855
rect -3190 5835 -3170 5855
rect -3150 5835 -3130 5855
rect -3110 5835 -3095 5855
rect -5595 5825 -3095 5835
rect -2045 5855 455 5865
rect -2045 5835 -2030 5855
rect -2010 5835 -1990 5855
rect -1970 5835 -1950 5855
rect -1930 5835 -1910 5855
rect -1890 5835 -1870 5855
rect -1850 5835 -1830 5855
rect -1810 5835 -1790 5855
rect -1770 5835 -1750 5855
rect -1730 5835 -1710 5855
rect -1690 5835 -1670 5855
rect -1650 5835 -1630 5855
rect -1610 5835 -1590 5855
rect -1570 5835 -1550 5855
rect -1530 5835 -1510 5855
rect -1490 5835 -1470 5855
rect -1450 5835 -1430 5855
rect -1410 5835 -1390 5855
rect -1370 5835 -1350 5855
rect -1330 5835 -1310 5855
rect -1290 5835 -1270 5855
rect -1250 5835 -1230 5855
rect -1210 5835 -1190 5855
rect -1170 5835 -1150 5855
rect -1130 5835 -1110 5855
rect -1090 5835 -1070 5855
rect -1050 5835 -1030 5855
rect -1010 5835 -990 5855
rect -970 5835 -950 5855
rect -930 5835 -910 5855
rect -890 5835 -870 5855
rect -850 5835 -830 5855
rect -810 5835 -790 5855
rect -770 5835 -750 5855
rect -730 5835 -710 5855
rect -690 5835 -670 5855
rect -650 5835 -630 5855
rect -610 5835 -590 5855
rect -570 5835 -550 5855
rect -530 5835 -510 5855
rect -490 5835 -470 5855
rect -450 5835 -430 5855
rect -410 5835 -390 5855
rect -370 5835 -350 5855
rect -330 5835 -310 5855
rect -290 5835 -270 5855
rect -250 5835 -230 5855
rect -210 5835 -190 5855
rect -170 5835 -150 5855
rect -130 5835 -110 5855
rect -90 5835 -70 5855
rect -50 5835 -30 5855
rect -10 5835 10 5855
rect 30 5835 50 5855
rect 70 5835 90 5855
rect 110 5835 130 5855
rect 150 5835 170 5855
rect 190 5835 210 5855
rect 230 5835 250 5855
rect 270 5835 290 5855
rect 310 5835 330 5855
rect 350 5835 370 5855
rect 390 5835 410 5855
rect 440 5835 455 5855
rect -2045 5825 455 5835
rect -3075 5810 -2920 5820
rect -3050 5785 -3030 5810
rect -3010 5785 -2990 5810
rect -2970 5785 -2950 5810
rect -2930 5785 -2920 5810
rect -3075 5775 -2920 5785
rect -2220 5810 -2065 5820
rect -2220 5785 -2210 5810
rect -2190 5785 -2170 5810
rect -2150 5785 -2130 5810
rect -2110 5785 -2090 5810
rect -2220 5775 -2065 5785
rect -5595 5760 -3095 5770
rect -5595 5740 -5580 5760
rect -5550 5740 -5530 5760
rect -5510 5740 -5490 5760
rect -5470 5740 -5450 5760
rect -5430 5740 -5410 5760
rect -5390 5740 -5370 5760
rect -5350 5740 -5330 5760
rect -5310 5740 -5290 5760
rect -5270 5740 -5250 5760
rect -5230 5740 -5210 5760
rect -5190 5740 -5170 5760
rect -5150 5740 -5130 5760
rect -5110 5740 -5090 5760
rect -5070 5740 -5050 5760
rect -5030 5740 -5010 5760
rect -4990 5740 -4970 5760
rect -4950 5740 -4930 5760
rect -4910 5740 -4890 5760
rect -4870 5740 -4850 5760
rect -4830 5740 -4810 5760
rect -4790 5740 -4770 5760
rect -4750 5740 -4730 5760
rect -4710 5740 -4690 5760
rect -4670 5740 -4650 5760
rect -4630 5740 -4610 5760
rect -4590 5740 -4570 5760
rect -4550 5740 -4530 5760
rect -4510 5740 -4490 5760
rect -4470 5740 -4450 5760
rect -4430 5740 -4410 5760
rect -4390 5740 -4370 5760
rect -4350 5740 -4330 5760
rect -4310 5740 -4290 5760
rect -4270 5740 -4250 5760
rect -4230 5740 -4210 5760
rect -4190 5740 -4170 5760
rect -4150 5740 -4130 5760
rect -4110 5740 -4090 5760
rect -4070 5740 -4050 5760
rect -4030 5740 -4010 5760
rect -3990 5740 -3970 5760
rect -3950 5740 -3930 5760
rect -3910 5740 -3890 5760
rect -3870 5740 -3850 5760
rect -3830 5740 -3810 5760
rect -3790 5740 -3770 5760
rect -3750 5740 -3730 5760
rect -3710 5740 -3690 5760
rect -3670 5740 -3650 5760
rect -3630 5740 -3610 5760
rect -3590 5740 -3570 5760
rect -3550 5740 -3530 5760
rect -3510 5740 -3490 5760
rect -3470 5740 -3450 5760
rect -3430 5740 -3410 5760
rect -3390 5740 -3370 5760
rect -3350 5740 -3330 5760
rect -3310 5740 -3290 5760
rect -3270 5740 -3250 5760
rect -3230 5740 -3210 5760
rect -3190 5740 -3170 5760
rect -3150 5740 -3130 5760
rect -3110 5740 -3095 5760
rect -5595 5730 -3095 5740
rect -2045 5760 455 5770
rect -2045 5740 -2030 5760
rect -2010 5740 -1990 5760
rect -1970 5740 -1950 5760
rect -1930 5740 -1910 5760
rect -1890 5740 -1870 5760
rect -1850 5740 -1830 5760
rect -1810 5740 -1790 5760
rect -1770 5740 -1750 5760
rect -1730 5740 -1710 5760
rect -1690 5740 -1670 5760
rect -1650 5740 -1630 5760
rect -1610 5740 -1590 5760
rect -1570 5740 -1550 5760
rect -1530 5740 -1510 5760
rect -1490 5740 -1470 5760
rect -1450 5740 -1430 5760
rect -1410 5740 -1390 5760
rect -1370 5740 -1350 5760
rect -1330 5740 -1310 5760
rect -1290 5740 -1270 5760
rect -1250 5740 -1230 5760
rect -1210 5740 -1190 5760
rect -1170 5740 -1150 5760
rect -1130 5740 -1110 5760
rect -1090 5740 -1070 5760
rect -1050 5740 -1030 5760
rect -1010 5740 -990 5760
rect -970 5740 -950 5760
rect -930 5740 -910 5760
rect -890 5740 -870 5760
rect -850 5740 -830 5760
rect -810 5740 -790 5760
rect -770 5740 -750 5760
rect -730 5740 -710 5760
rect -690 5740 -670 5760
rect -650 5740 -630 5760
rect -610 5740 -590 5760
rect -570 5740 -550 5760
rect -530 5740 -510 5760
rect -490 5740 -470 5760
rect -450 5740 -430 5760
rect -410 5740 -390 5760
rect -370 5740 -350 5760
rect -330 5740 -310 5760
rect -290 5740 -270 5760
rect -250 5740 -230 5760
rect -210 5740 -190 5760
rect -170 5740 -150 5760
rect -130 5740 -110 5760
rect -90 5740 -70 5760
rect -50 5740 -30 5760
rect -10 5740 10 5760
rect 30 5740 50 5760
rect 70 5740 90 5760
rect 110 5740 130 5760
rect 150 5740 170 5760
rect 190 5740 210 5760
rect 230 5740 250 5760
rect 270 5740 290 5760
rect 310 5740 330 5760
rect 350 5740 370 5760
rect 390 5740 410 5760
rect 440 5740 455 5760
rect -2045 5730 455 5740
rect -3075 5715 -2920 5725
rect -3050 5690 -3030 5715
rect -3010 5690 -2990 5715
rect -2970 5690 -2950 5715
rect -2930 5690 -2920 5715
rect -3075 5680 -2920 5690
rect -2220 5715 -2065 5725
rect -2220 5690 -2210 5715
rect -2190 5690 -2170 5715
rect -2150 5690 -2130 5715
rect -2110 5690 -2090 5715
rect -2220 5680 -2065 5690
rect -5595 5665 -3095 5675
rect -5595 5645 -5580 5665
rect -5550 5645 -5530 5665
rect -5510 5645 -5490 5665
rect -5470 5645 -5450 5665
rect -5430 5645 -5410 5665
rect -5390 5645 -5370 5665
rect -5350 5645 -5330 5665
rect -5310 5645 -5290 5665
rect -5270 5645 -5250 5665
rect -5230 5645 -5210 5665
rect -5190 5645 -5170 5665
rect -5150 5645 -5130 5665
rect -5110 5645 -5090 5665
rect -5070 5645 -5050 5665
rect -5030 5645 -5010 5665
rect -4990 5645 -4970 5665
rect -4950 5645 -4930 5665
rect -4910 5645 -4890 5665
rect -4870 5645 -4850 5665
rect -4830 5645 -4810 5665
rect -4790 5645 -4770 5665
rect -4750 5645 -4730 5665
rect -4710 5645 -4690 5665
rect -4670 5645 -4650 5665
rect -4630 5645 -4610 5665
rect -4590 5645 -4570 5665
rect -4550 5645 -4530 5665
rect -4510 5645 -4490 5665
rect -4470 5645 -4450 5665
rect -4430 5645 -4410 5665
rect -4390 5645 -4370 5665
rect -4350 5645 -4330 5665
rect -4310 5645 -4290 5665
rect -4270 5645 -4250 5665
rect -4230 5645 -4210 5665
rect -4190 5645 -4170 5665
rect -4150 5645 -4130 5665
rect -4110 5645 -4090 5665
rect -4070 5645 -4050 5665
rect -4030 5645 -4010 5665
rect -3990 5645 -3970 5665
rect -3950 5645 -3930 5665
rect -3910 5645 -3890 5665
rect -3870 5645 -3850 5665
rect -3830 5645 -3810 5665
rect -3790 5645 -3770 5665
rect -3750 5645 -3730 5665
rect -3710 5645 -3690 5665
rect -3670 5645 -3650 5665
rect -3630 5645 -3610 5665
rect -3590 5645 -3570 5665
rect -3550 5645 -3530 5665
rect -3510 5645 -3490 5665
rect -3470 5645 -3450 5665
rect -3430 5645 -3410 5665
rect -3390 5645 -3370 5665
rect -3350 5645 -3330 5665
rect -3310 5645 -3290 5665
rect -3270 5645 -3250 5665
rect -3230 5645 -3210 5665
rect -3190 5645 -3170 5665
rect -3150 5645 -3130 5665
rect -3110 5645 -3095 5665
rect -5595 5635 -3095 5645
rect -2045 5665 455 5675
rect -2045 5645 -2030 5665
rect -2010 5645 -1990 5665
rect -1970 5645 -1950 5665
rect -1930 5645 -1910 5665
rect -1890 5645 -1870 5665
rect -1850 5645 -1830 5665
rect -1810 5645 -1790 5665
rect -1770 5645 -1750 5665
rect -1730 5645 -1710 5665
rect -1690 5645 -1670 5665
rect -1650 5645 -1630 5665
rect -1610 5645 -1590 5665
rect -1570 5645 -1550 5665
rect -1530 5645 -1510 5665
rect -1490 5645 -1470 5665
rect -1450 5645 -1430 5665
rect -1410 5645 -1390 5665
rect -1370 5645 -1350 5665
rect -1330 5645 -1310 5665
rect -1290 5645 -1270 5665
rect -1250 5645 -1230 5665
rect -1210 5645 -1190 5665
rect -1170 5645 -1150 5665
rect -1130 5645 -1110 5665
rect -1090 5645 -1070 5665
rect -1050 5645 -1030 5665
rect -1010 5645 -990 5665
rect -970 5645 -950 5665
rect -930 5645 -910 5665
rect -890 5645 -870 5665
rect -850 5645 -830 5665
rect -810 5645 -790 5665
rect -770 5645 -750 5665
rect -730 5645 -710 5665
rect -690 5645 -670 5665
rect -650 5645 -630 5665
rect -610 5645 -590 5665
rect -570 5645 -550 5665
rect -530 5645 -510 5665
rect -490 5645 -470 5665
rect -450 5645 -430 5665
rect -410 5645 -390 5665
rect -370 5645 -350 5665
rect -330 5645 -310 5665
rect -290 5645 -270 5665
rect -250 5645 -230 5665
rect -210 5645 -190 5665
rect -170 5645 -150 5665
rect -130 5645 -110 5665
rect -90 5645 -70 5665
rect -50 5645 -30 5665
rect -10 5645 10 5665
rect 30 5645 50 5665
rect 70 5645 90 5665
rect 110 5645 130 5665
rect 150 5645 170 5665
rect 190 5645 210 5665
rect 230 5645 250 5665
rect 270 5645 290 5665
rect 310 5645 330 5665
rect 350 5645 370 5665
rect 390 5645 410 5665
rect 440 5645 455 5665
rect -2045 5635 455 5645
rect -3075 5620 -2920 5630
rect -3050 5595 -3030 5620
rect -3010 5595 -2990 5620
rect -2970 5595 -2950 5620
rect -2930 5595 -2920 5620
rect -3075 5585 -2920 5595
rect -2220 5620 -2065 5630
rect -2220 5595 -2210 5620
rect -2190 5595 -2170 5620
rect -2150 5595 -2130 5620
rect -2110 5595 -2090 5620
rect -2220 5585 -2065 5595
rect -5595 5570 -3095 5580
rect -5595 5550 -5580 5570
rect -5550 5550 -5530 5570
rect -5510 5550 -5490 5570
rect -5470 5550 -5450 5570
rect -5430 5550 -5410 5570
rect -5390 5550 -5370 5570
rect -5350 5550 -5330 5570
rect -5310 5550 -5290 5570
rect -5270 5550 -5250 5570
rect -5230 5550 -5210 5570
rect -5190 5550 -5170 5570
rect -5150 5550 -5130 5570
rect -5110 5550 -5090 5570
rect -5070 5550 -5050 5570
rect -5030 5550 -5010 5570
rect -4990 5550 -4970 5570
rect -4950 5550 -4930 5570
rect -4910 5550 -4890 5570
rect -4870 5550 -4850 5570
rect -4830 5550 -4810 5570
rect -4790 5550 -4770 5570
rect -4750 5550 -4730 5570
rect -4710 5550 -4690 5570
rect -4670 5550 -4650 5570
rect -4630 5550 -4610 5570
rect -4590 5550 -4570 5570
rect -4550 5550 -4530 5570
rect -4510 5550 -4490 5570
rect -4470 5550 -4450 5570
rect -4430 5550 -4410 5570
rect -4390 5550 -4370 5570
rect -4350 5550 -4330 5570
rect -4310 5550 -4290 5570
rect -4270 5550 -4250 5570
rect -4230 5550 -4210 5570
rect -4190 5550 -4170 5570
rect -4150 5550 -4130 5570
rect -4110 5550 -4090 5570
rect -4070 5550 -4050 5570
rect -4030 5550 -4010 5570
rect -3990 5550 -3970 5570
rect -3950 5550 -3930 5570
rect -3910 5550 -3890 5570
rect -3870 5550 -3850 5570
rect -3830 5550 -3810 5570
rect -3790 5550 -3770 5570
rect -3750 5550 -3730 5570
rect -3710 5550 -3690 5570
rect -3670 5550 -3650 5570
rect -3630 5550 -3610 5570
rect -3590 5550 -3570 5570
rect -3550 5550 -3530 5570
rect -3510 5550 -3490 5570
rect -3470 5550 -3450 5570
rect -3430 5550 -3410 5570
rect -3390 5550 -3370 5570
rect -3350 5550 -3330 5570
rect -3310 5550 -3290 5570
rect -3270 5550 -3250 5570
rect -3230 5550 -3210 5570
rect -3190 5550 -3170 5570
rect -3150 5550 -3130 5570
rect -3110 5550 -3095 5570
rect -5595 5540 -3095 5550
rect -2045 5570 455 5580
rect -2045 5550 -2030 5570
rect -2010 5550 -1990 5570
rect -1970 5550 -1950 5570
rect -1930 5550 -1910 5570
rect -1890 5550 -1870 5570
rect -1850 5550 -1830 5570
rect -1810 5550 -1790 5570
rect -1770 5550 -1750 5570
rect -1730 5550 -1710 5570
rect -1690 5550 -1670 5570
rect -1650 5550 -1630 5570
rect -1610 5550 -1590 5570
rect -1570 5550 -1550 5570
rect -1530 5550 -1510 5570
rect -1490 5550 -1470 5570
rect -1450 5550 -1430 5570
rect -1410 5550 -1390 5570
rect -1370 5550 -1350 5570
rect -1330 5550 -1310 5570
rect -1290 5550 -1270 5570
rect -1250 5550 -1230 5570
rect -1210 5550 -1190 5570
rect -1170 5550 -1150 5570
rect -1130 5550 -1110 5570
rect -1090 5550 -1070 5570
rect -1050 5550 -1030 5570
rect -1010 5550 -990 5570
rect -970 5550 -950 5570
rect -930 5550 -910 5570
rect -890 5550 -870 5570
rect -850 5550 -830 5570
rect -810 5550 -790 5570
rect -770 5550 -750 5570
rect -730 5550 -710 5570
rect -690 5550 -670 5570
rect -650 5550 -630 5570
rect -610 5550 -590 5570
rect -570 5550 -550 5570
rect -530 5550 -510 5570
rect -490 5550 -470 5570
rect -450 5550 -430 5570
rect -410 5550 -390 5570
rect -370 5550 -350 5570
rect -330 5550 -310 5570
rect -290 5550 -270 5570
rect -250 5550 -230 5570
rect -210 5550 -190 5570
rect -170 5550 -150 5570
rect -130 5550 -110 5570
rect -90 5550 -70 5570
rect -50 5550 -30 5570
rect -10 5550 10 5570
rect 30 5550 50 5570
rect 70 5550 90 5570
rect 110 5550 130 5570
rect 150 5550 170 5570
rect 190 5550 210 5570
rect 230 5550 250 5570
rect 270 5550 290 5570
rect 310 5550 330 5570
rect 350 5550 370 5570
rect 390 5550 410 5570
rect 440 5550 455 5570
rect -2045 5540 455 5550
rect -3075 5525 -2920 5535
rect -3050 5500 -3030 5525
rect -3010 5500 -2990 5525
rect -2970 5500 -2950 5525
rect -2930 5500 -2920 5525
rect -3075 5490 -2920 5500
rect -2220 5525 -2065 5535
rect -2220 5500 -2210 5525
rect -2190 5500 -2170 5525
rect -2150 5500 -2130 5525
rect -2110 5500 -2090 5525
rect -2220 5490 -2065 5500
rect -5595 5475 -3095 5485
rect -5595 5455 -5580 5475
rect -5550 5455 -5530 5475
rect -5510 5455 -5490 5475
rect -5470 5455 -5450 5475
rect -5430 5455 -5410 5475
rect -5390 5455 -5370 5475
rect -5350 5455 -5330 5475
rect -5310 5455 -5290 5475
rect -5270 5455 -5250 5475
rect -5230 5455 -5210 5475
rect -5190 5455 -5170 5475
rect -5150 5455 -5130 5475
rect -5110 5455 -5090 5475
rect -5070 5455 -5050 5475
rect -5030 5455 -5010 5475
rect -4990 5455 -4970 5475
rect -4950 5455 -4930 5475
rect -4910 5455 -4890 5475
rect -4870 5455 -4850 5475
rect -4830 5455 -4810 5475
rect -4790 5455 -4770 5475
rect -4750 5455 -4730 5475
rect -4710 5455 -4690 5475
rect -4670 5455 -4650 5475
rect -4630 5455 -4610 5475
rect -4590 5455 -4570 5475
rect -4550 5455 -4530 5475
rect -4510 5455 -4490 5475
rect -4470 5455 -4450 5475
rect -4430 5455 -4410 5475
rect -4390 5455 -4370 5475
rect -4350 5455 -4330 5475
rect -4310 5455 -4290 5475
rect -4270 5455 -4250 5475
rect -4230 5455 -4210 5475
rect -4190 5455 -4170 5475
rect -4150 5455 -4130 5475
rect -4110 5455 -4090 5475
rect -4070 5455 -4050 5475
rect -4030 5455 -4010 5475
rect -3990 5455 -3970 5475
rect -3950 5455 -3930 5475
rect -3910 5455 -3890 5475
rect -3870 5455 -3850 5475
rect -3830 5455 -3810 5475
rect -3790 5455 -3770 5475
rect -3750 5455 -3730 5475
rect -3710 5455 -3690 5475
rect -3670 5455 -3650 5475
rect -3630 5455 -3610 5475
rect -3590 5455 -3570 5475
rect -3550 5455 -3530 5475
rect -3510 5455 -3490 5475
rect -3470 5455 -3450 5475
rect -3430 5455 -3410 5475
rect -3390 5455 -3370 5475
rect -3350 5455 -3330 5475
rect -3310 5455 -3290 5475
rect -3270 5455 -3250 5475
rect -3230 5455 -3210 5475
rect -3190 5455 -3170 5475
rect -3150 5455 -3130 5475
rect -3110 5455 -3095 5475
rect -5595 5445 -3095 5455
rect -2045 5475 455 5485
rect -2045 5455 -2030 5475
rect -2010 5455 -1990 5475
rect -1970 5455 -1950 5475
rect -1930 5455 -1910 5475
rect -1890 5455 -1870 5475
rect -1850 5455 -1830 5475
rect -1810 5455 -1790 5475
rect -1770 5455 -1750 5475
rect -1730 5455 -1710 5475
rect -1690 5455 -1670 5475
rect -1650 5455 -1630 5475
rect -1610 5455 -1590 5475
rect -1570 5455 -1550 5475
rect -1530 5455 -1510 5475
rect -1490 5455 -1470 5475
rect -1450 5455 -1430 5475
rect -1410 5455 -1390 5475
rect -1370 5455 -1350 5475
rect -1330 5455 -1310 5475
rect -1290 5455 -1270 5475
rect -1250 5455 -1230 5475
rect -1210 5455 -1190 5475
rect -1170 5455 -1150 5475
rect -1130 5455 -1110 5475
rect -1090 5455 -1070 5475
rect -1050 5455 -1030 5475
rect -1010 5455 -990 5475
rect -970 5455 -950 5475
rect -930 5455 -910 5475
rect -890 5455 -870 5475
rect -850 5455 -830 5475
rect -810 5455 -790 5475
rect -770 5455 -750 5475
rect -730 5455 -710 5475
rect -690 5455 -670 5475
rect -650 5455 -630 5475
rect -610 5455 -590 5475
rect -570 5455 -550 5475
rect -530 5455 -510 5475
rect -490 5455 -470 5475
rect -450 5455 -430 5475
rect -410 5455 -390 5475
rect -370 5455 -350 5475
rect -330 5455 -310 5475
rect -290 5455 -270 5475
rect -250 5455 -230 5475
rect -210 5455 -190 5475
rect -170 5455 -150 5475
rect -130 5455 -110 5475
rect -90 5455 -70 5475
rect -50 5455 -30 5475
rect -10 5455 10 5475
rect 30 5455 50 5475
rect 70 5455 90 5475
rect 110 5455 130 5475
rect 150 5455 170 5475
rect 190 5455 210 5475
rect 230 5455 250 5475
rect 270 5455 290 5475
rect 310 5455 330 5475
rect 350 5455 370 5475
rect 390 5455 410 5475
rect 440 5455 455 5475
rect -2045 5445 455 5455
rect -3075 5430 -2920 5440
rect -3050 5405 -3030 5430
rect -3010 5405 -2990 5430
rect -2970 5405 -2950 5430
rect -2930 5405 -2920 5430
rect -3075 5395 -2920 5405
rect -2220 5430 -2065 5440
rect -2220 5405 -2210 5430
rect -2190 5405 -2170 5430
rect -2150 5405 -2130 5430
rect -2110 5405 -2090 5430
rect -2220 5395 -2065 5405
rect -5595 5380 -3095 5390
rect -5595 5360 -5580 5380
rect -5550 5360 -5530 5380
rect -5510 5360 -5490 5380
rect -5470 5360 -5450 5380
rect -5430 5360 -5410 5380
rect -5390 5360 -5370 5380
rect -5350 5360 -5330 5380
rect -5310 5360 -5290 5380
rect -5270 5360 -5250 5380
rect -5230 5360 -5210 5380
rect -5190 5360 -5170 5380
rect -5150 5360 -5130 5380
rect -5110 5360 -5090 5380
rect -5070 5360 -5050 5380
rect -5030 5360 -5010 5380
rect -4990 5360 -4970 5380
rect -4950 5360 -4930 5380
rect -4910 5360 -4890 5380
rect -4870 5360 -4850 5380
rect -4830 5360 -4810 5380
rect -4790 5360 -4770 5380
rect -4750 5360 -4730 5380
rect -4710 5360 -4690 5380
rect -4670 5360 -4650 5380
rect -4630 5360 -4610 5380
rect -4590 5360 -4570 5380
rect -4550 5360 -4530 5380
rect -4510 5360 -4490 5380
rect -4470 5360 -4450 5380
rect -4430 5360 -4410 5380
rect -4390 5360 -4370 5380
rect -4350 5360 -4330 5380
rect -4310 5360 -4290 5380
rect -4270 5360 -4250 5380
rect -4230 5360 -4210 5380
rect -4190 5360 -4170 5380
rect -4150 5360 -4130 5380
rect -4110 5360 -4090 5380
rect -4070 5360 -4050 5380
rect -4030 5360 -4010 5380
rect -3990 5360 -3970 5380
rect -3950 5360 -3930 5380
rect -3910 5360 -3890 5380
rect -3870 5360 -3850 5380
rect -3830 5360 -3810 5380
rect -3790 5360 -3770 5380
rect -3750 5360 -3730 5380
rect -3710 5360 -3690 5380
rect -3670 5360 -3650 5380
rect -3630 5360 -3610 5380
rect -3590 5360 -3570 5380
rect -3550 5360 -3530 5380
rect -3510 5360 -3490 5380
rect -3470 5360 -3450 5380
rect -3430 5360 -3410 5380
rect -3390 5360 -3370 5380
rect -3350 5360 -3330 5380
rect -3310 5360 -3290 5380
rect -3270 5360 -3250 5380
rect -3230 5360 -3210 5380
rect -3190 5360 -3170 5380
rect -3150 5360 -3130 5380
rect -3110 5360 -3095 5380
rect -5595 5350 -3095 5360
rect -2045 5380 455 5390
rect -2045 5360 -2030 5380
rect -2010 5360 -1990 5380
rect -1970 5360 -1950 5380
rect -1930 5360 -1910 5380
rect -1890 5360 -1870 5380
rect -1850 5360 -1830 5380
rect -1810 5360 -1790 5380
rect -1770 5360 -1750 5380
rect -1730 5360 -1710 5380
rect -1690 5360 -1670 5380
rect -1650 5360 -1630 5380
rect -1610 5360 -1590 5380
rect -1570 5360 -1550 5380
rect -1530 5360 -1510 5380
rect -1490 5360 -1470 5380
rect -1450 5360 -1430 5380
rect -1410 5360 -1390 5380
rect -1370 5360 -1350 5380
rect -1330 5360 -1310 5380
rect -1290 5360 -1270 5380
rect -1250 5360 -1230 5380
rect -1210 5360 -1190 5380
rect -1170 5360 -1150 5380
rect -1130 5360 -1110 5380
rect -1090 5360 -1070 5380
rect -1050 5360 -1030 5380
rect -1010 5360 -990 5380
rect -970 5360 -950 5380
rect -930 5360 -910 5380
rect -890 5360 -870 5380
rect -850 5360 -830 5380
rect -810 5360 -790 5380
rect -770 5360 -750 5380
rect -730 5360 -710 5380
rect -690 5360 -670 5380
rect -650 5360 -630 5380
rect -610 5360 -590 5380
rect -570 5360 -550 5380
rect -530 5360 -510 5380
rect -490 5360 -470 5380
rect -450 5360 -430 5380
rect -410 5360 -390 5380
rect -370 5360 -350 5380
rect -330 5360 -310 5380
rect -290 5360 -270 5380
rect -250 5360 -230 5380
rect -210 5360 -190 5380
rect -170 5360 -150 5380
rect -130 5360 -110 5380
rect -90 5360 -70 5380
rect -50 5360 -30 5380
rect -10 5360 10 5380
rect 30 5360 50 5380
rect 70 5360 90 5380
rect 110 5360 130 5380
rect 150 5360 170 5380
rect 190 5360 210 5380
rect 230 5360 250 5380
rect 270 5360 290 5380
rect 310 5360 330 5380
rect 350 5360 370 5380
rect 390 5360 410 5380
rect 440 5360 455 5380
rect -2045 5350 455 5360
rect -3075 5335 -2920 5345
rect -3050 5310 -3030 5335
rect -3010 5310 -2990 5335
rect -2970 5310 -2950 5335
rect -2930 5310 -2920 5335
rect -3075 5300 -2920 5310
rect -2220 5335 -2065 5345
rect -2220 5310 -2210 5335
rect -2190 5310 -2170 5335
rect -2150 5310 -2130 5335
rect -2110 5310 -2090 5335
rect -2220 5300 -2065 5310
rect -5595 5285 -3095 5295
rect -5595 5265 -5580 5285
rect -5550 5265 -5530 5285
rect -5510 5265 -5490 5285
rect -5470 5265 -5450 5285
rect -5430 5265 -5410 5285
rect -5390 5265 -5370 5285
rect -5350 5265 -5330 5285
rect -5310 5265 -5290 5285
rect -5270 5265 -5250 5285
rect -5230 5265 -5210 5285
rect -5190 5265 -5170 5285
rect -5150 5265 -5130 5285
rect -5110 5265 -5090 5285
rect -5070 5265 -5050 5285
rect -5030 5265 -5010 5285
rect -4990 5265 -4970 5285
rect -4950 5265 -4930 5285
rect -4910 5265 -4890 5285
rect -4870 5265 -4850 5285
rect -4830 5265 -4810 5285
rect -4790 5265 -4770 5285
rect -4750 5265 -4730 5285
rect -4710 5265 -4690 5285
rect -4670 5265 -4650 5285
rect -4630 5265 -4610 5285
rect -4590 5265 -4570 5285
rect -4550 5265 -4530 5285
rect -4510 5265 -4490 5285
rect -4470 5265 -4450 5285
rect -4430 5265 -4410 5285
rect -4390 5265 -4370 5285
rect -4350 5265 -4330 5285
rect -4310 5265 -4290 5285
rect -4270 5265 -4250 5285
rect -4230 5265 -4210 5285
rect -4190 5265 -4170 5285
rect -4150 5265 -4130 5285
rect -4110 5265 -4090 5285
rect -4070 5265 -4050 5285
rect -4030 5265 -4010 5285
rect -3990 5265 -3970 5285
rect -3950 5265 -3930 5285
rect -3910 5265 -3890 5285
rect -3870 5265 -3850 5285
rect -3830 5265 -3810 5285
rect -3790 5265 -3770 5285
rect -3750 5265 -3730 5285
rect -3710 5265 -3690 5285
rect -3670 5265 -3650 5285
rect -3630 5265 -3610 5285
rect -3590 5265 -3570 5285
rect -3550 5265 -3530 5285
rect -3510 5265 -3490 5285
rect -3470 5265 -3450 5285
rect -3430 5265 -3410 5285
rect -3390 5265 -3370 5285
rect -3350 5265 -3330 5285
rect -3310 5265 -3290 5285
rect -3270 5265 -3250 5285
rect -3230 5265 -3210 5285
rect -3190 5265 -3170 5285
rect -3150 5265 -3130 5285
rect -3110 5265 -3095 5285
rect -5595 5255 -3095 5265
rect -2045 5285 455 5295
rect -2045 5265 -2030 5285
rect -2010 5265 -1990 5285
rect -1970 5265 -1950 5285
rect -1930 5265 -1910 5285
rect -1890 5265 -1870 5285
rect -1850 5265 -1830 5285
rect -1810 5265 -1790 5285
rect -1770 5265 -1750 5285
rect -1730 5265 -1710 5285
rect -1690 5265 -1670 5285
rect -1650 5265 -1630 5285
rect -1610 5265 -1590 5285
rect -1570 5265 -1550 5285
rect -1530 5265 -1510 5285
rect -1490 5265 -1470 5285
rect -1450 5265 -1430 5285
rect -1410 5265 -1390 5285
rect -1370 5265 -1350 5285
rect -1330 5265 -1310 5285
rect -1290 5265 -1270 5285
rect -1250 5265 -1230 5285
rect -1210 5265 -1190 5285
rect -1170 5265 -1150 5285
rect -1130 5265 -1110 5285
rect -1090 5265 -1070 5285
rect -1050 5265 -1030 5285
rect -1010 5265 -990 5285
rect -970 5265 -950 5285
rect -930 5265 -910 5285
rect -890 5265 -870 5285
rect -850 5265 -830 5285
rect -810 5265 -790 5285
rect -770 5265 -750 5285
rect -730 5265 -710 5285
rect -690 5265 -670 5285
rect -650 5265 -630 5285
rect -610 5265 -590 5285
rect -570 5265 -550 5285
rect -530 5265 -510 5285
rect -490 5265 -470 5285
rect -450 5265 -430 5285
rect -410 5265 -390 5285
rect -370 5265 -350 5285
rect -330 5265 -310 5285
rect -290 5265 -270 5285
rect -250 5265 -230 5285
rect -210 5265 -190 5285
rect -170 5265 -150 5285
rect -130 5265 -110 5285
rect -90 5265 -70 5285
rect -50 5265 -30 5285
rect -10 5265 10 5285
rect 30 5265 50 5285
rect 70 5265 90 5285
rect 110 5265 130 5285
rect 150 5265 170 5285
rect 190 5265 210 5285
rect 230 5265 250 5285
rect 270 5265 290 5285
rect 310 5265 330 5285
rect 350 5265 370 5285
rect 390 5265 410 5285
rect 440 5265 455 5285
rect -2045 5255 455 5265
rect -3075 5240 -2920 5250
rect -3050 5215 -3030 5240
rect -3010 5215 -2990 5240
rect -2970 5215 -2950 5240
rect -2930 5215 -2920 5240
rect -3075 5205 -2920 5215
rect -2220 5240 -2065 5250
rect -2220 5215 -2210 5240
rect -2190 5215 -2170 5240
rect -2150 5215 -2130 5240
rect -2110 5215 -2090 5240
rect -2220 5205 -2065 5215
rect -5595 5190 -3095 5200
rect -5595 5170 -5580 5190
rect -5550 5170 -5530 5190
rect -5510 5170 -5490 5190
rect -5470 5170 -5450 5190
rect -5430 5170 -5410 5190
rect -5390 5170 -5370 5190
rect -5350 5170 -5330 5190
rect -5310 5170 -5290 5190
rect -5270 5170 -5250 5190
rect -5230 5170 -5210 5190
rect -5190 5170 -5170 5190
rect -5150 5170 -5130 5190
rect -5110 5170 -5090 5190
rect -5070 5170 -5050 5190
rect -5030 5170 -5010 5190
rect -4990 5170 -4970 5190
rect -4950 5170 -4930 5190
rect -4910 5170 -4890 5190
rect -4870 5170 -4850 5190
rect -4830 5170 -4810 5190
rect -4790 5170 -4770 5190
rect -4750 5170 -4730 5190
rect -4710 5170 -4690 5190
rect -4670 5170 -4650 5190
rect -4630 5170 -4610 5190
rect -4590 5170 -4570 5190
rect -4550 5170 -4530 5190
rect -4510 5170 -4490 5190
rect -4470 5170 -4450 5190
rect -4430 5170 -4410 5190
rect -4390 5170 -4370 5190
rect -4350 5170 -4330 5190
rect -4310 5170 -4290 5190
rect -4270 5170 -4250 5190
rect -4230 5170 -4210 5190
rect -4190 5170 -4170 5190
rect -4150 5170 -4130 5190
rect -4110 5170 -4090 5190
rect -4070 5170 -4050 5190
rect -4030 5170 -4010 5190
rect -3990 5170 -3970 5190
rect -3950 5170 -3930 5190
rect -3910 5170 -3890 5190
rect -3870 5170 -3850 5190
rect -3830 5170 -3810 5190
rect -3790 5170 -3770 5190
rect -3750 5170 -3730 5190
rect -3710 5170 -3690 5190
rect -3670 5170 -3650 5190
rect -3630 5170 -3610 5190
rect -3590 5170 -3570 5190
rect -3550 5170 -3530 5190
rect -3510 5170 -3490 5190
rect -3470 5170 -3450 5190
rect -3430 5170 -3410 5190
rect -3390 5170 -3370 5190
rect -3350 5170 -3330 5190
rect -3310 5170 -3290 5190
rect -3270 5170 -3250 5190
rect -3230 5170 -3210 5190
rect -3190 5170 -3170 5190
rect -3150 5170 -3130 5190
rect -3110 5170 -3095 5190
rect -5595 5160 -3095 5170
rect -2045 5190 455 5200
rect -2045 5170 -2030 5190
rect -2010 5170 -1990 5190
rect -1970 5170 -1950 5190
rect -1930 5170 -1910 5190
rect -1890 5170 -1870 5190
rect -1850 5170 -1830 5190
rect -1810 5170 -1790 5190
rect -1770 5170 -1750 5190
rect -1730 5170 -1710 5190
rect -1690 5170 -1670 5190
rect -1650 5170 -1630 5190
rect -1610 5170 -1590 5190
rect -1570 5170 -1550 5190
rect -1530 5170 -1510 5190
rect -1490 5170 -1470 5190
rect -1450 5170 -1430 5190
rect -1410 5170 -1390 5190
rect -1370 5170 -1350 5190
rect -1330 5170 -1310 5190
rect -1290 5170 -1270 5190
rect -1250 5170 -1230 5190
rect -1210 5170 -1190 5190
rect -1170 5170 -1150 5190
rect -1130 5170 -1110 5190
rect -1090 5170 -1070 5190
rect -1050 5170 -1030 5190
rect -1010 5170 -990 5190
rect -970 5170 -950 5190
rect -930 5170 -910 5190
rect -890 5170 -870 5190
rect -850 5170 -830 5190
rect -810 5170 -790 5190
rect -770 5170 -750 5190
rect -730 5170 -710 5190
rect -690 5170 -670 5190
rect -650 5170 -630 5190
rect -610 5170 -590 5190
rect -570 5170 -550 5190
rect -530 5170 -510 5190
rect -490 5170 -470 5190
rect -450 5170 -430 5190
rect -410 5170 -390 5190
rect -370 5170 -350 5190
rect -330 5170 -310 5190
rect -290 5170 -270 5190
rect -250 5170 -230 5190
rect -210 5170 -190 5190
rect -170 5170 -150 5190
rect -130 5170 -110 5190
rect -90 5170 -70 5190
rect -50 5170 -30 5190
rect -10 5170 10 5190
rect 30 5170 50 5190
rect 70 5170 90 5190
rect 110 5170 130 5190
rect 150 5170 170 5190
rect 190 5170 210 5190
rect 230 5170 250 5190
rect 270 5170 290 5190
rect 310 5170 330 5190
rect 350 5170 370 5190
rect 390 5170 410 5190
rect 440 5170 455 5190
rect -2045 5160 455 5170
rect -3075 5145 -2920 5155
rect -3050 5120 -3030 5145
rect -3010 5120 -2990 5145
rect -2970 5120 -2950 5145
rect -2930 5120 -2920 5145
rect -3075 5110 -2920 5120
rect -2220 5145 -2065 5155
rect -2220 5120 -2210 5145
rect -2190 5120 -2170 5145
rect -2150 5120 -2130 5145
rect -2110 5120 -2090 5145
rect -2220 5110 -2065 5120
rect -5595 5095 -3095 5105
rect -5595 5075 -5580 5095
rect -5550 5075 -5530 5095
rect -5510 5075 -5490 5095
rect -5470 5075 -5450 5095
rect -5430 5075 -5410 5095
rect -5390 5075 -5370 5095
rect -5350 5075 -5330 5095
rect -5310 5075 -5290 5095
rect -5270 5075 -5250 5095
rect -5230 5075 -5210 5095
rect -5190 5075 -5170 5095
rect -5150 5075 -5130 5095
rect -5110 5075 -5090 5095
rect -5070 5075 -5050 5095
rect -5030 5075 -5010 5095
rect -4990 5075 -4970 5095
rect -4950 5075 -4930 5095
rect -4910 5075 -4890 5095
rect -4870 5075 -4850 5095
rect -4830 5075 -4810 5095
rect -4790 5075 -4770 5095
rect -4750 5075 -4730 5095
rect -4710 5075 -4690 5095
rect -4670 5075 -4650 5095
rect -4630 5075 -4610 5095
rect -4590 5075 -4570 5095
rect -4550 5075 -4530 5095
rect -4510 5075 -4490 5095
rect -4470 5075 -4450 5095
rect -4430 5075 -4410 5095
rect -4390 5075 -4370 5095
rect -4350 5075 -4330 5095
rect -4310 5075 -4290 5095
rect -4270 5075 -4250 5095
rect -4230 5075 -4210 5095
rect -4190 5075 -4170 5095
rect -4150 5075 -4130 5095
rect -4110 5075 -4090 5095
rect -4070 5075 -4050 5095
rect -4030 5075 -4010 5095
rect -3990 5075 -3970 5095
rect -3950 5075 -3930 5095
rect -3910 5075 -3890 5095
rect -3870 5075 -3850 5095
rect -3830 5075 -3810 5095
rect -3790 5075 -3770 5095
rect -3750 5075 -3730 5095
rect -3710 5075 -3690 5095
rect -3670 5075 -3650 5095
rect -3630 5075 -3610 5095
rect -3590 5075 -3570 5095
rect -3550 5075 -3530 5095
rect -3510 5075 -3490 5095
rect -3470 5075 -3450 5095
rect -3430 5075 -3410 5095
rect -3390 5075 -3370 5095
rect -3350 5075 -3330 5095
rect -3310 5075 -3290 5095
rect -3270 5075 -3250 5095
rect -3230 5075 -3210 5095
rect -3190 5075 -3170 5095
rect -3150 5075 -3130 5095
rect -3110 5075 -3095 5095
rect -5595 5065 -3095 5075
rect -2045 5095 455 5105
rect -2045 5075 -2030 5095
rect -2010 5075 -1990 5095
rect -1970 5075 -1950 5095
rect -1930 5075 -1910 5095
rect -1890 5075 -1870 5095
rect -1850 5075 -1830 5095
rect -1810 5075 -1790 5095
rect -1770 5075 -1750 5095
rect -1730 5075 -1710 5095
rect -1690 5075 -1670 5095
rect -1650 5075 -1630 5095
rect -1610 5075 -1590 5095
rect -1570 5075 -1550 5095
rect -1530 5075 -1510 5095
rect -1490 5075 -1470 5095
rect -1450 5075 -1430 5095
rect -1410 5075 -1390 5095
rect -1370 5075 -1350 5095
rect -1330 5075 -1310 5095
rect -1290 5075 -1270 5095
rect -1250 5075 -1230 5095
rect -1210 5075 -1190 5095
rect -1170 5075 -1150 5095
rect -1130 5075 -1110 5095
rect -1090 5075 -1070 5095
rect -1050 5075 -1030 5095
rect -1010 5075 -990 5095
rect -970 5075 -950 5095
rect -930 5075 -910 5095
rect -890 5075 -870 5095
rect -850 5075 -830 5095
rect -810 5075 -790 5095
rect -770 5075 -750 5095
rect -730 5075 -710 5095
rect -690 5075 -670 5095
rect -650 5075 -630 5095
rect -610 5075 -590 5095
rect -570 5075 -550 5095
rect -530 5075 -510 5095
rect -490 5075 -470 5095
rect -450 5075 -430 5095
rect -410 5075 -390 5095
rect -370 5075 -350 5095
rect -330 5075 -310 5095
rect -290 5075 -270 5095
rect -250 5075 -230 5095
rect -210 5075 -190 5095
rect -170 5075 -150 5095
rect -130 5075 -110 5095
rect -90 5075 -70 5095
rect -50 5075 -30 5095
rect -10 5075 10 5095
rect 30 5075 50 5095
rect 70 5075 90 5095
rect 110 5075 130 5095
rect 150 5075 170 5095
rect 190 5075 210 5095
rect 230 5075 250 5095
rect 270 5075 290 5095
rect 310 5075 330 5095
rect 350 5075 370 5095
rect 390 5075 410 5095
rect 440 5075 455 5095
rect -2045 5065 455 5075
rect -3075 5050 -2920 5060
rect -3050 5025 -3030 5050
rect -3010 5025 -2990 5050
rect -2970 5025 -2950 5050
rect -2930 5025 -2920 5050
rect -3075 5015 -2920 5025
rect -2220 5050 -2065 5060
rect -2220 5025 -2210 5050
rect -2190 5025 -2170 5050
rect -2150 5025 -2130 5050
rect -2110 5025 -2090 5050
rect -2220 5015 -2065 5025
rect -5595 5000 -3095 5010
rect -5595 4980 -5580 5000
rect -5550 4980 -5530 5000
rect -5510 4980 -5490 5000
rect -5470 4980 -5450 5000
rect -5430 4980 -5410 5000
rect -5390 4980 -5370 5000
rect -5350 4980 -5330 5000
rect -5310 4980 -5290 5000
rect -5270 4980 -5250 5000
rect -5230 4980 -5210 5000
rect -5190 4980 -5170 5000
rect -5150 4980 -5130 5000
rect -5110 4980 -5090 5000
rect -5070 4980 -5050 5000
rect -5030 4980 -5010 5000
rect -4990 4980 -4970 5000
rect -4950 4980 -4930 5000
rect -4910 4980 -4890 5000
rect -4870 4980 -4850 5000
rect -4830 4980 -4810 5000
rect -4790 4980 -4770 5000
rect -4750 4980 -4730 5000
rect -4710 4980 -4690 5000
rect -4670 4980 -4650 5000
rect -4630 4980 -4610 5000
rect -4590 4980 -4570 5000
rect -4550 4980 -4530 5000
rect -4510 4980 -4490 5000
rect -4470 4980 -4450 5000
rect -4430 4980 -4410 5000
rect -4390 4980 -4370 5000
rect -4350 4980 -4330 5000
rect -4310 4980 -4290 5000
rect -4270 4980 -4250 5000
rect -4230 4980 -4210 5000
rect -4190 4980 -4170 5000
rect -4150 4980 -4130 5000
rect -4110 4980 -4090 5000
rect -4070 4980 -4050 5000
rect -4030 4980 -4010 5000
rect -3990 4980 -3970 5000
rect -3950 4980 -3930 5000
rect -3910 4980 -3890 5000
rect -3870 4980 -3850 5000
rect -3830 4980 -3810 5000
rect -3790 4980 -3770 5000
rect -3750 4980 -3730 5000
rect -3710 4980 -3690 5000
rect -3670 4980 -3650 5000
rect -3630 4980 -3610 5000
rect -3590 4980 -3570 5000
rect -3550 4980 -3530 5000
rect -3510 4980 -3490 5000
rect -3470 4980 -3450 5000
rect -3430 4980 -3410 5000
rect -3390 4980 -3370 5000
rect -3350 4980 -3330 5000
rect -3310 4980 -3290 5000
rect -3270 4980 -3250 5000
rect -3230 4980 -3210 5000
rect -3190 4980 -3170 5000
rect -3150 4980 -3130 5000
rect -3110 4980 -3095 5000
rect -5595 4970 -3095 4980
rect -2045 5000 455 5010
rect -2045 4980 -2030 5000
rect -2010 4980 -1990 5000
rect -1970 4980 -1950 5000
rect -1930 4980 -1910 5000
rect -1890 4980 -1870 5000
rect -1850 4980 -1830 5000
rect -1810 4980 -1790 5000
rect -1770 4980 -1750 5000
rect -1730 4980 -1710 5000
rect -1690 4980 -1670 5000
rect -1650 4980 -1630 5000
rect -1610 4980 -1590 5000
rect -1570 4980 -1550 5000
rect -1530 4980 -1510 5000
rect -1490 4980 -1470 5000
rect -1450 4980 -1430 5000
rect -1410 4980 -1390 5000
rect -1370 4980 -1350 5000
rect -1330 4980 -1310 5000
rect -1290 4980 -1270 5000
rect -1250 4980 -1230 5000
rect -1210 4980 -1190 5000
rect -1170 4980 -1150 5000
rect -1130 4980 -1110 5000
rect -1090 4980 -1070 5000
rect -1050 4980 -1030 5000
rect -1010 4980 -990 5000
rect -970 4980 -950 5000
rect -930 4980 -910 5000
rect -890 4980 -870 5000
rect -850 4980 -830 5000
rect -810 4980 -790 5000
rect -770 4980 -750 5000
rect -730 4980 -710 5000
rect -690 4980 -670 5000
rect -650 4980 -630 5000
rect -610 4980 -590 5000
rect -570 4980 -550 5000
rect -530 4980 -510 5000
rect -490 4980 -470 5000
rect -450 4980 -430 5000
rect -410 4980 -390 5000
rect -370 4980 -350 5000
rect -330 4980 -310 5000
rect -290 4980 -270 5000
rect -250 4980 -230 5000
rect -210 4980 -190 5000
rect -170 4980 -150 5000
rect -130 4980 -110 5000
rect -90 4980 -70 5000
rect -50 4980 -30 5000
rect -10 4980 10 5000
rect 30 4980 50 5000
rect 70 4980 90 5000
rect 110 4980 130 5000
rect 150 4980 170 5000
rect 190 4980 210 5000
rect 230 4980 250 5000
rect 270 4980 290 5000
rect 310 4980 330 5000
rect 350 4980 370 5000
rect 390 4980 410 5000
rect 440 4980 455 5000
rect -2045 4970 455 4980
rect -3075 4955 -2920 4965
rect -3050 4930 -3030 4955
rect -3010 4930 -2990 4955
rect -2970 4930 -2950 4955
rect -2930 4930 -2920 4955
rect -3075 4920 -2920 4930
rect -2220 4955 -2065 4965
rect -2220 4930 -2210 4955
rect -2190 4930 -2170 4955
rect -2150 4930 -2130 4955
rect -2110 4930 -2090 4955
rect -2220 4920 -2065 4930
rect -5595 4905 -3095 4915
rect -5595 4885 -5580 4905
rect -5550 4885 -5530 4905
rect -5510 4885 -5490 4905
rect -5470 4885 -5450 4905
rect -5430 4885 -5410 4905
rect -5390 4885 -5370 4905
rect -5350 4885 -5330 4905
rect -5310 4885 -5290 4905
rect -5270 4885 -5250 4905
rect -5230 4885 -5210 4905
rect -5190 4885 -5170 4905
rect -5150 4885 -5130 4905
rect -5110 4885 -5090 4905
rect -5070 4885 -5050 4905
rect -5030 4885 -5010 4905
rect -4990 4885 -4970 4905
rect -4950 4885 -4930 4905
rect -4910 4885 -4890 4905
rect -4870 4885 -4850 4905
rect -4830 4885 -4810 4905
rect -4790 4885 -4770 4905
rect -4750 4885 -4730 4905
rect -4710 4885 -4690 4905
rect -4670 4885 -4650 4905
rect -4630 4885 -4610 4905
rect -4590 4885 -4570 4905
rect -4550 4885 -4530 4905
rect -4510 4885 -4490 4905
rect -4470 4885 -4450 4905
rect -4430 4885 -4410 4905
rect -4390 4885 -4370 4905
rect -4350 4885 -4330 4905
rect -4310 4885 -4290 4905
rect -4270 4885 -4250 4905
rect -4230 4885 -4210 4905
rect -4190 4885 -4170 4905
rect -4150 4885 -4130 4905
rect -4110 4885 -4090 4905
rect -4070 4885 -4050 4905
rect -4030 4885 -4010 4905
rect -3990 4885 -3970 4905
rect -3950 4885 -3930 4905
rect -3910 4885 -3890 4905
rect -3870 4885 -3850 4905
rect -3830 4885 -3810 4905
rect -3790 4885 -3770 4905
rect -3750 4885 -3730 4905
rect -3710 4885 -3690 4905
rect -3670 4885 -3650 4905
rect -3630 4885 -3610 4905
rect -3590 4885 -3570 4905
rect -3550 4885 -3530 4905
rect -3510 4885 -3490 4905
rect -3470 4885 -3450 4905
rect -3430 4885 -3410 4905
rect -3390 4885 -3370 4905
rect -3350 4885 -3330 4905
rect -3310 4885 -3290 4905
rect -3270 4885 -3250 4905
rect -3230 4885 -3210 4905
rect -3190 4885 -3170 4905
rect -3150 4885 -3130 4905
rect -3110 4885 -3095 4905
rect -5595 4875 -3095 4885
rect -2045 4905 455 4915
rect -2045 4885 -2030 4905
rect -2010 4885 -1990 4905
rect -1970 4885 -1950 4905
rect -1930 4885 -1910 4905
rect -1890 4885 -1870 4905
rect -1850 4885 -1830 4905
rect -1810 4885 -1790 4905
rect -1770 4885 -1750 4905
rect -1730 4885 -1710 4905
rect -1690 4885 -1670 4905
rect -1650 4885 -1630 4905
rect -1610 4885 -1590 4905
rect -1570 4885 -1550 4905
rect -1530 4885 -1510 4905
rect -1490 4885 -1470 4905
rect -1450 4885 -1430 4905
rect -1410 4885 -1390 4905
rect -1370 4885 -1350 4905
rect -1330 4885 -1310 4905
rect -1290 4885 -1270 4905
rect -1250 4885 -1230 4905
rect -1210 4885 -1190 4905
rect -1170 4885 -1150 4905
rect -1130 4885 -1110 4905
rect -1090 4885 -1070 4905
rect -1050 4885 -1030 4905
rect -1010 4885 -990 4905
rect -970 4885 -950 4905
rect -930 4885 -910 4905
rect -890 4885 -870 4905
rect -850 4885 -830 4905
rect -810 4885 -790 4905
rect -770 4885 -750 4905
rect -730 4885 -710 4905
rect -690 4885 -670 4905
rect -650 4885 -630 4905
rect -610 4885 -590 4905
rect -570 4885 -550 4905
rect -530 4885 -510 4905
rect -490 4885 -470 4905
rect -450 4885 -430 4905
rect -410 4885 -390 4905
rect -370 4885 -350 4905
rect -330 4885 -310 4905
rect -290 4885 -270 4905
rect -250 4885 -230 4905
rect -210 4885 -190 4905
rect -170 4885 -150 4905
rect -130 4885 -110 4905
rect -90 4885 -70 4905
rect -50 4885 -30 4905
rect -10 4885 10 4905
rect 30 4885 50 4905
rect 70 4885 90 4905
rect 110 4885 130 4905
rect 150 4885 170 4905
rect 190 4885 210 4905
rect 230 4885 250 4905
rect 270 4885 290 4905
rect 310 4885 330 4905
rect 350 4885 370 4905
rect 390 4885 410 4905
rect 440 4885 455 4905
rect -2045 4875 455 4885
rect -3075 4860 -2920 4870
rect -3050 4835 -3030 4860
rect -3010 4835 -2990 4860
rect -2970 4835 -2950 4860
rect -2930 4835 -2920 4860
rect -3075 4825 -2920 4835
rect -2220 4860 -2065 4870
rect -2220 4835 -2210 4860
rect -2190 4835 -2170 4860
rect -2150 4835 -2130 4860
rect -2110 4835 -2090 4860
rect -2220 4825 -2065 4835
rect -5595 4810 -3095 4820
rect -5595 4790 -5580 4810
rect -5550 4790 -5530 4810
rect -5510 4790 -5490 4810
rect -5470 4790 -5450 4810
rect -5430 4790 -5410 4810
rect -5390 4790 -5370 4810
rect -5350 4790 -5330 4810
rect -5310 4790 -5290 4810
rect -5270 4790 -5250 4810
rect -5230 4790 -5210 4810
rect -5190 4790 -5170 4810
rect -5150 4790 -5130 4810
rect -5110 4790 -5090 4810
rect -5070 4790 -5050 4810
rect -5030 4790 -5010 4810
rect -4990 4790 -4970 4810
rect -4950 4790 -4930 4810
rect -4910 4790 -4890 4810
rect -4870 4790 -4850 4810
rect -4830 4790 -4810 4810
rect -4790 4790 -4770 4810
rect -4750 4790 -4730 4810
rect -4710 4790 -4690 4810
rect -4670 4790 -4650 4810
rect -4630 4790 -4610 4810
rect -4590 4790 -4570 4810
rect -4550 4790 -4530 4810
rect -4510 4790 -4490 4810
rect -4470 4790 -4450 4810
rect -4430 4790 -4410 4810
rect -4390 4790 -4370 4810
rect -4350 4790 -4330 4810
rect -4310 4790 -4290 4810
rect -4270 4790 -4250 4810
rect -4230 4790 -4210 4810
rect -4190 4790 -4170 4810
rect -4150 4790 -4130 4810
rect -4110 4790 -4090 4810
rect -4070 4790 -4050 4810
rect -4030 4790 -4010 4810
rect -3990 4790 -3970 4810
rect -3950 4790 -3930 4810
rect -3910 4790 -3890 4810
rect -3870 4790 -3850 4810
rect -3830 4790 -3810 4810
rect -3790 4790 -3770 4810
rect -3750 4790 -3730 4810
rect -3710 4790 -3690 4810
rect -3670 4790 -3650 4810
rect -3630 4790 -3610 4810
rect -3590 4790 -3570 4810
rect -3550 4790 -3530 4810
rect -3510 4790 -3490 4810
rect -3470 4790 -3450 4810
rect -3430 4790 -3410 4810
rect -3390 4790 -3370 4810
rect -3350 4790 -3330 4810
rect -3310 4790 -3290 4810
rect -3270 4790 -3250 4810
rect -3230 4790 -3210 4810
rect -3190 4790 -3170 4810
rect -3150 4790 -3130 4810
rect -3110 4790 -3095 4810
rect -5595 4780 -3095 4790
rect -2045 4810 455 4820
rect -2045 4790 -2030 4810
rect -2010 4790 -1990 4810
rect -1970 4790 -1950 4810
rect -1930 4790 -1910 4810
rect -1890 4790 -1870 4810
rect -1850 4790 -1830 4810
rect -1810 4790 -1790 4810
rect -1770 4790 -1750 4810
rect -1730 4790 -1710 4810
rect -1690 4790 -1670 4810
rect -1650 4790 -1630 4810
rect -1610 4790 -1590 4810
rect -1570 4790 -1550 4810
rect -1530 4790 -1510 4810
rect -1490 4790 -1470 4810
rect -1450 4790 -1430 4810
rect -1410 4790 -1390 4810
rect -1370 4790 -1350 4810
rect -1330 4790 -1310 4810
rect -1290 4790 -1270 4810
rect -1250 4790 -1230 4810
rect -1210 4790 -1190 4810
rect -1170 4790 -1150 4810
rect -1130 4790 -1110 4810
rect -1090 4790 -1070 4810
rect -1050 4790 -1030 4810
rect -1010 4790 -990 4810
rect -970 4790 -950 4810
rect -930 4790 -910 4810
rect -890 4790 -870 4810
rect -850 4790 -830 4810
rect -810 4790 -790 4810
rect -770 4790 -750 4810
rect -730 4790 -710 4810
rect -690 4790 -670 4810
rect -650 4790 -630 4810
rect -610 4790 -590 4810
rect -570 4790 -550 4810
rect -530 4790 -510 4810
rect -490 4790 -470 4810
rect -450 4790 -430 4810
rect -410 4790 -390 4810
rect -370 4790 -350 4810
rect -330 4790 -310 4810
rect -290 4790 -270 4810
rect -250 4790 -230 4810
rect -210 4790 -190 4810
rect -170 4790 -150 4810
rect -130 4790 -110 4810
rect -90 4790 -70 4810
rect -50 4790 -30 4810
rect -10 4790 10 4810
rect 30 4790 50 4810
rect 70 4790 90 4810
rect 110 4790 130 4810
rect 150 4790 170 4810
rect 190 4790 210 4810
rect 230 4790 250 4810
rect 270 4790 290 4810
rect 310 4790 330 4810
rect 350 4790 370 4810
rect 390 4790 410 4810
rect 440 4790 455 4810
rect -2045 4780 455 4790
rect -3075 4765 -2920 4775
rect -3050 4740 -3030 4765
rect -3010 4740 -2990 4765
rect -2970 4740 -2950 4765
rect -2930 4740 -2920 4765
rect -3075 4730 -2920 4740
rect -2220 4765 -2065 4775
rect -2220 4740 -2210 4765
rect -2190 4740 -2170 4765
rect -2150 4740 -2130 4765
rect -2110 4740 -2090 4765
rect -2220 4730 -2065 4740
rect -5595 4715 -3095 4725
rect -5595 4695 -5580 4715
rect -5550 4695 -5530 4715
rect -5510 4695 -5490 4715
rect -5470 4695 -5450 4715
rect -5430 4695 -5410 4715
rect -5390 4695 -5370 4715
rect -5350 4695 -5330 4715
rect -5310 4695 -5290 4715
rect -5270 4695 -5250 4715
rect -5230 4695 -5210 4715
rect -5190 4695 -5170 4715
rect -5150 4695 -5130 4715
rect -5110 4695 -5090 4715
rect -5070 4695 -5050 4715
rect -5030 4695 -5010 4715
rect -4990 4695 -4970 4715
rect -4950 4695 -4930 4715
rect -4910 4695 -4890 4715
rect -4870 4695 -4850 4715
rect -4830 4695 -4810 4715
rect -4790 4695 -4770 4715
rect -4750 4695 -4730 4715
rect -4710 4695 -4690 4715
rect -4670 4695 -4650 4715
rect -4630 4695 -4610 4715
rect -4590 4695 -4570 4715
rect -4550 4695 -4530 4715
rect -4510 4695 -4490 4715
rect -4470 4695 -4450 4715
rect -4430 4695 -4410 4715
rect -4390 4695 -4370 4715
rect -4350 4695 -4330 4715
rect -4310 4695 -4290 4715
rect -4270 4695 -4250 4715
rect -4230 4695 -4210 4715
rect -4190 4695 -4170 4715
rect -4150 4695 -4130 4715
rect -4110 4695 -4090 4715
rect -4070 4695 -4050 4715
rect -4030 4695 -4010 4715
rect -3990 4695 -3970 4715
rect -3950 4695 -3930 4715
rect -3910 4695 -3890 4715
rect -3870 4695 -3850 4715
rect -3830 4695 -3810 4715
rect -3790 4695 -3770 4715
rect -3750 4695 -3730 4715
rect -3710 4695 -3690 4715
rect -3670 4695 -3650 4715
rect -3630 4695 -3610 4715
rect -3590 4695 -3570 4715
rect -3550 4695 -3530 4715
rect -3510 4695 -3490 4715
rect -3470 4695 -3450 4715
rect -3430 4695 -3410 4715
rect -3390 4695 -3370 4715
rect -3350 4695 -3330 4715
rect -3310 4695 -3290 4715
rect -3270 4695 -3250 4715
rect -3230 4695 -3210 4715
rect -3190 4695 -3170 4715
rect -3150 4695 -3130 4715
rect -3110 4695 -3095 4715
rect -5595 4685 -3095 4695
rect -2045 4715 455 4725
rect -2045 4695 -2030 4715
rect -2010 4695 -1990 4715
rect -1970 4695 -1950 4715
rect -1930 4695 -1910 4715
rect -1890 4695 -1870 4715
rect -1850 4695 -1830 4715
rect -1810 4695 -1790 4715
rect -1770 4695 -1750 4715
rect -1730 4695 -1710 4715
rect -1690 4695 -1670 4715
rect -1650 4695 -1630 4715
rect -1610 4695 -1590 4715
rect -1570 4695 -1550 4715
rect -1530 4695 -1510 4715
rect -1490 4695 -1470 4715
rect -1450 4695 -1430 4715
rect -1410 4695 -1390 4715
rect -1370 4695 -1350 4715
rect -1330 4695 -1310 4715
rect -1290 4695 -1270 4715
rect -1250 4695 -1230 4715
rect -1210 4695 -1190 4715
rect -1170 4695 -1150 4715
rect -1130 4695 -1110 4715
rect -1090 4695 -1070 4715
rect -1050 4695 -1030 4715
rect -1010 4695 -990 4715
rect -970 4695 -950 4715
rect -930 4695 -910 4715
rect -890 4695 -870 4715
rect -850 4695 -830 4715
rect -810 4695 -790 4715
rect -770 4695 -750 4715
rect -730 4695 -710 4715
rect -690 4695 -670 4715
rect -650 4695 -630 4715
rect -610 4695 -590 4715
rect -570 4695 -550 4715
rect -530 4695 -510 4715
rect -490 4695 -470 4715
rect -450 4695 -430 4715
rect -410 4695 -390 4715
rect -370 4695 -350 4715
rect -330 4695 -310 4715
rect -290 4695 -270 4715
rect -250 4695 -230 4715
rect -210 4695 -190 4715
rect -170 4695 -150 4715
rect -130 4695 -110 4715
rect -90 4695 -70 4715
rect -50 4695 -30 4715
rect -10 4695 10 4715
rect 30 4695 50 4715
rect 70 4695 90 4715
rect 110 4695 130 4715
rect 150 4695 170 4715
rect 190 4695 210 4715
rect 230 4695 250 4715
rect 270 4695 290 4715
rect 310 4695 330 4715
rect 350 4695 370 4715
rect 390 4695 410 4715
rect 440 4695 455 4715
rect -2045 4685 455 4695
rect -3075 4670 -2920 4680
rect -3050 4645 -3030 4670
rect -3010 4645 -2990 4670
rect -2970 4645 -2950 4670
rect -2930 4645 -2920 4670
rect -3075 4635 -2920 4645
rect -2220 4670 -2065 4680
rect -2220 4645 -2210 4670
rect -2190 4645 -2170 4670
rect -2150 4645 -2130 4670
rect -2110 4645 -2090 4670
rect -2220 4635 -2065 4645
rect -5595 4620 -3095 4630
rect -5595 4600 -5580 4620
rect -5550 4600 -5530 4620
rect -5510 4600 -5490 4620
rect -5470 4600 -5450 4620
rect -5430 4600 -5410 4620
rect -5390 4600 -5370 4620
rect -5350 4600 -5330 4620
rect -5310 4600 -5290 4620
rect -5270 4600 -5250 4620
rect -5230 4600 -5210 4620
rect -5190 4600 -5170 4620
rect -5150 4600 -5130 4620
rect -5110 4600 -5090 4620
rect -5070 4600 -5050 4620
rect -5030 4600 -5010 4620
rect -4990 4600 -4970 4620
rect -4950 4600 -4930 4620
rect -4910 4600 -4890 4620
rect -4870 4600 -4850 4620
rect -4830 4600 -4810 4620
rect -4790 4600 -4770 4620
rect -4750 4600 -4730 4620
rect -4710 4600 -4690 4620
rect -4670 4600 -4650 4620
rect -4630 4600 -4610 4620
rect -4590 4600 -4570 4620
rect -4550 4600 -4530 4620
rect -4510 4600 -4490 4620
rect -4470 4600 -4450 4620
rect -4430 4600 -4410 4620
rect -4390 4600 -4370 4620
rect -4350 4600 -4330 4620
rect -4310 4600 -4290 4620
rect -4270 4600 -4250 4620
rect -4230 4600 -4210 4620
rect -4190 4600 -4170 4620
rect -4150 4600 -4130 4620
rect -4110 4600 -4090 4620
rect -4070 4600 -4050 4620
rect -4030 4600 -4010 4620
rect -3990 4600 -3970 4620
rect -3950 4600 -3930 4620
rect -3910 4600 -3890 4620
rect -3870 4600 -3850 4620
rect -3830 4600 -3810 4620
rect -3790 4600 -3770 4620
rect -3750 4600 -3730 4620
rect -3710 4600 -3690 4620
rect -3670 4600 -3650 4620
rect -3630 4600 -3610 4620
rect -3590 4600 -3570 4620
rect -3550 4600 -3530 4620
rect -3510 4600 -3490 4620
rect -3470 4600 -3450 4620
rect -3430 4600 -3410 4620
rect -3390 4600 -3370 4620
rect -3350 4600 -3330 4620
rect -3310 4600 -3290 4620
rect -3270 4600 -3250 4620
rect -3230 4600 -3210 4620
rect -3190 4600 -3170 4620
rect -3150 4600 -3130 4620
rect -3110 4600 -3095 4620
rect -5595 4590 -3095 4600
rect -2045 4620 455 4630
rect -2045 4600 -2030 4620
rect -2010 4600 -1990 4620
rect -1970 4600 -1950 4620
rect -1930 4600 -1910 4620
rect -1890 4600 -1870 4620
rect -1850 4600 -1830 4620
rect -1810 4600 -1790 4620
rect -1770 4600 -1750 4620
rect -1730 4600 -1710 4620
rect -1690 4600 -1670 4620
rect -1650 4600 -1630 4620
rect -1610 4600 -1590 4620
rect -1570 4600 -1550 4620
rect -1530 4600 -1510 4620
rect -1490 4600 -1470 4620
rect -1450 4600 -1430 4620
rect -1410 4600 -1390 4620
rect -1370 4600 -1350 4620
rect -1330 4600 -1310 4620
rect -1290 4600 -1270 4620
rect -1250 4600 -1230 4620
rect -1210 4600 -1190 4620
rect -1170 4600 -1150 4620
rect -1130 4600 -1110 4620
rect -1090 4600 -1070 4620
rect -1050 4600 -1030 4620
rect -1010 4600 -990 4620
rect -970 4600 -950 4620
rect -930 4600 -910 4620
rect -890 4600 -870 4620
rect -850 4600 -830 4620
rect -810 4600 -790 4620
rect -770 4600 -750 4620
rect -730 4600 -710 4620
rect -690 4600 -670 4620
rect -650 4600 -630 4620
rect -610 4600 -590 4620
rect -570 4600 -550 4620
rect -530 4600 -510 4620
rect -490 4600 -470 4620
rect -450 4600 -430 4620
rect -410 4600 -390 4620
rect -370 4600 -350 4620
rect -330 4600 -310 4620
rect -290 4600 -270 4620
rect -250 4600 -230 4620
rect -210 4600 -190 4620
rect -170 4600 -150 4620
rect -130 4600 -110 4620
rect -90 4600 -70 4620
rect -50 4600 -30 4620
rect -10 4600 10 4620
rect 30 4600 50 4620
rect 70 4600 90 4620
rect 110 4600 130 4620
rect 150 4600 170 4620
rect 190 4600 210 4620
rect 230 4600 250 4620
rect 270 4600 290 4620
rect 310 4600 330 4620
rect 350 4600 370 4620
rect 390 4600 410 4620
rect 440 4600 455 4620
rect -2045 4590 455 4600
rect -3075 4575 -2920 4585
rect -3050 4550 -3030 4575
rect -3010 4550 -2990 4575
rect -2970 4550 -2950 4575
rect -2930 4550 -2920 4575
rect -3075 4540 -2920 4550
rect -2220 4575 -2065 4585
rect -2220 4550 -2210 4575
rect -2190 4550 -2170 4575
rect -2150 4550 -2130 4575
rect -2110 4550 -2090 4575
rect -2220 4540 -2065 4550
rect -5595 4525 -3095 4535
rect -5595 4505 -5580 4525
rect -5550 4505 -5530 4525
rect -5510 4505 -5490 4525
rect -5470 4505 -5450 4525
rect -5430 4505 -5410 4525
rect -5390 4505 -5370 4525
rect -5350 4505 -5330 4525
rect -5310 4505 -5290 4525
rect -5270 4505 -5250 4525
rect -5230 4505 -5210 4525
rect -5190 4505 -5170 4525
rect -5150 4505 -5130 4525
rect -5110 4505 -5090 4525
rect -5070 4505 -5050 4525
rect -5030 4505 -5010 4525
rect -4990 4505 -4970 4525
rect -4950 4505 -4930 4525
rect -4910 4505 -4890 4525
rect -4870 4505 -4850 4525
rect -4830 4505 -4810 4525
rect -4790 4505 -4770 4525
rect -4750 4505 -4730 4525
rect -4710 4505 -4690 4525
rect -4670 4505 -4650 4525
rect -4630 4505 -4610 4525
rect -4590 4505 -4570 4525
rect -4550 4505 -4530 4525
rect -4510 4505 -4490 4525
rect -4470 4505 -4450 4525
rect -4430 4505 -4410 4525
rect -4390 4505 -4370 4525
rect -4350 4505 -4330 4525
rect -4310 4505 -4290 4525
rect -4270 4505 -4250 4525
rect -4230 4505 -4210 4525
rect -4190 4505 -4170 4525
rect -4150 4505 -4130 4525
rect -4110 4505 -4090 4525
rect -4070 4505 -4050 4525
rect -4030 4505 -4010 4525
rect -3990 4505 -3970 4525
rect -3950 4505 -3930 4525
rect -3910 4505 -3890 4525
rect -3870 4505 -3850 4525
rect -3830 4505 -3810 4525
rect -3790 4505 -3770 4525
rect -3750 4505 -3730 4525
rect -3710 4505 -3690 4525
rect -3670 4505 -3650 4525
rect -3630 4505 -3610 4525
rect -3590 4505 -3570 4525
rect -3550 4505 -3530 4525
rect -3510 4505 -3490 4525
rect -3470 4505 -3450 4525
rect -3430 4505 -3410 4525
rect -3390 4505 -3370 4525
rect -3350 4505 -3330 4525
rect -3310 4505 -3290 4525
rect -3270 4505 -3250 4525
rect -3230 4505 -3210 4525
rect -3190 4505 -3170 4525
rect -3150 4505 -3130 4525
rect -3110 4505 -3095 4525
rect -5595 4495 -3095 4505
rect -2045 4525 455 4535
rect -2045 4505 -2030 4525
rect -2010 4505 -1990 4525
rect -1970 4505 -1950 4525
rect -1930 4505 -1910 4525
rect -1890 4505 -1870 4525
rect -1850 4505 -1830 4525
rect -1810 4505 -1790 4525
rect -1770 4505 -1750 4525
rect -1730 4505 -1710 4525
rect -1690 4505 -1670 4525
rect -1650 4505 -1630 4525
rect -1610 4505 -1590 4525
rect -1570 4505 -1550 4525
rect -1530 4505 -1510 4525
rect -1490 4505 -1470 4525
rect -1450 4505 -1430 4525
rect -1410 4505 -1390 4525
rect -1370 4505 -1350 4525
rect -1330 4505 -1310 4525
rect -1290 4505 -1270 4525
rect -1250 4505 -1230 4525
rect -1210 4505 -1190 4525
rect -1170 4505 -1150 4525
rect -1130 4505 -1110 4525
rect -1090 4505 -1070 4525
rect -1050 4505 -1030 4525
rect -1010 4505 -990 4525
rect -970 4505 -950 4525
rect -930 4505 -910 4525
rect -890 4505 -870 4525
rect -850 4505 -830 4525
rect -810 4505 -790 4525
rect -770 4505 -750 4525
rect -730 4505 -710 4525
rect -690 4505 -670 4525
rect -650 4505 -630 4525
rect -610 4505 -590 4525
rect -570 4505 -550 4525
rect -530 4505 -510 4525
rect -490 4505 -470 4525
rect -450 4505 -430 4525
rect -410 4505 -390 4525
rect -370 4505 -350 4525
rect -330 4505 -310 4525
rect -290 4505 -270 4525
rect -250 4505 -230 4525
rect -210 4505 -190 4525
rect -170 4505 -150 4525
rect -130 4505 -110 4525
rect -90 4505 -70 4525
rect -50 4505 -30 4525
rect -10 4505 10 4525
rect 30 4505 50 4525
rect 70 4505 90 4525
rect 110 4505 130 4525
rect 150 4505 170 4525
rect 190 4505 210 4525
rect 230 4505 250 4525
rect 270 4505 290 4525
rect 310 4505 330 4525
rect 350 4505 370 4525
rect 390 4505 410 4525
rect 440 4505 455 4525
rect -2045 4495 455 4505
rect -3075 4480 -2920 4490
rect -3050 4455 -3030 4480
rect -3010 4455 -2990 4480
rect -2970 4455 -2950 4480
rect -2930 4455 -2920 4480
rect -3075 4445 -2920 4455
rect -2220 4480 -2065 4490
rect -2220 4455 -2210 4480
rect -2190 4455 -2170 4480
rect -2150 4455 -2130 4480
rect -2110 4455 -2090 4480
rect -2220 4445 -2065 4455
rect -5595 4430 -3095 4440
rect -5595 4410 -5580 4430
rect -5550 4410 -5530 4430
rect -5510 4410 -5490 4430
rect -5470 4410 -5450 4430
rect -5430 4410 -5410 4430
rect -5390 4410 -5370 4430
rect -5350 4410 -5330 4430
rect -5310 4410 -5290 4430
rect -5270 4410 -5250 4430
rect -5230 4410 -5210 4430
rect -5190 4410 -5170 4430
rect -5150 4410 -5130 4430
rect -5110 4410 -5090 4430
rect -5070 4410 -5050 4430
rect -5030 4410 -5010 4430
rect -4990 4410 -4970 4430
rect -4950 4410 -4930 4430
rect -4910 4410 -4890 4430
rect -4870 4410 -4850 4430
rect -4830 4410 -4810 4430
rect -4790 4410 -4770 4430
rect -4750 4410 -4730 4430
rect -4710 4410 -4690 4430
rect -4670 4410 -4650 4430
rect -4630 4410 -4610 4430
rect -4590 4410 -4570 4430
rect -4550 4410 -4530 4430
rect -4510 4410 -4490 4430
rect -4470 4410 -4450 4430
rect -4430 4410 -4410 4430
rect -4390 4410 -4370 4430
rect -4350 4410 -4330 4430
rect -4310 4410 -4290 4430
rect -4270 4410 -4250 4430
rect -4230 4410 -4210 4430
rect -4190 4410 -4170 4430
rect -4150 4410 -4130 4430
rect -4110 4410 -4090 4430
rect -4070 4410 -4050 4430
rect -4030 4410 -4010 4430
rect -3990 4410 -3970 4430
rect -3950 4410 -3930 4430
rect -3910 4410 -3890 4430
rect -3870 4410 -3850 4430
rect -3830 4410 -3810 4430
rect -3790 4410 -3770 4430
rect -3750 4410 -3730 4430
rect -3710 4410 -3690 4430
rect -3670 4410 -3650 4430
rect -3630 4410 -3610 4430
rect -3590 4410 -3570 4430
rect -3550 4410 -3530 4430
rect -3510 4410 -3490 4430
rect -3470 4410 -3450 4430
rect -3430 4410 -3410 4430
rect -3390 4410 -3370 4430
rect -3350 4410 -3330 4430
rect -3310 4410 -3290 4430
rect -3270 4410 -3250 4430
rect -3230 4410 -3210 4430
rect -3190 4410 -3170 4430
rect -3150 4410 -3130 4430
rect -3110 4410 -3095 4430
rect -5595 4400 -3095 4410
rect -2045 4430 455 4440
rect -2045 4410 -2030 4430
rect -2010 4410 -1990 4430
rect -1970 4410 -1950 4430
rect -1930 4410 -1910 4430
rect -1890 4410 -1870 4430
rect -1850 4410 -1830 4430
rect -1810 4410 -1790 4430
rect -1770 4410 -1750 4430
rect -1730 4410 -1710 4430
rect -1690 4410 -1670 4430
rect -1650 4410 -1630 4430
rect -1610 4410 -1590 4430
rect -1570 4410 -1550 4430
rect -1530 4410 -1510 4430
rect -1490 4410 -1470 4430
rect -1450 4410 -1430 4430
rect -1410 4410 -1390 4430
rect -1370 4410 -1350 4430
rect -1330 4410 -1310 4430
rect -1290 4410 -1270 4430
rect -1250 4410 -1230 4430
rect -1210 4410 -1190 4430
rect -1170 4410 -1150 4430
rect -1130 4410 -1110 4430
rect -1090 4410 -1070 4430
rect -1050 4410 -1030 4430
rect -1010 4410 -990 4430
rect -970 4410 -950 4430
rect -930 4410 -910 4430
rect -890 4410 -870 4430
rect -850 4410 -830 4430
rect -810 4410 -790 4430
rect -770 4410 -750 4430
rect -730 4410 -710 4430
rect -690 4410 -670 4430
rect -650 4410 -630 4430
rect -610 4410 -590 4430
rect -570 4410 -550 4430
rect -530 4410 -510 4430
rect -490 4410 -470 4430
rect -450 4410 -430 4430
rect -410 4410 -390 4430
rect -370 4410 -350 4430
rect -330 4410 -310 4430
rect -290 4410 -270 4430
rect -250 4410 -230 4430
rect -210 4410 -190 4430
rect -170 4410 -150 4430
rect -130 4410 -110 4430
rect -90 4410 -70 4430
rect -50 4410 -30 4430
rect -10 4410 10 4430
rect 30 4410 50 4430
rect 70 4410 90 4430
rect 110 4410 130 4430
rect 150 4410 170 4430
rect 190 4410 210 4430
rect 230 4410 250 4430
rect 270 4410 290 4430
rect 310 4410 330 4430
rect 350 4410 370 4430
rect 390 4410 410 4430
rect 440 4410 455 4430
rect -2045 4400 455 4410
rect -3075 4385 -2920 4395
rect -3050 4360 -3030 4385
rect -3010 4360 -2990 4385
rect -2970 4360 -2950 4385
rect -2930 4360 -2920 4385
rect -3075 4350 -2920 4360
rect -2220 4385 -2065 4395
rect -2220 4360 -2210 4385
rect -2190 4360 -2170 4385
rect -2150 4360 -2130 4385
rect -2110 4360 -2090 4385
rect -2220 4350 -2065 4360
rect -5595 4335 -3095 4345
rect -5595 4315 -5580 4335
rect -5550 4315 -5530 4335
rect -5510 4315 -5490 4335
rect -5470 4315 -5450 4335
rect -5430 4315 -5410 4335
rect -5390 4315 -5370 4335
rect -5350 4315 -5330 4335
rect -5310 4315 -5290 4335
rect -5270 4315 -5250 4335
rect -5230 4315 -5210 4335
rect -5190 4315 -5170 4335
rect -5150 4315 -5130 4335
rect -5110 4315 -5090 4335
rect -5070 4315 -5050 4335
rect -5030 4315 -5010 4335
rect -4990 4315 -4970 4335
rect -4950 4315 -4930 4335
rect -4910 4315 -4890 4335
rect -4870 4315 -4850 4335
rect -4830 4315 -4810 4335
rect -4790 4315 -4770 4335
rect -4750 4315 -4730 4335
rect -4710 4315 -4690 4335
rect -4670 4315 -4650 4335
rect -4630 4315 -4610 4335
rect -4590 4315 -4570 4335
rect -4550 4315 -4530 4335
rect -4510 4315 -4490 4335
rect -4470 4315 -4450 4335
rect -4430 4315 -4410 4335
rect -4390 4315 -4370 4335
rect -4350 4315 -4330 4335
rect -4310 4315 -4290 4335
rect -4270 4315 -4250 4335
rect -4230 4315 -4210 4335
rect -4190 4315 -4170 4335
rect -4150 4315 -4130 4335
rect -4110 4315 -4090 4335
rect -4070 4315 -4050 4335
rect -4030 4315 -4010 4335
rect -3990 4315 -3970 4335
rect -3950 4315 -3930 4335
rect -3910 4315 -3890 4335
rect -3870 4315 -3850 4335
rect -3830 4315 -3810 4335
rect -3790 4315 -3770 4335
rect -3750 4315 -3730 4335
rect -3710 4315 -3690 4335
rect -3670 4315 -3650 4335
rect -3630 4315 -3610 4335
rect -3590 4315 -3570 4335
rect -3550 4315 -3530 4335
rect -3510 4315 -3490 4335
rect -3470 4315 -3450 4335
rect -3430 4315 -3410 4335
rect -3390 4315 -3370 4335
rect -3350 4315 -3330 4335
rect -3310 4315 -3290 4335
rect -3270 4315 -3250 4335
rect -3230 4315 -3210 4335
rect -3190 4315 -3170 4335
rect -3150 4315 -3130 4335
rect -3110 4315 -3095 4335
rect -5595 4305 -3095 4315
rect -2045 4335 455 4345
rect -2045 4315 -2030 4335
rect -2010 4315 -1990 4335
rect -1970 4315 -1950 4335
rect -1930 4315 -1910 4335
rect -1890 4315 -1870 4335
rect -1850 4315 -1830 4335
rect -1810 4315 -1790 4335
rect -1770 4315 -1750 4335
rect -1730 4315 -1710 4335
rect -1690 4315 -1670 4335
rect -1650 4315 -1630 4335
rect -1610 4315 -1590 4335
rect -1570 4315 -1550 4335
rect -1530 4315 -1510 4335
rect -1490 4315 -1470 4335
rect -1450 4315 -1430 4335
rect -1410 4315 -1390 4335
rect -1370 4315 -1350 4335
rect -1330 4315 -1310 4335
rect -1290 4315 -1270 4335
rect -1250 4315 -1230 4335
rect -1210 4315 -1190 4335
rect -1170 4315 -1150 4335
rect -1130 4315 -1110 4335
rect -1090 4315 -1070 4335
rect -1050 4315 -1030 4335
rect -1010 4315 -990 4335
rect -970 4315 -950 4335
rect -930 4315 -910 4335
rect -890 4315 -870 4335
rect -850 4315 -830 4335
rect -810 4315 -790 4335
rect -770 4315 -750 4335
rect -730 4315 -710 4335
rect -690 4315 -670 4335
rect -650 4315 -630 4335
rect -610 4315 -590 4335
rect -570 4315 -550 4335
rect -530 4315 -510 4335
rect -490 4315 -470 4335
rect -450 4315 -430 4335
rect -410 4315 -390 4335
rect -370 4315 -350 4335
rect -330 4315 -310 4335
rect -290 4315 -270 4335
rect -250 4315 -230 4335
rect -210 4315 -190 4335
rect -170 4315 -150 4335
rect -130 4315 -110 4335
rect -90 4315 -70 4335
rect -50 4315 -30 4335
rect -10 4315 10 4335
rect 30 4315 50 4335
rect 70 4315 90 4335
rect 110 4315 130 4335
rect 150 4315 170 4335
rect 190 4315 210 4335
rect 230 4315 250 4335
rect 270 4315 290 4335
rect 310 4315 330 4335
rect 350 4315 370 4335
rect 390 4315 410 4335
rect 440 4315 455 4335
rect -2045 4305 455 4315
rect -3075 4290 -2920 4300
rect -3050 4265 -3030 4290
rect -3010 4265 -2990 4290
rect -2970 4265 -2950 4290
rect -2930 4265 -2920 4290
rect -3075 4255 -2920 4265
rect -2220 4290 -2065 4300
rect -2220 4265 -2210 4290
rect -2190 4265 -2170 4290
rect -2150 4265 -2130 4290
rect -2110 4265 -2090 4290
rect -2220 4255 -2065 4265
rect -5595 4240 -3095 4250
rect -5595 4220 -5580 4240
rect -5550 4220 -5530 4240
rect -5510 4220 -5490 4240
rect -5470 4220 -5450 4240
rect -5430 4220 -5410 4240
rect -5390 4220 -5370 4240
rect -5350 4220 -5330 4240
rect -5310 4220 -5290 4240
rect -5270 4220 -5250 4240
rect -5230 4220 -5210 4240
rect -5190 4220 -5170 4240
rect -5150 4220 -5130 4240
rect -5110 4220 -5090 4240
rect -5070 4220 -5050 4240
rect -5030 4220 -5010 4240
rect -4990 4220 -4970 4240
rect -4950 4220 -4930 4240
rect -4910 4220 -4890 4240
rect -4870 4220 -4850 4240
rect -4830 4220 -4810 4240
rect -4790 4220 -4770 4240
rect -4750 4220 -4730 4240
rect -4710 4220 -4690 4240
rect -4670 4220 -4650 4240
rect -4630 4220 -4610 4240
rect -4590 4220 -4570 4240
rect -4550 4220 -4530 4240
rect -4510 4220 -4490 4240
rect -4470 4220 -4450 4240
rect -4430 4220 -4410 4240
rect -4390 4220 -4370 4240
rect -4350 4220 -4330 4240
rect -4310 4220 -4290 4240
rect -4270 4220 -4250 4240
rect -4230 4220 -4210 4240
rect -4190 4220 -4170 4240
rect -4150 4220 -4130 4240
rect -4110 4220 -4090 4240
rect -4070 4220 -4050 4240
rect -4030 4220 -4010 4240
rect -3990 4220 -3970 4240
rect -3950 4220 -3930 4240
rect -3910 4220 -3890 4240
rect -3870 4220 -3850 4240
rect -3830 4220 -3810 4240
rect -3790 4220 -3770 4240
rect -3750 4220 -3730 4240
rect -3710 4220 -3690 4240
rect -3670 4220 -3650 4240
rect -3630 4220 -3610 4240
rect -3590 4220 -3570 4240
rect -3550 4220 -3530 4240
rect -3510 4220 -3490 4240
rect -3470 4220 -3450 4240
rect -3430 4220 -3410 4240
rect -3390 4220 -3370 4240
rect -3350 4220 -3330 4240
rect -3310 4220 -3290 4240
rect -3270 4220 -3250 4240
rect -3230 4220 -3210 4240
rect -3190 4220 -3170 4240
rect -3150 4220 -3130 4240
rect -3110 4220 -3095 4240
rect -5595 4210 -3095 4220
rect -2045 4240 455 4250
rect -2045 4220 -2030 4240
rect -2010 4220 -1990 4240
rect -1970 4220 -1950 4240
rect -1930 4220 -1910 4240
rect -1890 4220 -1870 4240
rect -1850 4220 -1830 4240
rect -1810 4220 -1790 4240
rect -1770 4220 -1750 4240
rect -1730 4220 -1710 4240
rect -1690 4220 -1670 4240
rect -1650 4220 -1630 4240
rect -1610 4220 -1590 4240
rect -1570 4220 -1550 4240
rect -1530 4220 -1510 4240
rect -1490 4220 -1470 4240
rect -1450 4220 -1430 4240
rect -1410 4220 -1390 4240
rect -1370 4220 -1350 4240
rect -1330 4220 -1310 4240
rect -1290 4220 -1270 4240
rect -1250 4220 -1230 4240
rect -1210 4220 -1190 4240
rect -1170 4220 -1150 4240
rect -1130 4220 -1110 4240
rect -1090 4220 -1070 4240
rect -1050 4220 -1030 4240
rect -1010 4220 -990 4240
rect -970 4220 -950 4240
rect -930 4220 -910 4240
rect -890 4220 -870 4240
rect -850 4220 -830 4240
rect -810 4220 -790 4240
rect -770 4220 -750 4240
rect -730 4220 -710 4240
rect -690 4220 -670 4240
rect -650 4220 -630 4240
rect -610 4220 -590 4240
rect -570 4220 -550 4240
rect -530 4220 -510 4240
rect -490 4220 -470 4240
rect -450 4220 -430 4240
rect -410 4220 -390 4240
rect -370 4220 -350 4240
rect -330 4220 -310 4240
rect -290 4220 -270 4240
rect -250 4220 -230 4240
rect -210 4220 -190 4240
rect -170 4220 -150 4240
rect -130 4220 -110 4240
rect -90 4220 -70 4240
rect -50 4220 -30 4240
rect -10 4220 10 4240
rect 30 4220 50 4240
rect 70 4220 90 4240
rect 110 4220 130 4240
rect 150 4220 170 4240
rect 190 4220 210 4240
rect 230 4220 250 4240
rect 270 4220 290 4240
rect 310 4220 330 4240
rect 350 4220 370 4240
rect 390 4220 410 4240
rect 440 4220 455 4240
rect -2045 4210 455 4220
rect -3075 4195 -2920 4205
rect -3050 4170 -3030 4195
rect -3010 4170 -2990 4195
rect -2970 4170 -2950 4195
rect -2930 4170 -2920 4195
rect -3075 4160 -2920 4170
rect -2220 4195 -2065 4205
rect -2220 4170 -2210 4195
rect -2190 4170 -2170 4195
rect -2150 4170 -2130 4195
rect -2110 4170 -2090 4195
rect -2220 4160 -2065 4170
rect -5595 4145 -3095 4155
rect -5595 4125 -5580 4145
rect -5550 4125 -5530 4145
rect -5510 4125 -5490 4145
rect -5470 4125 -5450 4145
rect -5430 4125 -5410 4145
rect -5390 4125 -5370 4145
rect -5350 4125 -5330 4145
rect -5310 4125 -5290 4145
rect -5270 4125 -5250 4145
rect -5230 4125 -5210 4145
rect -5190 4125 -5170 4145
rect -5150 4125 -5130 4145
rect -5110 4125 -5090 4145
rect -5070 4125 -5050 4145
rect -5030 4125 -5010 4145
rect -4990 4125 -4970 4145
rect -4950 4125 -4930 4145
rect -4910 4125 -4890 4145
rect -4870 4125 -4850 4145
rect -4830 4125 -4810 4145
rect -4790 4125 -4770 4145
rect -4750 4125 -4730 4145
rect -4710 4125 -4690 4145
rect -4670 4125 -4650 4145
rect -4630 4125 -4610 4145
rect -4590 4125 -4570 4145
rect -4550 4125 -4530 4145
rect -4510 4125 -4490 4145
rect -4470 4125 -4450 4145
rect -4430 4125 -4410 4145
rect -4390 4125 -4370 4145
rect -4350 4125 -4330 4145
rect -4310 4125 -4290 4145
rect -4270 4125 -4250 4145
rect -4230 4125 -4210 4145
rect -4190 4125 -4170 4145
rect -4150 4125 -4130 4145
rect -4110 4125 -4090 4145
rect -4070 4125 -4050 4145
rect -4030 4125 -4010 4145
rect -3990 4125 -3970 4145
rect -3950 4125 -3930 4145
rect -3910 4125 -3890 4145
rect -3870 4125 -3850 4145
rect -3830 4125 -3810 4145
rect -3790 4125 -3770 4145
rect -3750 4125 -3730 4145
rect -3710 4125 -3690 4145
rect -3670 4125 -3650 4145
rect -3630 4125 -3610 4145
rect -3590 4125 -3570 4145
rect -3550 4125 -3530 4145
rect -3510 4125 -3490 4145
rect -3470 4125 -3450 4145
rect -3430 4125 -3410 4145
rect -3390 4125 -3370 4145
rect -3350 4125 -3330 4145
rect -3310 4125 -3290 4145
rect -3270 4125 -3250 4145
rect -3230 4125 -3210 4145
rect -3190 4125 -3170 4145
rect -3150 4125 -3130 4145
rect -3110 4125 -3095 4145
rect -5595 4115 -3095 4125
rect -2045 4145 455 4155
rect -2045 4125 -2030 4145
rect -2010 4125 -1990 4145
rect -1970 4125 -1950 4145
rect -1930 4125 -1910 4145
rect -1890 4125 -1870 4145
rect -1850 4125 -1830 4145
rect -1810 4125 -1790 4145
rect -1770 4125 -1750 4145
rect -1730 4125 -1710 4145
rect -1690 4125 -1670 4145
rect -1650 4125 -1630 4145
rect -1610 4125 -1590 4145
rect -1570 4125 -1550 4145
rect -1530 4125 -1510 4145
rect -1490 4125 -1470 4145
rect -1450 4125 -1430 4145
rect -1410 4125 -1390 4145
rect -1370 4125 -1350 4145
rect -1330 4125 -1310 4145
rect -1290 4125 -1270 4145
rect -1250 4125 -1230 4145
rect -1210 4125 -1190 4145
rect -1170 4125 -1150 4145
rect -1130 4125 -1110 4145
rect -1090 4125 -1070 4145
rect -1050 4125 -1030 4145
rect -1010 4125 -990 4145
rect -970 4125 -950 4145
rect -930 4125 -910 4145
rect -890 4125 -870 4145
rect -850 4125 -830 4145
rect -810 4125 -790 4145
rect -770 4125 -750 4145
rect -730 4125 -710 4145
rect -690 4125 -670 4145
rect -650 4125 -630 4145
rect -610 4125 -590 4145
rect -570 4125 -550 4145
rect -530 4125 -510 4145
rect -490 4125 -470 4145
rect -450 4125 -430 4145
rect -410 4125 -390 4145
rect -370 4125 -350 4145
rect -330 4125 -310 4145
rect -290 4125 -270 4145
rect -250 4125 -230 4145
rect -210 4125 -190 4145
rect -170 4125 -150 4145
rect -130 4125 -110 4145
rect -90 4125 -70 4145
rect -50 4125 -30 4145
rect -10 4125 10 4145
rect 30 4125 50 4145
rect 70 4125 90 4145
rect 110 4125 130 4145
rect 150 4125 170 4145
rect 190 4125 210 4145
rect 230 4125 250 4145
rect 270 4125 290 4145
rect 310 4125 330 4145
rect 350 4125 370 4145
rect 390 4125 410 4145
rect 440 4125 455 4145
rect -2045 4115 455 4125
rect -3075 4100 -2920 4110
rect -3050 4075 -3030 4100
rect -3010 4075 -2990 4100
rect -2970 4075 -2950 4100
rect -2930 4075 -2920 4100
rect -3075 4065 -2920 4075
rect -2220 4100 -2065 4110
rect -2220 4075 -2210 4100
rect -2190 4075 -2170 4100
rect -2150 4075 -2130 4100
rect -2110 4075 -2090 4100
rect -2220 4065 -2065 4075
rect -5595 4050 -3095 4060
rect -5595 4030 -5580 4050
rect -5550 4030 -5530 4050
rect -5510 4030 -5490 4050
rect -5470 4030 -5450 4050
rect -5430 4030 -5410 4050
rect -5390 4030 -5370 4050
rect -5350 4030 -5330 4050
rect -5310 4030 -5290 4050
rect -5270 4030 -5250 4050
rect -5230 4030 -5210 4050
rect -5190 4030 -5170 4050
rect -5150 4030 -5130 4050
rect -5110 4030 -5090 4050
rect -5070 4030 -5050 4050
rect -5030 4030 -5010 4050
rect -4990 4030 -4970 4050
rect -4950 4030 -4930 4050
rect -4910 4030 -4890 4050
rect -4870 4030 -4850 4050
rect -4830 4030 -4810 4050
rect -4790 4030 -4770 4050
rect -4750 4030 -4730 4050
rect -4710 4030 -4690 4050
rect -4670 4030 -4650 4050
rect -4630 4030 -4610 4050
rect -4590 4030 -4570 4050
rect -4550 4030 -4530 4050
rect -4510 4030 -4490 4050
rect -4470 4030 -4450 4050
rect -4430 4030 -4410 4050
rect -4390 4030 -4370 4050
rect -4350 4030 -4330 4050
rect -4310 4030 -4290 4050
rect -4270 4030 -4250 4050
rect -4230 4030 -4210 4050
rect -4190 4030 -4170 4050
rect -4150 4030 -4130 4050
rect -4110 4030 -4090 4050
rect -4070 4030 -4050 4050
rect -4030 4030 -4010 4050
rect -3990 4030 -3970 4050
rect -3950 4030 -3930 4050
rect -3910 4030 -3890 4050
rect -3870 4030 -3850 4050
rect -3830 4030 -3810 4050
rect -3790 4030 -3770 4050
rect -3750 4030 -3730 4050
rect -3710 4030 -3690 4050
rect -3670 4030 -3650 4050
rect -3630 4030 -3610 4050
rect -3590 4030 -3570 4050
rect -3550 4030 -3530 4050
rect -3510 4030 -3490 4050
rect -3470 4030 -3450 4050
rect -3430 4030 -3410 4050
rect -3390 4030 -3370 4050
rect -3350 4030 -3330 4050
rect -3310 4030 -3290 4050
rect -3270 4030 -3250 4050
rect -3230 4030 -3210 4050
rect -3190 4030 -3170 4050
rect -3150 4030 -3130 4050
rect -3110 4030 -3095 4050
rect -5595 4020 -3095 4030
rect -2045 4050 455 4060
rect -2045 4030 -2030 4050
rect -2010 4030 -1990 4050
rect -1970 4030 -1950 4050
rect -1930 4030 -1910 4050
rect -1890 4030 -1870 4050
rect -1850 4030 -1830 4050
rect -1810 4030 -1790 4050
rect -1770 4030 -1750 4050
rect -1730 4030 -1710 4050
rect -1690 4030 -1670 4050
rect -1650 4030 -1630 4050
rect -1610 4030 -1590 4050
rect -1570 4030 -1550 4050
rect -1530 4030 -1510 4050
rect -1490 4030 -1470 4050
rect -1450 4030 -1430 4050
rect -1410 4030 -1390 4050
rect -1370 4030 -1350 4050
rect -1330 4030 -1310 4050
rect -1290 4030 -1270 4050
rect -1250 4030 -1230 4050
rect -1210 4030 -1190 4050
rect -1170 4030 -1150 4050
rect -1130 4030 -1110 4050
rect -1090 4030 -1070 4050
rect -1050 4030 -1030 4050
rect -1010 4030 -990 4050
rect -970 4030 -950 4050
rect -930 4030 -910 4050
rect -890 4030 -870 4050
rect -850 4030 -830 4050
rect -810 4030 -790 4050
rect -770 4030 -750 4050
rect -730 4030 -710 4050
rect -690 4030 -670 4050
rect -650 4030 -630 4050
rect -610 4030 -590 4050
rect -570 4030 -550 4050
rect -530 4030 -510 4050
rect -490 4030 -470 4050
rect -450 4030 -430 4050
rect -410 4030 -390 4050
rect -370 4030 -350 4050
rect -330 4030 -310 4050
rect -290 4030 -270 4050
rect -250 4030 -230 4050
rect -210 4030 -190 4050
rect -170 4030 -150 4050
rect -130 4030 -110 4050
rect -90 4030 -70 4050
rect -50 4030 -30 4050
rect -10 4030 10 4050
rect 30 4030 50 4050
rect 70 4030 90 4050
rect 110 4030 130 4050
rect 150 4030 170 4050
rect 190 4030 210 4050
rect 230 4030 250 4050
rect 270 4030 290 4050
rect 310 4030 330 4050
rect 350 4030 370 4050
rect 390 4030 410 4050
rect 440 4030 455 4050
rect -2045 4020 455 4030
rect -3075 4005 -2920 4015
rect -3050 3980 -3030 4005
rect -3010 3980 -2990 4005
rect -2970 3980 -2950 4005
rect -2930 3980 -2920 4005
rect -3075 3970 -2920 3980
rect -2220 4005 -2065 4015
rect -2220 3980 -2210 4005
rect -2190 3980 -2170 4005
rect -2150 3980 -2130 4005
rect -2110 3980 -2090 4005
rect -2220 3970 -2065 3980
rect -5595 3955 -3095 3965
rect -5595 3935 -5580 3955
rect -5550 3935 -5530 3955
rect -5510 3935 -5490 3955
rect -5470 3935 -5450 3955
rect -5430 3935 -5410 3955
rect -5390 3935 -5370 3955
rect -5350 3935 -5330 3955
rect -5310 3935 -5290 3955
rect -5270 3935 -5250 3955
rect -5230 3935 -5210 3955
rect -5190 3935 -5170 3955
rect -5150 3935 -5130 3955
rect -5110 3935 -5090 3955
rect -5070 3935 -5050 3955
rect -5030 3935 -5010 3955
rect -4990 3935 -4970 3955
rect -4950 3935 -4930 3955
rect -4910 3935 -4890 3955
rect -4870 3935 -4850 3955
rect -4830 3935 -4810 3955
rect -4790 3935 -4770 3955
rect -4750 3935 -4730 3955
rect -4710 3935 -4690 3955
rect -4670 3935 -4650 3955
rect -4630 3935 -4610 3955
rect -4590 3935 -4570 3955
rect -4550 3935 -4530 3955
rect -4510 3935 -4490 3955
rect -4470 3935 -4450 3955
rect -4430 3935 -4410 3955
rect -4390 3935 -4370 3955
rect -4350 3935 -4330 3955
rect -4310 3935 -4290 3955
rect -4270 3935 -4250 3955
rect -4230 3935 -4210 3955
rect -4190 3935 -4170 3955
rect -4150 3935 -4130 3955
rect -4110 3935 -4090 3955
rect -4070 3935 -4050 3955
rect -4030 3935 -4010 3955
rect -3990 3935 -3970 3955
rect -3950 3935 -3930 3955
rect -3910 3935 -3890 3955
rect -3870 3935 -3850 3955
rect -3830 3935 -3810 3955
rect -3790 3935 -3770 3955
rect -3750 3935 -3730 3955
rect -3710 3935 -3690 3955
rect -3670 3935 -3650 3955
rect -3630 3935 -3610 3955
rect -3590 3935 -3570 3955
rect -3550 3935 -3530 3955
rect -3510 3935 -3490 3955
rect -3470 3935 -3450 3955
rect -3430 3935 -3410 3955
rect -3390 3935 -3370 3955
rect -3350 3935 -3330 3955
rect -3310 3935 -3290 3955
rect -3270 3935 -3250 3955
rect -3230 3935 -3210 3955
rect -3190 3935 -3170 3955
rect -3150 3935 -3130 3955
rect -3110 3935 -3095 3955
rect -5595 3925 -3095 3935
rect -2045 3955 455 3965
rect -2045 3935 -2030 3955
rect -2010 3935 -1990 3955
rect -1970 3935 -1950 3955
rect -1930 3935 -1910 3955
rect -1890 3935 -1870 3955
rect -1850 3935 -1830 3955
rect -1810 3935 -1790 3955
rect -1770 3935 -1750 3955
rect -1730 3935 -1710 3955
rect -1690 3935 -1670 3955
rect -1650 3935 -1630 3955
rect -1610 3935 -1590 3955
rect -1570 3935 -1550 3955
rect -1530 3935 -1510 3955
rect -1490 3935 -1470 3955
rect -1450 3935 -1430 3955
rect -1410 3935 -1390 3955
rect -1370 3935 -1350 3955
rect -1330 3935 -1310 3955
rect -1290 3935 -1270 3955
rect -1250 3935 -1230 3955
rect -1210 3935 -1190 3955
rect -1170 3935 -1150 3955
rect -1130 3935 -1110 3955
rect -1090 3935 -1070 3955
rect -1050 3935 -1030 3955
rect -1010 3935 -990 3955
rect -970 3935 -950 3955
rect -930 3935 -910 3955
rect -890 3935 -870 3955
rect -850 3935 -830 3955
rect -810 3935 -790 3955
rect -770 3935 -750 3955
rect -730 3935 -710 3955
rect -690 3935 -670 3955
rect -650 3935 -630 3955
rect -610 3935 -590 3955
rect -570 3935 -550 3955
rect -530 3935 -510 3955
rect -490 3935 -470 3955
rect -450 3935 -430 3955
rect -410 3935 -390 3955
rect -370 3935 -350 3955
rect -330 3935 -310 3955
rect -290 3935 -270 3955
rect -250 3935 -230 3955
rect -210 3935 -190 3955
rect -170 3935 -150 3955
rect -130 3935 -110 3955
rect -90 3935 -70 3955
rect -50 3935 -30 3955
rect -10 3935 10 3955
rect 30 3935 50 3955
rect 70 3935 90 3955
rect 110 3935 130 3955
rect 150 3935 170 3955
rect 190 3935 210 3955
rect 230 3935 250 3955
rect 270 3935 290 3955
rect 310 3935 330 3955
rect 350 3935 370 3955
rect 390 3935 410 3955
rect 440 3935 455 3955
rect -2045 3925 455 3935
rect -3075 3910 -2920 3920
rect -3050 3885 -3030 3910
rect -3010 3885 -2990 3910
rect -2970 3885 -2950 3910
rect -2930 3885 -2920 3910
rect -3075 3875 -2920 3885
rect -2220 3910 -2065 3920
rect -2220 3885 -2210 3910
rect -2190 3885 -2170 3910
rect -2150 3885 -2130 3910
rect -2110 3885 -2090 3910
rect -2220 3875 -2065 3885
rect -5595 3860 -3095 3870
rect -5595 3840 -5580 3860
rect -5550 3840 -5530 3860
rect -5510 3840 -5490 3860
rect -5470 3840 -5450 3860
rect -5430 3840 -5410 3860
rect -5390 3840 -5370 3860
rect -5350 3840 -5330 3860
rect -5310 3840 -5290 3860
rect -5270 3840 -5250 3860
rect -5230 3840 -5210 3860
rect -5190 3840 -5170 3860
rect -5150 3840 -5130 3860
rect -5110 3840 -5090 3860
rect -5070 3840 -5050 3860
rect -5030 3840 -5010 3860
rect -4990 3840 -4970 3860
rect -4950 3840 -4930 3860
rect -4910 3840 -4890 3860
rect -4870 3840 -4850 3860
rect -4830 3840 -4810 3860
rect -4790 3840 -4770 3860
rect -4750 3840 -4730 3860
rect -4710 3840 -4690 3860
rect -4670 3840 -4650 3860
rect -4630 3840 -4610 3860
rect -4590 3840 -4570 3860
rect -4550 3840 -4530 3860
rect -4510 3840 -4490 3860
rect -4470 3840 -4450 3860
rect -4430 3840 -4410 3860
rect -4390 3840 -4370 3860
rect -4350 3840 -4330 3860
rect -4310 3840 -4290 3860
rect -4270 3840 -4250 3860
rect -4230 3840 -4210 3860
rect -4190 3840 -4170 3860
rect -4150 3840 -4130 3860
rect -4110 3840 -4090 3860
rect -4070 3840 -4050 3860
rect -4030 3840 -4010 3860
rect -3990 3840 -3970 3860
rect -3950 3840 -3930 3860
rect -3910 3840 -3890 3860
rect -3870 3840 -3850 3860
rect -3830 3840 -3810 3860
rect -3790 3840 -3770 3860
rect -3750 3840 -3730 3860
rect -3710 3840 -3690 3860
rect -3670 3840 -3650 3860
rect -3630 3840 -3610 3860
rect -3590 3840 -3570 3860
rect -3550 3840 -3530 3860
rect -3510 3840 -3490 3860
rect -3470 3840 -3450 3860
rect -3430 3840 -3410 3860
rect -3390 3840 -3370 3860
rect -3350 3840 -3330 3860
rect -3310 3840 -3290 3860
rect -3270 3840 -3250 3860
rect -3230 3840 -3210 3860
rect -3190 3840 -3170 3860
rect -3150 3840 -3130 3860
rect -3110 3840 -3095 3860
rect -5595 3830 -3095 3840
rect -2045 3860 455 3870
rect -2045 3840 -2030 3860
rect -2010 3840 -1990 3860
rect -1970 3840 -1950 3860
rect -1930 3840 -1910 3860
rect -1890 3840 -1870 3860
rect -1850 3840 -1830 3860
rect -1810 3840 -1790 3860
rect -1770 3840 -1750 3860
rect -1730 3840 -1710 3860
rect -1690 3840 -1670 3860
rect -1650 3840 -1630 3860
rect -1610 3840 -1590 3860
rect -1570 3840 -1550 3860
rect -1530 3840 -1510 3860
rect -1490 3840 -1470 3860
rect -1450 3840 -1430 3860
rect -1410 3840 -1390 3860
rect -1370 3840 -1350 3860
rect -1330 3840 -1310 3860
rect -1290 3840 -1270 3860
rect -1250 3840 -1230 3860
rect -1210 3840 -1190 3860
rect -1170 3840 -1150 3860
rect -1130 3840 -1110 3860
rect -1090 3840 -1070 3860
rect -1050 3840 -1030 3860
rect -1010 3840 -990 3860
rect -970 3840 -950 3860
rect -930 3840 -910 3860
rect -890 3840 -870 3860
rect -850 3840 -830 3860
rect -810 3840 -790 3860
rect -770 3840 -750 3860
rect -730 3840 -710 3860
rect -690 3840 -670 3860
rect -650 3840 -630 3860
rect -610 3840 -590 3860
rect -570 3840 -550 3860
rect -530 3840 -510 3860
rect -490 3840 -470 3860
rect -450 3840 -430 3860
rect -410 3840 -390 3860
rect -370 3840 -350 3860
rect -330 3840 -310 3860
rect -290 3840 -270 3860
rect -250 3840 -230 3860
rect -210 3840 -190 3860
rect -170 3840 -150 3860
rect -130 3840 -110 3860
rect -90 3840 -70 3860
rect -50 3840 -30 3860
rect -10 3840 10 3860
rect 30 3840 50 3860
rect 70 3840 90 3860
rect 110 3840 130 3860
rect 150 3840 170 3860
rect 190 3840 210 3860
rect 230 3840 250 3860
rect 270 3840 290 3860
rect 310 3840 330 3860
rect 350 3840 370 3860
rect 390 3840 410 3860
rect 440 3840 455 3860
rect -2045 3830 455 3840
rect -3075 3815 -2920 3825
rect -3050 3790 -3030 3815
rect -3010 3790 -2990 3815
rect -2970 3790 -2950 3815
rect -2930 3790 -2920 3815
rect -3075 3780 -2920 3790
rect -2220 3815 -2065 3825
rect -2220 3790 -2210 3815
rect -2190 3790 -2170 3815
rect -2150 3790 -2130 3815
rect -2110 3790 -2090 3815
rect -2220 3780 -2065 3790
rect -5595 3765 -3095 3775
rect -5595 3745 -5580 3765
rect -5550 3745 -5530 3765
rect -5510 3745 -5490 3765
rect -5470 3745 -5450 3765
rect -5430 3745 -5410 3765
rect -5390 3745 -5370 3765
rect -5350 3745 -5330 3765
rect -5310 3745 -5290 3765
rect -5270 3745 -5250 3765
rect -5230 3745 -5210 3765
rect -5190 3745 -5170 3765
rect -5150 3745 -5130 3765
rect -5110 3745 -5090 3765
rect -5070 3745 -5050 3765
rect -5030 3745 -5010 3765
rect -4990 3745 -4970 3765
rect -4950 3745 -4930 3765
rect -4910 3745 -4890 3765
rect -4870 3745 -4850 3765
rect -4830 3745 -4810 3765
rect -4790 3745 -4770 3765
rect -4750 3745 -4730 3765
rect -4710 3745 -4690 3765
rect -4670 3745 -4650 3765
rect -4630 3745 -4610 3765
rect -4590 3745 -4570 3765
rect -4550 3745 -4530 3765
rect -4510 3745 -4490 3765
rect -4470 3745 -4450 3765
rect -4430 3745 -4410 3765
rect -4390 3745 -4370 3765
rect -4350 3745 -4330 3765
rect -4310 3745 -4290 3765
rect -4270 3745 -4250 3765
rect -4230 3745 -4210 3765
rect -4190 3745 -4170 3765
rect -4150 3745 -4130 3765
rect -4110 3745 -4090 3765
rect -4070 3745 -4050 3765
rect -4030 3745 -4010 3765
rect -3990 3745 -3970 3765
rect -3950 3745 -3930 3765
rect -3910 3745 -3890 3765
rect -3870 3745 -3850 3765
rect -3830 3745 -3810 3765
rect -3790 3745 -3770 3765
rect -3750 3745 -3730 3765
rect -3710 3745 -3690 3765
rect -3670 3745 -3650 3765
rect -3630 3745 -3610 3765
rect -3590 3745 -3570 3765
rect -3550 3745 -3530 3765
rect -3510 3745 -3490 3765
rect -3470 3745 -3450 3765
rect -3430 3745 -3410 3765
rect -3390 3745 -3370 3765
rect -3350 3745 -3330 3765
rect -3310 3745 -3290 3765
rect -3270 3745 -3250 3765
rect -3230 3745 -3210 3765
rect -3190 3745 -3170 3765
rect -3150 3745 -3130 3765
rect -3110 3745 -3095 3765
rect -5595 3735 -3095 3745
rect -2045 3765 455 3775
rect -2045 3745 -2030 3765
rect -2010 3745 -1990 3765
rect -1970 3745 -1950 3765
rect -1930 3745 -1910 3765
rect -1890 3745 -1870 3765
rect -1850 3745 -1830 3765
rect -1810 3745 -1790 3765
rect -1770 3745 -1750 3765
rect -1730 3745 -1710 3765
rect -1690 3745 -1670 3765
rect -1650 3745 -1630 3765
rect -1610 3745 -1590 3765
rect -1570 3745 -1550 3765
rect -1530 3745 -1510 3765
rect -1490 3745 -1470 3765
rect -1450 3745 -1430 3765
rect -1410 3745 -1390 3765
rect -1370 3745 -1350 3765
rect -1330 3745 -1310 3765
rect -1290 3745 -1270 3765
rect -1250 3745 -1230 3765
rect -1210 3745 -1190 3765
rect -1170 3745 -1150 3765
rect -1130 3745 -1110 3765
rect -1090 3745 -1070 3765
rect -1050 3745 -1030 3765
rect -1010 3745 -990 3765
rect -970 3745 -950 3765
rect -930 3745 -910 3765
rect -890 3745 -870 3765
rect -850 3745 -830 3765
rect -810 3745 -790 3765
rect -770 3745 -750 3765
rect -730 3745 -710 3765
rect -690 3745 -670 3765
rect -650 3745 -630 3765
rect -610 3745 -590 3765
rect -570 3745 -550 3765
rect -530 3745 -510 3765
rect -490 3745 -470 3765
rect -450 3745 -430 3765
rect -410 3745 -390 3765
rect -370 3745 -350 3765
rect -330 3745 -310 3765
rect -290 3745 -270 3765
rect -250 3745 -230 3765
rect -210 3745 -190 3765
rect -170 3745 -150 3765
rect -130 3745 -110 3765
rect -90 3745 -70 3765
rect -50 3745 -30 3765
rect -10 3745 10 3765
rect 30 3745 50 3765
rect 70 3745 90 3765
rect 110 3745 130 3765
rect 150 3745 170 3765
rect 190 3745 210 3765
rect 230 3745 250 3765
rect 270 3745 290 3765
rect 310 3745 330 3765
rect 350 3745 370 3765
rect 390 3745 410 3765
rect 440 3745 455 3765
rect -2045 3735 455 3745
rect -3075 3720 -2920 3730
rect -3050 3695 -3030 3720
rect -3010 3695 -2990 3720
rect -2970 3695 -2950 3720
rect -2930 3695 -2920 3720
rect -3075 3685 -2920 3695
rect -2220 3720 -2065 3730
rect -2220 3695 -2210 3720
rect -2190 3695 -2170 3720
rect -2150 3695 -2130 3720
rect -2110 3695 -2090 3720
rect -2220 3685 -2065 3695
rect -5595 3670 -3095 3680
rect -5595 3650 -5580 3670
rect -5550 3650 -5530 3670
rect -5510 3650 -5490 3670
rect -5470 3650 -5450 3670
rect -5430 3650 -5410 3670
rect -5390 3650 -5370 3670
rect -5350 3650 -5330 3670
rect -5310 3650 -5290 3670
rect -5270 3650 -5250 3670
rect -5230 3650 -5210 3670
rect -5190 3650 -5170 3670
rect -5150 3650 -5130 3670
rect -5110 3650 -5090 3670
rect -5070 3650 -5050 3670
rect -5030 3650 -5010 3670
rect -4990 3650 -4970 3670
rect -4950 3650 -4930 3670
rect -4910 3650 -4890 3670
rect -4870 3650 -4850 3670
rect -4830 3650 -4810 3670
rect -4790 3650 -4770 3670
rect -4750 3650 -4730 3670
rect -4710 3650 -4690 3670
rect -4670 3650 -4650 3670
rect -4630 3650 -4610 3670
rect -4590 3650 -4570 3670
rect -4550 3650 -4530 3670
rect -4510 3650 -4490 3670
rect -4470 3650 -4450 3670
rect -4430 3650 -4410 3670
rect -4390 3650 -4370 3670
rect -4350 3650 -4330 3670
rect -4310 3650 -4290 3670
rect -4270 3650 -4250 3670
rect -4230 3650 -4210 3670
rect -4190 3650 -4170 3670
rect -4150 3650 -4130 3670
rect -4110 3650 -4090 3670
rect -4070 3650 -4050 3670
rect -4030 3650 -4010 3670
rect -3990 3650 -3970 3670
rect -3950 3650 -3930 3670
rect -3910 3650 -3890 3670
rect -3870 3650 -3850 3670
rect -3830 3650 -3810 3670
rect -3790 3650 -3770 3670
rect -3750 3650 -3730 3670
rect -3710 3650 -3690 3670
rect -3670 3650 -3650 3670
rect -3630 3650 -3610 3670
rect -3590 3650 -3570 3670
rect -3550 3650 -3530 3670
rect -3510 3650 -3490 3670
rect -3470 3650 -3450 3670
rect -3430 3650 -3410 3670
rect -3390 3650 -3370 3670
rect -3350 3650 -3330 3670
rect -3310 3650 -3290 3670
rect -3270 3650 -3250 3670
rect -3230 3650 -3210 3670
rect -3190 3650 -3170 3670
rect -3150 3650 -3130 3670
rect -3110 3650 -3095 3670
rect -5595 3640 -3095 3650
rect -2045 3670 455 3680
rect -2045 3650 -2030 3670
rect -2010 3650 -1990 3670
rect -1970 3650 -1950 3670
rect -1930 3650 -1910 3670
rect -1890 3650 -1870 3670
rect -1850 3650 -1830 3670
rect -1810 3650 -1790 3670
rect -1770 3650 -1750 3670
rect -1730 3650 -1710 3670
rect -1690 3650 -1670 3670
rect -1650 3650 -1630 3670
rect -1610 3650 -1590 3670
rect -1570 3650 -1550 3670
rect -1530 3650 -1510 3670
rect -1490 3650 -1470 3670
rect -1450 3650 -1430 3670
rect -1410 3650 -1390 3670
rect -1370 3650 -1350 3670
rect -1330 3650 -1310 3670
rect -1290 3650 -1270 3670
rect -1250 3650 -1230 3670
rect -1210 3650 -1190 3670
rect -1170 3650 -1150 3670
rect -1130 3650 -1110 3670
rect -1090 3650 -1070 3670
rect -1050 3650 -1030 3670
rect -1010 3650 -990 3670
rect -970 3650 -950 3670
rect -930 3650 -910 3670
rect -890 3650 -870 3670
rect -850 3650 -830 3670
rect -810 3650 -790 3670
rect -770 3650 -750 3670
rect -730 3650 -710 3670
rect -690 3650 -670 3670
rect -650 3650 -630 3670
rect -610 3650 -590 3670
rect -570 3650 -550 3670
rect -530 3650 -510 3670
rect -490 3650 -470 3670
rect -450 3650 -430 3670
rect -410 3650 -390 3670
rect -370 3650 -350 3670
rect -330 3650 -310 3670
rect -290 3650 -270 3670
rect -250 3650 -230 3670
rect -210 3650 -190 3670
rect -170 3650 -150 3670
rect -130 3650 -110 3670
rect -90 3650 -70 3670
rect -50 3650 -30 3670
rect -10 3650 10 3670
rect 30 3650 50 3670
rect 70 3650 90 3670
rect 110 3650 130 3670
rect 150 3650 170 3670
rect 190 3650 210 3670
rect 230 3650 250 3670
rect 270 3650 290 3670
rect 310 3650 330 3670
rect 350 3650 370 3670
rect 390 3650 410 3670
rect 440 3650 455 3670
rect -2045 3640 455 3650
rect -3075 3625 -2920 3635
rect -3050 3600 -3030 3625
rect -3010 3600 -2990 3625
rect -2970 3600 -2950 3625
rect -2930 3600 -2920 3625
rect -3075 3590 -2920 3600
rect -2220 3625 -2065 3635
rect -2220 3600 -2210 3625
rect -2190 3600 -2170 3625
rect -2150 3600 -2130 3625
rect -2110 3600 -2090 3625
rect -2220 3590 -2065 3600
rect -5595 3575 -3095 3585
rect -5595 3555 -5580 3575
rect -5550 3555 -5530 3575
rect -5510 3555 -5490 3575
rect -5470 3555 -5450 3575
rect -5430 3555 -5410 3575
rect -5390 3555 -5370 3575
rect -5350 3555 -5330 3575
rect -5310 3555 -5290 3575
rect -5270 3555 -5250 3575
rect -5230 3555 -5210 3575
rect -5190 3555 -5170 3575
rect -5150 3555 -5130 3575
rect -5110 3555 -5090 3575
rect -5070 3555 -5050 3575
rect -5030 3555 -5010 3575
rect -4990 3555 -4970 3575
rect -4950 3555 -4930 3575
rect -4910 3555 -4890 3575
rect -4870 3555 -4850 3575
rect -4830 3555 -4810 3575
rect -4790 3555 -4770 3575
rect -4750 3555 -4730 3575
rect -4710 3555 -4690 3575
rect -4670 3555 -4650 3575
rect -4630 3555 -4610 3575
rect -4590 3555 -4570 3575
rect -4550 3555 -4530 3575
rect -4510 3555 -4490 3575
rect -4470 3555 -4450 3575
rect -4430 3555 -4410 3575
rect -4390 3555 -4370 3575
rect -4350 3555 -4330 3575
rect -4310 3555 -4290 3575
rect -4270 3555 -4250 3575
rect -4230 3555 -4210 3575
rect -4190 3555 -4170 3575
rect -4150 3555 -4130 3575
rect -4110 3555 -4090 3575
rect -4070 3555 -4050 3575
rect -4030 3555 -4010 3575
rect -3990 3555 -3970 3575
rect -3950 3555 -3930 3575
rect -3910 3555 -3890 3575
rect -3870 3555 -3850 3575
rect -3830 3555 -3810 3575
rect -3790 3555 -3770 3575
rect -3750 3555 -3730 3575
rect -3710 3555 -3690 3575
rect -3670 3555 -3650 3575
rect -3630 3555 -3610 3575
rect -3590 3555 -3570 3575
rect -3550 3555 -3530 3575
rect -3510 3555 -3490 3575
rect -3470 3555 -3450 3575
rect -3430 3555 -3410 3575
rect -3390 3555 -3370 3575
rect -3350 3555 -3330 3575
rect -3310 3555 -3290 3575
rect -3270 3555 -3250 3575
rect -3230 3555 -3210 3575
rect -3190 3555 -3170 3575
rect -3150 3555 -3130 3575
rect -3110 3555 -3095 3575
rect -5595 3535 -3095 3555
rect -5595 3515 -5580 3535
rect -5550 3515 -5530 3535
rect -5510 3515 -5490 3535
rect -5470 3515 -5450 3535
rect -5430 3515 -5410 3535
rect -5390 3515 -5370 3535
rect -5350 3515 -5330 3535
rect -5310 3515 -5290 3535
rect -5270 3515 -5250 3535
rect -5230 3515 -5210 3535
rect -5190 3515 -5170 3535
rect -5150 3515 -5130 3535
rect -5110 3515 -5090 3535
rect -5070 3515 -5050 3535
rect -5030 3515 -5010 3535
rect -4990 3515 -4970 3535
rect -4950 3515 -4930 3535
rect -4910 3515 -4890 3535
rect -4870 3515 -4850 3535
rect -4830 3515 -4810 3535
rect -4790 3515 -4770 3535
rect -4750 3515 -4730 3535
rect -4710 3515 -4690 3535
rect -4670 3515 -4650 3535
rect -4630 3515 -4610 3535
rect -4590 3515 -4570 3535
rect -4550 3515 -4530 3535
rect -4510 3515 -4490 3535
rect -4470 3515 -4450 3535
rect -4430 3515 -4410 3535
rect -4390 3515 -4370 3535
rect -4350 3515 -4330 3535
rect -4310 3515 -4290 3535
rect -4270 3515 -4250 3535
rect -4230 3515 -4210 3535
rect -4190 3515 -4170 3535
rect -4150 3515 -4130 3535
rect -4110 3515 -4090 3535
rect -4070 3515 -4050 3535
rect -4030 3515 -4010 3535
rect -3990 3515 -3970 3535
rect -3950 3515 -3930 3535
rect -3910 3515 -3890 3535
rect -3870 3515 -3850 3535
rect -3830 3515 -3810 3535
rect -3790 3515 -3770 3535
rect -3750 3515 -3730 3535
rect -3710 3515 -3690 3535
rect -3670 3515 -3650 3535
rect -3630 3515 -3610 3535
rect -3590 3515 -3570 3535
rect -3550 3515 -3530 3535
rect -3510 3515 -3490 3535
rect -3470 3515 -3450 3535
rect -3430 3515 -3410 3535
rect -3390 3515 -3370 3535
rect -3350 3515 -3330 3535
rect -3310 3515 -3290 3535
rect -3270 3515 -3250 3535
rect -3230 3515 -3210 3535
rect -3190 3515 -3170 3535
rect -3150 3515 -3130 3535
rect -3110 3515 -3095 3535
rect -5595 3505 -3095 3515
rect -2045 3575 455 3585
rect -2045 3555 -2030 3575
rect -2010 3555 -1990 3575
rect -1970 3555 -1950 3575
rect -1930 3555 -1910 3575
rect -1890 3555 -1870 3575
rect -1850 3555 -1830 3575
rect -1810 3555 -1790 3575
rect -1770 3555 -1750 3575
rect -1730 3555 -1710 3575
rect -1690 3555 -1670 3575
rect -1650 3555 -1630 3575
rect -1610 3555 -1590 3575
rect -1570 3555 -1550 3575
rect -1530 3555 -1510 3575
rect -1490 3555 -1470 3575
rect -1450 3555 -1430 3575
rect -1410 3555 -1390 3575
rect -1370 3555 -1350 3575
rect -1330 3555 -1310 3575
rect -1290 3555 -1270 3575
rect -1250 3555 -1230 3575
rect -1210 3555 -1190 3575
rect -1170 3555 -1150 3575
rect -1130 3555 -1110 3575
rect -1090 3555 -1070 3575
rect -1050 3555 -1030 3575
rect -1010 3555 -990 3575
rect -970 3555 -950 3575
rect -930 3555 -910 3575
rect -890 3555 -870 3575
rect -850 3555 -830 3575
rect -810 3555 -790 3575
rect -770 3555 -750 3575
rect -730 3555 -710 3575
rect -690 3555 -670 3575
rect -650 3555 -630 3575
rect -610 3555 -590 3575
rect -570 3555 -550 3575
rect -530 3555 -510 3575
rect -490 3555 -470 3575
rect -450 3555 -430 3575
rect -410 3555 -390 3575
rect -370 3555 -350 3575
rect -330 3555 -310 3575
rect -290 3555 -270 3575
rect -250 3555 -230 3575
rect -210 3555 -190 3575
rect -170 3555 -150 3575
rect -130 3555 -110 3575
rect -90 3555 -70 3575
rect -50 3555 -30 3575
rect -10 3555 10 3575
rect 30 3555 50 3575
rect 70 3555 90 3575
rect 110 3555 130 3575
rect 150 3555 170 3575
rect 190 3555 210 3575
rect 230 3555 250 3575
rect 270 3555 290 3575
rect 310 3555 330 3575
rect 350 3555 370 3575
rect 390 3555 410 3575
rect 440 3555 455 3575
rect -2045 3535 455 3555
rect -2045 3515 -2030 3535
rect -2010 3515 -1990 3535
rect -1970 3515 -1950 3535
rect -1930 3515 -1910 3535
rect -1890 3515 -1870 3535
rect -1850 3515 -1830 3535
rect -1810 3515 -1790 3535
rect -1770 3515 -1750 3535
rect -1730 3515 -1710 3535
rect -1690 3515 -1670 3535
rect -1650 3515 -1630 3535
rect -1610 3515 -1590 3535
rect -1570 3515 -1550 3535
rect -1530 3515 -1510 3535
rect -1490 3515 -1470 3535
rect -1450 3515 -1430 3535
rect -1410 3515 -1390 3535
rect -1370 3515 -1350 3535
rect -1330 3515 -1310 3535
rect -1290 3515 -1270 3535
rect -1250 3515 -1230 3535
rect -1210 3515 -1190 3535
rect -1170 3515 -1150 3535
rect -1130 3515 -1110 3535
rect -1090 3515 -1070 3535
rect -1050 3515 -1030 3535
rect -1010 3515 -990 3535
rect -970 3515 -950 3535
rect -930 3515 -910 3535
rect -890 3515 -870 3535
rect -850 3515 -830 3535
rect -810 3515 -790 3535
rect -770 3515 -750 3535
rect -730 3515 -710 3535
rect -690 3515 -670 3535
rect -650 3515 -630 3535
rect -610 3515 -590 3535
rect -570 3515 -550 3535
rect -530 3515 -510 3535
rect -490 3515 -470 3535
rect -450 3515 -430 3535
rect -410 3515 -390 3535
rect -370 3515 -350 3535
rect -330 3515 -310 3535
rect -290 3515 -270 3535
rect -250 3515 -230 3535
rect -210 3515 -190 3535
rect -170 3515 -150 3535
rect -130 3515 -110 3535
rect -90 3515 -70 3535
rect -50 3515 -30 3535
rect -10 3515 10 3535
rect 30 3515 50 3535
rect 70 3515 90 3535
rect 110 3515 130 3535
rect 150 3515 170 3535
rect 190 3515 210 3535
rect 230 3515 250 3535
rect 270 3515 290 3535
rect 310 3515 330 3535
rect 350 3515 370 3535
rect 390 3515 410 3535
rect 440 3515 455 3535
rect -2045 3505 455 3515
<< viali >>
rect -5510 8585 -5490 8605
rect -5470 8585 -5450 8605
rect -5430 8585 -5410 8605
rect -5390 8585 -5370 8605
rect -5350 8585 -5330 8605
rect -5310 8585 -5290 8605
rect -5270 8585 -5250 8605
rect -5230 8585 -5210 8605
rect -5190 8585 -5170 8605
rect -5150 8585 -5130 8605
rect -5110 8585 -5090 8605
rect -5070 8585 -5050 8605
rect -5030 8585 -5010 8605
rect -4990 8585 -4970 8605
rect -4950 8585 -4930 8605
rect -4910 8585 -4890 8605
rect -4870 8585 -4850 8605
rect -4830 8585 -4810 8605
rect -4790 8585 -4770 8605
rect -4450 8500 -4430 8520
rect -4410 8500 -4390 8520
rect -4370 8500 -4350 8520
rect -4330 8500 -4310 8520
rect -4290 8500 -4270 8520
rect -4250 8500 -4230 8520
rect -4210 8500 -4190 8520
rect -4170 8500 -4150 8520
rect -4130 8500 -4110 8520
rect -4090 8500 -4070 8520
rect -4050 8500 -4030 8520
rect -4010 8500 -3990 8520
rect -3970 8500 -3950 8520
rect -3930 8500 -3910 8520
rect -3890 8500 -3870 8520
rect -3850 8500 -3830 8520
rect -3810 8500 -3790 8520
rect -3770 8500 -3750 8520
rect -3730 8500 -3710 8520
rect -3690 8500 -3670 8520
rect -4450 8457 -4430 8477
rect -4410 8457 -4390 8477
rect -4370 8457 -4350 8477
rect -4330 8457 -4310 8477
rect -4290 8457 -4270 8477
rect -4250 8457 -4230 8477
rect -4210 8457 -4190 8477
rect -4170 8457 -4150 8477
rect -4130 8457 -4110 8477
rect -4090 8457 -4070 8477
rect -4050 8457 -4030 8477
rect -4010 8457 -3990 8477
rect -3970 8457 -3950 8477
rect -3930 8457 -3910 8477
rect -3890 8457 -3870 8477
rect -3850 8457 -3830 8477
rect -3810 8457 -3790 8477
rect -3770 8457 -3750 8477
rect -3730 8457 -3710 8477
rect -3690 8457 -3670 8477
rect -3140 8415 -3120 8435
rect -3100 8415 -3080 8435
rect -3060 8415 -3040 8435
rect -3020 8415 -3000 8435
rect -5530 8375 -5510 8395
rect -5490 8375 -5470 8395
rect -5450 8375 -5430 8395
rect -5410 8375 -5390 8395
rect -5370 8375 -5350 8395
rect -5330 8375 -5310 8395
rect -5290 8375 -5270 8395
rect -5250 8375 -5230 8395
rect -5210 8375 -5190 8395
rect -5170 8375 -5150 8395
rect -5130 8375 -5110 8395
rect -5090 8375 -5070 8395
rect -5050 8375 -5030 8395
rect -5010 8375 -4990 8395
rect -4970 8375 -4950 8395
rect -4930 8375 -4910 8395
rect -4890 8375 -4870 8395
rect -4850 8375 -4830 8395
rect -4810 8375 -4790 8395
rect -4770 8375 -4750 8395
rect -3140 8335 -3120 8355
rect -3100 8335 -3080 8355
rect -3060 8335 -3040 8355
rect -3020 8335 -3000 8355
rect -4450 8293 -4430 8313
rect -4410 8293 -4390 8313
rect -4370 8293 -4350 8313
rect -4330 8293 -4310 8313
rect -4290 8293 -4270 8313
rect -4250 8293 -4230 8313
rect -4210 8293 -4190 8313
rect -4170 8293 -4150 8313
rect -4130 8293 -4110 8313
rect -4090 8293 -4070 8313
rect -4050 8293 -4030 8313
rect -4010 8293 -3990 8313
rect -3970 8293 -3950 8313
rect -3930 8293 -3910 8313
rect -3890 8293 -3870 8313
rect -3850 8293 -3830 8313
rect -3810 8293 -3790 8313
rect -3770 8293 -3750 8313
rect -3730 8293 -3710 8313
rect -3690 8293 -3670 8313
rect -3140 8250 -3120 8270
rect -3100 8250 -3080 8270
rect -3060 8250 -3040 8270
rect -3020 8250 -3000 8270
rect -5530 8211 -5510 8231
rect -5490 8211 -5470 8231
rect -5450 8211 -5430 8231
rect -5410 8211 -5390 8231
rect -5370 8211 -5350 8231
rect -5330 8211 -5310 8231
rect -5290 8211 -5270 8231
rect -5250 8211 -5230 8231
rect -5210 8211 -5190 8231
rect -5170 8211 -5150 8231
rect -5130 8211 -5110 8231
rect -5090 8211 -5070 8231
rect -5050 8211 -5030 8231
rect -5010 8211 -4990 8231
rect -4970 8211 -4950 8231
rect -4930 8211 -4910 8231
rect -4890 8211 -4870 8231
rect -4850 8211 -4830 8231
rect -4810 8211 -4790 8231
rect -4770 8211 -4750 8231
rect -3140 8170 -3120 8190
rect -3100 8170 -3080 8190
rect -3060 8170 -3040 8190
rect -3020 8170 -3000 8190
rect -4450 8129 -4430 8149
rect -4410 8129 -4390 8149
rect -4370 8129 -4350 8149
rect -4330 8129 -4310 8149
rect -4290 8129 -4270 8149
rect -4250 8129 -4230 8149
rect -4210 8129 -4190 8149
rect -4170 8129 -4150 8149
rect -4130 8129 -4110 8149
rect -4090 8129 -4070 8149
rect -4050 8129 -4030 8149
rect -4010 8129 -3990 8149
rect -3970 8129 -3950 8149
rect -3930 8129 -3910 8149
rect -3890 8129 -3870 8149
rect -3850 8129 -3830 8149
rect -3810 8129 -3790 8149
rect -3770 8129 -3750 8149
rect -3730 8129 -3710 8149
rect -3690 8129 -3670 8149
rect -3140 8090 -3120 8110
rect -3100 8090 -3080 8110
rect -3060 8090 -3040 8110
rect -3020 8090 -3000 8110
rect -5530 8047 -5510 8067
rect -5490 8047 -5470 8067
rect -5450 8047 -5430 8067
rect -5410 8047 -5390 8067
rect -5370 8047 -5350 8067
rect -5330 8047 -5310 8067
rect -5290 8047 -5270 8067
rect -5250 8047 -5230 8067
rect -5210 8047 -5190 8067
rect -5170 8047 -5150 8067
rect -5130 8047 -5110 8067
rect -5090 8047 -5070 8067
rect -5050 8047 -5030 8067
rect -5010 8047 -4990 8067
rect -4970 8047 -4950 8067
rect -4930 8047 -4910 8067
rect -4890 8047 -4870 8067
rect -4850 8047 -4830 8067
rect -4810 8047 -4790 8067
rect -4770 8047 -4750 8067
rect -3140 8005 -3120 8025
rect -3100 8005 -3080 8025
rect -3060 8005 -3040 8025
rect -3020 8005 -3000 8025
rect -4450 7965 -4430 7985
rect -4410 7965 -4390 7985
rect -4370 7965 -4350 7985
rect -4330 7965 -4310 7985
rect -4290 7965 -4270 7985
rect -4250 7965 -4230 7985
rect -4210 7965 -4190 7985
rect -4170 7965 -4150 7985
rect -4130 7965 -4110 7985
rect -4090 7965 -4070 7985
rect -4050 7965 -4030 7985
rect -4010 7965 -3990 7985
rect -3970 7965 -3950 7985
rect -3930 7965 -3910 7985
rect -3890 7965 -3870 7985
rect -3850 7965 -3830 7985
rect -3810 7965 -3790 7985
rect -3770 7965 -3750 7985
rect -3730 7965 -3710 7985
rect -3690 7965 -3670 7985
rect -3140 7925 -3120 7945
rect -3100 7925 -3080 7945
rect -3060 7925 -3040 7945
rect -3020 7925 -3000 7945
rect -5530 7883 -5510 7903
rect -5490 7883 -5470 7903
rect -5450 7883 -5430 7903
rect -5410 7883 -5390 7903
rect -5370 7883 -5350 7903
rect -5330 7883 -5310 7903
rect -5290 7883 -5270 7903
rect -5250 7883 -5230 7903
rect -5210 7883 -5190 7903
rect -5170 7883 -5150 7903
rect -5130 7883 -5110 7903
rect -5090 7883 -5070 7903
rect -5050 7883 -5030 7903
rect -5010 7883 -4990 7903
rect -4970 7883 -4950 7903
rect -4930 7883 -4910 7903
rect -4890 7883 -4870 7903
rect -4850 7883 -4830 7903
rect -4810 7883 -4790 7903
rect -4770 7883 -4750 7903
rect -3140 7840 -3120 7860
rect -3100 7840 -3080 7860
rect -3060 7840 -3040 7860
rect -3020 7840 -3000 7860
rect -4450 7801 -4430 7821
rect -4410 7801 -4390 7821
rect -4370 7801 -4350 7821
rect -4330 7801 -4310 7821
rect -4290 7801 -4270 7821
rect -4250 7801 -4230 7821
rect -4210 7801 -4190 7821
rect -4170 7801 -4150 7821
rect -4130 7801 -4110 7821
rect -4090 7801 -4070 7821
rect -4050 7801 -4030 7821
rect -4010 7801 -3990 7821
rect -3970 7801 -3950 7821
rect -3930 7801 -3910 7821
rect -3890 7801 -3870 7821
rect -3850 7801 -3830 7821
rect -3810 7801 -3790 7821
rect -3770 7801 -3750 7821
rect -3730 7801 -3710 7821
rect -3690 7801 -3670 7821
rect -3140 7760 -3120 7780
rect -3100 7760 -3080 7780
rect -3060 7760 -3040 7780
rect -3020 7760 -3000 7780
rect -5530 7719 -5510 7739
rect -5490 7719 -5470 7739
rect -5450 7719 -5430 7739
rect -5410 7719 -5390 7739
rect -5370 7719 -5350 7739
rect -5330 7719 -5310 7739
rect -5290 7719 -5270 7739
rect -5250 7719 -5230 7739
rect -5210 7719 -5190 7739
rect -5170 7719 -5150 7739
rect -5130 7719 -5110 7739
rect -5090 7719 -5070 7739
rect -5050 7719 -5030 7739
rect -5010 7719 -4990 7739
rect -4970 7719 -4950 7739
rect -4930 7719 -4910 7739
rect -4890 7719 -4870 7739
rect -4850 7719 -4830 7739
rect -4810 7719 -4790 7739
rect -4770 7719 -4750 7739
rect -3140 7680 -3120 7700
rect -3100 7680 -3080 7700
rect -3060 7680 -3040 7700
rect -3020 7680 -3000 7700
rect -4450 7637 -4430 7657
rect -4410 7637 -4390 7657
rect -4370 7637 -4350 7657
rect -4330 7637 -4310 7657
rect -4290 7637 -4270 7657
rect -4250 7637 -4230 7657
rect -4210 7637 -4190 7657
rect -4170 7637 -4150 7657
rect -4130 7637 -4110 7657
rect -4090 7637 -4070 7657
rect -4050 7637 -4030 7657
rect -4010 7637 -3990 7657
rect -3970 7637 -3950 7657
rect -3930 7637 -3910 7657
rect -3890 7637 -3870 7657
rect -3850 7637 -3830 7657
rect -3810 7637 -3790 7657
rect -3770 7637 -3750 7657
rect -3730 7637 -3710 7657
rect -3690 7637 -3670 7657
rect -3140 7595 -3120 7615
rect -3100 7595 -3080 7615
rect -3060 7595 -3040 7615
rect -3020 7595 -3000 7615
rect -5530 7555 -5510 7575
rect -5490 7555 -5470 7575
rect -5450 7555 -5430 7575
rect -5410 7555 -5390 7575
rect -5370 7555 -5350 7575
rect -5330 7555 -5310 7575
rect -5290 7555 -5270 7575
rect -5250 7555 -5230 7575
rect -5210 7555 -5190 7575
rect -5170 7555 -5150 7575
rect -5130 7555 -5110 7575
rect -5090 7555 -5070 7575
rect -5050 7555 -5030 7575
rect -5010 7555 -4990 7575
rect -4970 7555 -4950 7575
rect -4930 7555 -4910 7575
rect -4890 7555 -4870 7575
rect -4850 7555 -4830 7575
rect -4810 7555 -4790 7575
rect -4770 7555 -4750 7575
rect -3140 7515 -3120 7535
rect -3100 7515 -3080 7535
rect -3060 7515 -3040 7535
rect -3020 7515 -3000 7535
rect -4450 7473 -4430 7493
rect -4410 7473 -4390 7493
rect -4370 7473 -4350 7493
rect -4330 7473 -4310 7493
rect -4290 7473 -4270 7493
rect -4250 7473 -4230 7493
rect -4210 7473 -4190 7493
rect -4170 7473 -4150 7493
rect -4130 7473 -4110 7493
rect -4090 7473 -4070 7493
rect -4050 7473 -4030 7493
rect -4010 7473 -3990 7493
rect -3970 7473 -3950 7493
rect -3930 7473 -3910 7493
rect -3890 7473 -3870 7493
rect -3850 7473 -3830 7493
rect -3810 7473 -3790 7493
rect -3770 7473 -3750 7493
rect -3730 7473 -3710 7493
rect -3690 7473 -3670 7493
rect -3140 7430 -3120 7450
rect -3100 7430 -3080 7450
rect -3060 7430 -3040 7450
rect -3020 7430 -3000 7450
rect -5530 7391 -5510 7411
rect -5490 7391 -5470 7411
rect -5450 7391 -5430 7411
rect -5410 7391 -5390 7411
rect -5370 7391 -5350 7411
rect -5330 7391 -5310 7411
rect -5290 7391 -5270 7411
rect -5250 7391 -5230 7411
rect -5210 7391 -5190 7411
rect -5170 7391 -5150 7411
rect -5130 7391 -5110 7411
rect -5090 7391 -5070 7411
rect -5050 7391 -5030 7411
rect -5010 7391 -4990 7411
rect -4970 7391 -4950 7411
rect -4930 7391 -4910 7411
rect -4890 7391 -4870 7411
rect -4850 7391 -4830 7411
rect -4810 7391 -4790 7411
rect -4770 7391 -4750 7411
rect -3140 7350 -3120 7370
rect -3100 7350 -3080 7370
rect -3060 7350 -3040 7370
rect -3020 7350 -3000 7370
rect -4450 7309 -4430 7329
rect -4410 7309 -4390 7329
rect -4370 7309 -4350 7329
rect -4330 7309 -4310 7329
rect -4290 7309 -4270 7329
rect -4250 7309 -4230 7329
rect -4210 7309 -4190 7329
rect -4170 7309 -4150 7329
rect -4130 7309 -4110 7329
rect -4090 7309 -4070 7329
rect -4050 7309 -4030 7329
rect -4010 7309 -3990 7329
rect -3970 7309 -3950 7329
rect -3930 7309 -3910 7329
rect -3890 7309 -3870 7329
rect -3850 7309 -3830 7329
rect -3810 7309 -3790 7329
rect -3770 7309 -3750 7329
rect -3730 7309 -3710 7329
rect -3690 7309 -3670 7329
rect -3140 7270 -3120 7290
rect -3100 7270 -3080 7290
rect -3060 7270 -3040 7290
rect -3020 7270 -3000 7290
rect -5530 7227 -5510 7247
rect -5490 7227 -5470 7247
rect -5450 7227 -5430 7247
rect -5410 7227 -5390 7247
rect -5370 7227 -5350 7247
rect -5330 7227 -5310 7247
rect -5290 7227 -5270 7247
rect -5250 7227 -5230 7247
rect -5210 7227 -5190 7247
rect -5170 7227 -5150 7247
rect -5130 7227 -5110 7247
rect -5090 7227 -5070 7247
rect -5050 7227 -5030 7247
rect -5010 7227 -4990 7247
rect -4970 7227 -4950 7247
rect -4930 7227 -4910 7247
rect -4890 7227 -4870 7247
rect -4850 7227 -4830 7247
rect -4810 7227 -4790 7247
rect -4770 7227 -4750 7247
rect -3140 7185 -3120 7205
rect -3100 7185 -3080 7205
rect -3060 7185 -3040 7205
rect -3020 7185 -3000 7205
rect -4450 7145 -4430 7165
rect -4410 7145 -4390 7165
rect -4370 7145 -4350 7165
rect -4330 7145 -4310 7165
rect -4290 7145 -4270 7165
rect -4250 7145 -4230 7165
rect -4210 7145 -4190 7165
rect -4170 7145 -4150 7165
rect -4130 7145 -4110 7165
rect -4090 7145 -4070 7165
rect -4050 7145 -4030 7165
rect -4010 7145 -3990 7165
rect -3970 7145 -3950 7165
rect -3930 7145 -3910 7165
rect -3890 7145 -3870 7165
rect -3850 7145 -3830 7165
rect -3810 7145 -3790 7165
rect -3770 7145 -3750 7165
rect -3730 7145 -3710 7165
rect -3690 7145 -3670 7165
rect -3140 7105 -3120 7125
rect -3100 7105 -3080 7125
rect -3060 7105 -3040 7125
rect -3020 7105 -3000 7125
rect -5530 7063 -5510 7083
rect -5490 7063 -5470 7083
rect -5450 7063 -5430 7083
rect -5410 7063 -5390 7083
rect -5370 7063 -5350 7083
rect -5330 7063 -5310 7083
rect -5290 7063 -5270 7083
rect -5250 7063 -5230 7083
rect -5210 7063 -5190 7083
rect -5170 7063 -5150 7083
rect -5130 7063 -5110 7083
rect -5090 7063 -5070 7083
rect -5050 7063 -5030 7083
rect -5010 7063 -4990 7083
rect -4970 7063 -4950 7083
rect -4930 7063 -4910 7083
rect -4890 7063 -4870 7083
rect -4850 7063 -4830 7083
rect -4810 7063 -4790 7083
rect -4770 7063 -4750 7083
rect -3140 7020 -3120 7040
rect -3100 7020 -3080 7040
rect -3060 7020 -3040 7040
rect -3020 7020 -3000 7040
rect -4450 6981 -4430 7001
rect -4410 6981 -4390 7001
rect -4370 6981 -4350 7001
rect -4330 6981 -4310 7001
rect -4290 6981 -4270 7001
rect -4250 6981 -4230 7001
rect -4210 6981 -4190 7001
rect -4170 6981 -4150 7001
rect -4130 6981 -4110 7001
rect -4090 6981 -4070 7001
rect -4050 6981 -4030 7001
rect -4010 6981 -3990 7001
rect -3970 6981 -3950 7001
rect -3930 6981 -3910 7001
rect -3890 6981 -3870 7001
rect -3850 6981 -3830 7001
rect -3810 6981 -3790 7001
rect -3770 6981 -3750 7001
rect -3730 6981 -3710 7001
rect -3690 6981 -3670 7001
rect -3140 6940 -3120 6960
rect -3100 6940 -3080 6960
rect -3060 6940 -3040 6960
rect -3020 6940 -3000 6960
rect -5530 6899 -5510 6919
rect -5490 6899 -5470 6919
rect -5450 6899 -5430 6919
rect -5410 6899 -5390 6919
rect -5370 6899 -5350 6919
rect -5330 6899 -5310 6919
rect -5290 6899 -5270 6919
rect -5250 6899 -5230 6919
rect -5210 6899 -5190 6919
rect -5170 6899 -5150 6919
rect -5130 6899 -5110 6919
rect -5090 6899 -5070 6919
rect -5050 6899 -5030 6919
rect -5010 6899 -4990 6919
rect -4970 6899 -4950 6919
rect -4930 6899 -4910 6919
rect -4890 6899 -4870 6919
rect -4850 6899 -4830 6919
rect -4810 6899 -4790 6919
rect -4770 6899 -4750 6919
rect -3140 6860 -3120 6880
rect -3100 6860 -3080 6880
rect -3060 6860 -3040 6880
rect -3020 6860 -3000 6880
rect -4450 6817 -4430 6837
rect -4410 6817 -4390 6837
rect -4370 6817 -4350 6837
rect -4330 6817 -4310 6837
rect -4290 6817 -4270 6837
rect -4250 6817 -4230 6837
rect -4210 6817 -4190 6837
rect -4170 6817 -4150 6837
rect -4130 6817 -4110 6837
rect -4090 6817 -4070 6837
rect -4050 6817 -4030 6837
rect -4010 6817 -3990 6837
rect -3970 6817 -3950 6837
rect -3930 6817 -3910 6837
rect -3890 6817 -3870 6837
rect -3850 6817 -3830 6837
rect -3810 6817 -3790 6837
rect -3770 6817 -3750 6837
rect -3730 6817 -3710 6837
rect -3690 6817 -3670 6837
rect -3140 6775 -3120 6795
rect -3100 6775 -3080 6795
rect -3060 6775 -3040 6795
rect -3020 6775 -3000 6795
rect -5530 6735 -5510 6755
rect -5490 6735 -5470 6755
rect -5450 6735 -5430 6755
rect -5410 6735 -5390 6755
rect -5370 6735 -5350 6755
rect -5330 6735 -5310 6755
rect -5290 6735 -5270 6755
rect -5250 6735 -5230 6755
rect -5210 6735 -5190 6755
rect -5170 6735 -5150 6755
rect -5130 6735 -5110 6755
rect -5090 6735 -5070 6755
rect -5050 6735 -5030 6755
rect -5010 6735 -4990 6755
rect -4970 6735 -4950 6755
rect -4930 6735 -4910 6755
rect -4890 6735 -4870 6755
rect -4850 6735 -4830 6755
rect -4810 6735 -4790 6755
rect -4770 6735 -4750 6755
rect -3140 6695 -3120 6715
rect -3100 6695 -3080 6715
rect -3060 6695 -3040 6715
rect -3020 6695 -3000 6715
rect -4450 6653 -4430 6673
rect -4410 6653 -4390 6673
rect -4370 6653 -4350 6673
rect -4330 6653 -4310 6673
rect -4290 6653 -4270 6673
rect -4250 6653 -4230 6673
rect -4210 6653 -4190 6673
rect -4170 6653 -4150 6673
rect -4130 6653 -4110 6673
rect -4090 6653 -4070 6673
rect -4050 6653 -4030 6673
rect -4010 6653 -3990 6673
rect -3970 6653 -3950 6673
rect -3930 6653 -3910 6673
rect -3890 6653 -3870 6673
rect -3850 6653 -3830 6673
rect -3810 6653 -3790 6673
rect -3770 6653 -3750 6673
rect -3730 6653 -3710 6673
rect -3690 6653 -3670 6673
rect -3140 6615 -3120 6635
rect -3100 6615 -3080 6635
rect -3060 6615 -3040 6635
rect -3020 6615 -3000 6635
rect -5530 6571 -5510 6591
rect -5490 6571 -5470 6591
rect -5450 6571 -5430 6591
rect -5410 6571 -5390 6591
rect -5370 6571 -5350 6591
rect -5330 6571 -5310 6591
rect -5290 6571 -5270 6591
rect -5250 6571 -5230 6591
rect -5210 6571 -5190 6591
rect -5170 6571 -5150 6591
rect -5130 6571 -5110 6591
rect -5090 6571 -5070 6591
rect -5050 6571 -5030 6591
rect -5010 6571 -4990 6591
rect -4970 6571 -4950 6591
rect -4930 6571 -4910 6591
rect -4890 6571 -4870 6591
rect -4850 6571 -4830 6591
rect -4810 6571 -4790 6591
rect -4770 6571 -4750 6591
rect -3140 6530 -3120 6550
rect -3100 6530 -3080 6550
rect -3060 6530 -3040 6550
rect -3020 6530 -3000 6550
rect -4450 6489 -4430 6509
rect -4410 6489 -4390 6509
rect -4370 6489 -4350 6509
rect -4330 6489 -4310 6509
rect -4290 6489 -4270 6509
rect -4250 6489 -4230 6509
rect -4210 6489 -4190 6509
rect -4170 6489 -4150 6509
rect -4130 6489 -4110 6509
rect -4090 6489 -4070 6509
rect -4050 6489 -4030 6509
rect -4010 6489 -3990 6509
rect -3970 6489 -3950 6509
rect -3930 6489 -3910 6509
rect -3890 6489 -3870 6509
rect -3850 6489 -3830 6509
rect -3810 6489 -3790 6509
rect -3770 6489 -3750 6509
rect -3730 6489 -3710 6509
rect -3690 6489 -3670 6509
rect -3140 6450 -3120 6470
rect -3100 6450 -3080 6470
rect -3060 6450 -3040 6470
rect -3020 6450 -3000 6470
rect -5530 6407 -5510 6427
rect -5490 6407 -5470 6427
rect -5450 6407 -5430 6427
rect -5410 6407 -5390 6427
rect -5370 6407 -5350 6427
rect -5330 6407 -5310 6427
rect -5290 6407 -5270 6427
rect -5250 6407 -5230 6427
rect -5210 6407 -5190 6427
rect -5170 6407 -5150 6427
rect -5130 6407 -5110 6427
rect -5090 6407 -5070 6427
rect -5050 6407 -5030 6427
rect -5010 6407 -4990 6427
rect -4970 6407 -4950 6427
rect -4930 6407 -4910 6427
rect -4890 6407 -4870 6427
rect -4850 6407 -4830 6427
rect -4810 6407 -4790 6427
rect -4770 6407 -4750 6427
rect -3140 6370 -3120 6390
rect -3100 6370 -3080 6390
rect -3060 6370 -3040 6390
rect -3020 6370 -3000 6390
rect -4450 6325 -4430 6345
rect -4410 6325 -4390 6345
rect -4370 6325 -4350 6345
rect -4330 6325 -4310 6345
rect -4290 6325 -4270 6345
rect -4250 6325 -4230 6345
rect -4210 6325 -4190 6345
rect -4170 6325 -4150 6345
rect -4130 6325 -4110 6345
rect -4090 6325 -4070 6345
rect -4050 6325 -4030 6345
rect -4010 6325 -3990 6345
rect -3970 6325 -3950 6345
rect -3930 6325 -3910 6345
rect -3890 6325 -3870 6345
rect -3850 6325 -3830 6345
rect -3810 6325 -3790 6345
rect -3770 6325 -3750 6345
rect -3730 6325 -3710 6345
rect -3690 6325 -3670 6345
rect -4450 6285 -4430 6305
rect -4410 6285 -4390 6305
rect -4370 6285 -4350 6305
rect -4330 6285 -4310 6305
rect -4290 6285 -4270 6305
rect -4250 6285 -4230 6305
rect -4210 6285 -4190 6305
rect -4170 6285 -4150 6305
rect -4130 6285 -4110 6305
rect -4090 6285 -4070 6305
rect -4050 6285 -4030 6305
rect -4010 6285 -3990 6305
rect -3970 6285 -3950 6305
rect -3930 6285 -3910 6305
rect -3890 6285 -3870 6305
rect -3850 6285 -3830 6305
rect -3810 6285 -3790 6305
rect -3770 6285 -3750 6305
rect -3730 6285 -3710 6305
rect -3690 6285 -3670 6305
rect -370 8585 -350 8605
rect -330 8585 -310 8605
rect -290 8585 -270 8605
rect -250 8585 -230 8605
rect -210 8585 -190 8605
rect -170 8585 -150 8605
rect -130 8585 -110 8605
rect -90 8585 -70 8605
rect -50 8585 -30 8605
rect -10 8585 10 8605
rect 30 8585 50 8605
rect 70 8585 90 8605
rect 110 8585 130 8605
rect 150 8585 170 8605
rect 190 8585 210 8605
rect 230 8585 250 8605
rect 270 8585 290 8605
rect 310 8585 330 8605
rect 350 8585 370 8605
rect -1470 8500 -1450 8520
rect -1430 8500 -1410 8520
rect -1390 8500 -1370 8520
rect -1350 8500 -1330 8520
rect -1310 8500 -1290 8520
rect -1270 8500 -1250 8520
rect -1230 8500 -1210 8520
rect -1190 8500 -1170 8520
rect -1150 8500 -1130 8520
rect -1110 8500 -1090 8520
rect -1070 8500 -1050 8520
rect -1030 8500 -1010 8520
rect -990 8500 -970 8520
rect -950 8500 -930 8520
rect -910 8500 -890 8520
rect -870 8500 -850 8520
rect -830 8500 -810 8520
rect -790 8500 -770 8520
rect -750 8500 -730 8520
rect -710 8500 -690 8520
rect -1470 8457 -1450 8477
rect -1430 8457 -1410 8477
rect -1390 8457 -1370 8477
rect -1350 8457 -1330 8477
rect -1310 8457 -1290 8477
rect -1270 8457 -1250 8477
rect -1230 8457 -1210 8477
rect -1190 8457 -1170 8477
rect -1150 8457 -1130 8477
rect -1110 8457 -1090 8477
rect -1070 8457 -1050 8477
rect -1030 8457 -1010 8477
rect -990 8457 -970 8477
rect -950 8457 -930 8477
rect -910 8457 -890 8477
rect -870 8457 -850 8477
rect -830 8457 -810 8477
rect -790 8457 -770 8477
rect -750 8457 -730 8477
rect -710 8457 -690 8477
rect -2140 8415 -2120 8435
rect -2100 8415 -2080 8435
rect -2060 8415 -2040 8435
rect -2020 8415 -2000 8435
rect -390 8375 -370 8395
rect -350 8375 -330 8395
rect -310 8375 -290 8395
rect -270 8375 -250 8395
rect -230 8375 -210 8395
rect -190 8375 -170 8395
rect -150 8375 -130 8395
rect -110 8375 -90 8395
rect -70 8375 -50 8395
rect -30 8375 -10 8395
rect 10 8375 30 8395
rect 50 8375 70 8395
rect 90 8375 110 8395
rect 130 8375 150 8395
rect 170 8375 190 8395
rect 210 8375 230 8395
rect 250 8375 270 8395
rect 290 8375 310 8395
rect 330 8375 350 8395
rect 370 8375 390 8395
rect -2140 8335 -2120 8355
rect -2100 8335 -2080 8355
rect -2060 8335 -2040 8355
rect -2020 8335 -2000 8355
rect -1470 8293 -1450 8313
rect -1430 8293 -1410 8313
rect -1390 8293 -1370 8313
rect -1350 8293 -1330 8313
rect -1310 8293 -1290 8313
rect -1270 8293 -1250 8313
rect -1230 8293 -1210 8313
rect -1190 8293 -1170 8313
rect -1150 8293 -1130 8313
rect -1110 8293 -1090 8313
rect -1070 8293 -1050 8313
rect -1030 8293 -1010 8313
rect -990 8293 -970 8313
rect -950 8293 -930 8313
rect -910 8293 -890 8313
rect -870 8293 -850 8313
rect -830 8293 -810 8313
rect -790 8293 -770 8313
rect -750 8293 -730 8313
rect -710 8293 -690 8313
rect -2140 8250 -2120 8270
rect -2100 8250 -2080 8270
rect -2060 8250 -2040 8270
rect -2020 8250 -2000 8270
rect -390 8211 -370 8231
rect -350 8211 -330 8231
rect -310 8211 -290 8231
rect -270 8211 -250 8231
rect -230 8211 -210 8231
rect -190 8211 -170 8231
rect -150 8211 -130 8231
rect -110 8211 -90 8231
rect -70 8211 -50 8231
rect -30 8211 -10 8231
rect 10 8211 30 8231
rect 50 8211 70 8231
rect 90 8211 110 8231
rect 130 8211 150 8231
rect 170 8211 190 8231
rect 210 8211 230 8231
rect 250 8211 270 8231
rect 290 8211 310 8231
rect 330 8211 350 8231
rect 370 8211 390 8231
rect -2140 8170 -2120 8190
rect -2100 8170 -2080 8190
rect -2060 8170 -2040 8190
rect -2020 8170 -2000 8190
rect -1470 8129 -1450 8149
rect -1430 8129 -1410 8149
rect -1390 8129 -1370 8149
rect -1350 8129 -1330 8149
rect -1310 8129 -1290 8149
rect -1270 8129 -1250 8149
rect -1230 8129 -1210 8149
rect -1190 8129 -1170 8149
rect -1150 8129 -1130 8149
rect -1110 8129 -1090 8149
rect -1070 8129 -1050 8149
rect -1030 8129 -1010 8149
rect -990 8129 -970 8149
rect -950 8129 -930 8149
rect -910 8129 -890 8149
rect -870 8129 -850 8149
rect -830 8129 -810 8149
rect -790 8129 -770 8149
rect -750 8129 -730 8149
rect -710 8129 -690 8149
rect -2140 8090 -2120 8110
rect -2100 8090 -2080 8110
rect -2060 8090 -2040 8110
rect -2020 8090 -2000 8110
rect -390 8047 -370 8067
rect -350 8047 -330 8067
rect -310 8047 -290 8067
rect -270 8047 -250 8067
rect -230 8047 -210 8067
rect -190 8047 -170 8067
rect -150 8047 -130 8067
rect -110 8047 -90 8067
rect -70 8047 -50 8067
rect -30 8047 -10 8067
rect 10 8047 30 8067
rect 50 8047 70 8067
rect 90 8047 110 8067
rect 130 8047 150 8067
rect 170 8047 190 8067
rect 210 8047 230 8067
rect 250 8047 270 8067
rect 290 8047 310 8067
rect 330 8047 350 8067
rect 370 8047 390 8067
rect -2140 8005 -2120 8025
rect -2100 8005 -2080 8025
rect -2060 8005 -2040 8025
rect -2020 8005 -2000 8025
rect -1470 7965 -1450 7985
rect -1430 7965 -1410 7985
rect -1390 7965 -1370 7985
rect -1350 7965 -1330 7985
rect -1310 7965 -1290 7985
rect -1270 7965 -1250 7985
rect -1230 7965 -1210 7985
rect -1190 7965 -1170 7985
rect -1150 7965 -1130 7985
rect -1110 7965 -1090 7985
rect -1070 7965 -1050 7985
rect -1030 7965 -1010 7985
rect -990 7965 -970 7985
rect -950 7965 -930 7985
rect -910 7965 -890 7985
rect -870 7965 -850 7985
rect -830 7965 -810 7985
rect -790 7965 -770 7985
rect -750 7965 -730 7985
rect -710 7965 -690 7985
rect -2140 7925 -2120 7945
rect -2100 7925 -2080 7945
rect -2060 7925 -2040 7945
rect -2020 7925 -2000 7945
rect -390 7883 -370 7903
rect -350 7883 -330 7903
rect -310 7883 -290 7903
rect -270 7883 -250 7903
rect -230 7883 -210 7903
rect -190 7883 -170 7903
rect -150 7883 -130 7903
rect -110 7883 -90 7903
rect -70 7883 -50 7903
rect -30 7883 -10 7903
rect 10 7883 30 7903
rect 50 7883 70 7903
rect 90 7883 110 7903
rect 130 7883 150 7903
rect 170 7883 190 7903
rect 210 7883 230 7903
rect 250 7883 270 7903
rect 290 7883 310 7903
rect 330 7883 350 7903
rect 370 7883 390 7903
rect -2140 7840 -2120 7860
rect -2100 7840 -2080 7860
rect -2060 7840 -2040 7860
rect -2020 7840 -2000 7860
rect -1470 7801 -1450 7821
rect -1430 7801 -1410 7821
rect -1390 7801 -1370 7821
rect -1350 7801 -1330 7821
rect -1310 7801 -1290 7821
rect -1270 7801 -1250 7821
rect -1230 7801 -1210 7821
rect -1190 7801 -1170 7821
rect -1150 7801 -1130 7821
rect -1110 7801 -1090 7821
rect -1070 7801 -1050 7821
rect -1030 7801 -1010 7821
rect -990 7801 -970 7821
rect -950 7801 -930 7821
rect -910 7801 -890 7821
rect -870 7801 -850 7821
rect -830 7801 -810 7821
rect -790 7801 -770 7821
rect -750 7801 -730 7821
rect -710 7801 -690 7821
rect -2140 7760 -2120 7780
rect -2100 7760 -2080 7780
rect -2060 7760 -2040 7780
rect -2020 7760 -2000 7780
rect -390 7719 -370 7739
rect -350 7719 -330 7739
rect -310 7719 -290 7739
rect -270 7719 -250 7739
rect -230 7719 -210 7739
rect -190 7719 -170 7739
rect -150 7719 -130 7739
rect -110 7719 -90 7739
rect -70 7719 -50 7739
rect -30 7719 -10 7739
rect 10 7719 30 7739
rect 50 7719 70 7739
rect 90 7719 110 7739
rect 130 7719 150 7739
rect 170 7719 190 7739
rect 210 7719 230 7739
rect 250 7719 270 7739
rect 290 7719 310 7739
rect 330 7719 350 7739
rect 370 7719 390 7739
rect -2140 7680 -2120 7700
rect -2100 7680 -2080 7700
rect -2060 7680 -2040 7700
rect -2020 7680 -2000 7700
rect -1470 7637 -1450 7657
rect -1430 7637 -1410 7657
rect -1390 7637 -1370 7657
rect -1350 7637 -1330 7657
rect -1310 7637 -1290 7657
rect -1270 7637 -1250 7657
rect -1230 7637 -1210 7657
rect -1190 7637 -1170 7657
rect -1150 7637 -1130 7657
rect -1110 7637 -1090 7657
rect -1070 7637 -1050 7657
rect -1030 7637 -1010 7657
rect -990 7637 -970 7657
rect -950 7637 -930 7657
rect -910 7637 -890 7657
rect -870 7637 -850 7657
rect -830 7637 -810 7657
rect -790 7637 -770 7657
rect -750 7637 -730 7657
rect -710 7637 -690 7657
rect -2140 7595 -2120 7615
rect -2100 7595 -2080 7615
rect -2060 7595 -2040 7615
rect -2020 7595 -2000 7615
rect -390 7555 -370 7575
rect -350 7555 -330 7575
rect -310 7555 -290 7575
rect -270 7555 -250 7575
rect -230 7555 -210 7575
rect -190 7555 -170 7575
rect -150 7555 -130 7575
rect -110 7555 -90 7575
rect -70 7555 -50 7575
rect -30 7555 -10 7575
rect 10 7555 30 7575
rect 50 7555 70 7575
rect 90 7555 110 7575
rect 130 7555 150 7575
rect 170 7555 190 7575
rect 210 7555 230 7575
rect 250 7555 270 7575
rect 290 7555 310 7575
rect 330 7555 350 7575
rect 370 7555 390 7575
rect -2140 7515 -2120 7535
rect -2100 7515 -2080 7535
rect -2060 7515 -2040 7535
rect -2020 7515 -2000 7535
rect -1470 7473 -1450 7493
rect -1430 7473 -1410 7493
rect -1390 7473 -1370 7493
rect -1350 7473 -1330 7493
rect -1310 7473 -1290 7493
rect -1270 7473 -1250 7493
rect -1230 7473 -1210 7493
rect -1190 7473 -1170 7493
rect -1150 7473 -1130 7493
rect -1110 7473 -1090 7493
rect -1070 7473 -1050 7493
rect -1030 7473 -1010 7493
rect -990 7473 -970 7493
rect -950 7473 -930 7493
rect -910 7473 -890 7493
rect -870 7473 -850 7493
rect -830 7473 -810 7493
rect -790 7473 -770 7493
rect -750 7473 -730 7493
rect -710 7473 -690 7493
rect -2140 7430 -2120 7450
rect -2100 7430 -2080 7450
rect -2060 7430 -2040 7450
rect -2020 7430 -2000 7450
rect -390 7391 -370 7411
rect -350 7391 -330 7411
rect -310 7391 -290 7411
rect -270 7391 -250 7411
rect -230 7391 -210 7411
rect -190 7391 -170 7411
rect -150 7391 -130 7411
rect -110 7391 -90 7411
rect -70 7391 -50 7411
rect -30 7391 -10 7411
rect 10 7391 30 7411
rect 50 7391 70 7411
rect 90 7391 110 7411
rect 130 7391 150 7411
rect 170 7391 190 7411
rect 210 7391 230 7411
rect 250 7391 270 7411
rect 290 7391 310 7411
rect 330 7391 350 7411
rect 370 7391 390 7411
rect -2140 7350 -2120 7370
rect -2100 7350 -2080 7370
rect -2060 7350 -2040 7370
rect -2020 7350 -2000 7370
rect -1470 7309 -1450 7329
rect -1430 7309 -1410 7329
rect -1390 7309 -1370 7329
rect -1350 7309 -1330 7329
rect -1310 7309 -1290 7329
rect -1270 7309 -1250 7329
rect -1230 7309 -1210 7329
rect -1190 7309 -1170 7329
rect -1150 7309 -1130 7329
rect -1110 7309 -1090 7329
rect -1070 7309 -1050 7329
rect -1030 7309 -1010 7329
rect -990 7309 -970 7329
rect -950 7309 -930 7329
rect -910 7309 -890 7329
rect -870 7309 -850 7329
rect -830 7309 -810 7329
rect -790 7309 -770 7329
rect -750 7309 -730 7329
rect -710 7309 -690 7329
rect -2140 7270 -2120 7290
rect -2100 7270 -2080 7290
rect -2060 7270 -2040 7290
rect -2020 7270 -2000 7290
rect -390 7227 -370 7247
rect -350 7227 -330 7247
rect -310 7227 -290 7247
rect -270 7227 -250 7247
rect -230 7227 -210 7247
rect -190 7227 -170 7247
rect -150 7227 -130 7247
rect -110 7227 -90 7247
rect -70 7227 -50 7247
rect -30 7227 -10 7247
rect 10 7227 30 7247
rect 50 7227 70 7247
rect 90 7227 110 7247
rect 130 7227 150 7247
rect 170 7227 190 7247
rect 210 7227 230 7247
rect 250 7227 270 7247
rect 290 7227 310 7247
rect 330 7227 350 7247
rect 370 7227 390 7247
rect -2140 7185 -2120 7205
rect -2100 7185 -2080 7205
rect -2060 7185 -2040 7205
rect -2020 7185 -2000 7205
rect -1470 7145 -1450 7165
rect -1430 7145 -1410 7165
rect -1390 7145 -1370 7165
rect -1350 7145 -1330 7165
rect -1310 7145 -1290 7165
rect -1270 7145 -1250 7165
rect -1230 7145 -1210 7165
rect -1190 7145 -1170 7165
rect -1150 7145 -1130 7165
rect -1110 7145 -1090 7165
rect -1070 7145 -1050 7165
rect -1030 7145 -1010 7165
rect -990 7145 -970 7165
rect -950 7145 -930 7165
rect -910 7145 -890 7165
rect -870 7145 -850 7165
rect -830 7145 -810 7165
rect -790 7145 -770 7165
rect -750 7145 -730 7165
rect -710 7145 -690 7165
rect -2140 7105 -2120 7125
rect -2100 7105 -2080 7125
rect -2060 7105 -2040 7125
rect -2020 7105 -2000 7125
rect -390 7063 -370 7083
rect -350 7063 -330 7083
rect -310 7063 -290 7083
rect -270 7063 -250 7083
rect -230 7063 -210 7083
rect -190 7063 -170 7083
rect -150 7063 -130 7083
rect -110 7063 -90 7083
rect -70 7063 -50 7083
rect -30 7063 -10 7083
rect 10 7063 30 7083
rect 50 7063 70 7083
rect 90 7063 110 7083
rect 130 7063 150 7083
rect 170 7063 190 7083
rect 210 7063 230 7083
rect 250 7063 270 7083
rect 290 7063 310 7083
rect 330 7063 350 7083
rect 370 7063 390 7083
rect -2140 7020 -2120 7040
rect -2100 7020 -2080 7040
rect -2060 7020 -2040 7040
rect -2020 7020 -2000 7040
rect -1470 6981 -1450 7001
rect -1430 6981 -1410 7001
rect -1390 6981 -1370 7001
rect -1350 6981 -1330 7001
rect -1310 6981 -1290 7001
rect -1270 6981 -1250 7001
rect -1230 6981 -1210 7001
rect -1190 6981 -1170 7001
rect -1150 6981 -1130 7001
rect -1110 6981 -1090 7001
rect -1070 6981 -1050 7001
rect -1030 6981 -1010 7001
rect -990 6981 -970 7001
rect -950 6981 -930 7001
rect -910 6981 -890 7001
rect -870 6981 -850 7001
rect -830 6981 -810 7001
rect -790 6981 -770 7001
rect -750 6981 -730 7001
rect -710 6981 -690 7001
rect -2140 6940 -2120 6960
rect -2100 6940 -2080 6960
rect -2060 6940 -2040 6960
rect -2020 6940 -2000 6960
rect -390 6899 -370 6919
rect -350 6899 -330 6919
rect -310 6899 -290 6919
rect -270 6899 -250 6919
rect -230 6899 -210 6919
rect -190 6899 -170 6919
rect -150 6899 -130 6919
rect -110 6899 -90 6919
rect -70 6899 -50 6919
rect -30 6899 -10 6919
rect 10 6899 30 6919
rect 50 6899 70 6919
rect 90 6899 110 6919
rect 130 6899 150 6919
rect 170 6899 190 6919
rect 210 6899 230 6919
rect 250 6899 270 6919
rect 290 6899 310 6919
rect 330 6899 350 6919
rect 370 6899 390 6919
rect -2140 6860 -2120 6880
rect -2100 6860 -2080 6880
rect -2060 6860 -2040 6880
rect -2020 6860 -2000 6880
rect -1470 6817 -1450 6837
rect -1430 6817 -1410 6837
rect -1390 6817 -1370 6837
rect -1350 6817 -1330 6837
rect -1310 6817 -1290 6837
rect -1270 6817 -1250 6837
rect -1230 6817 -1210 6837
rect -1190 6817 -1170 6837
rect -1150 6817 -1130 6837
rect -1110 6817 -1090 6837
rect -1070 6817 -1050 6837
rect -1030 6817 -1010 6837
rect -990 6817 -970 6837
rect -950 6817 -930 6837
rect -910 6817 -890 6837
rect -870 6817 -850 6837
rect -830 6817 -810 6837
rect -790 6817 -770 6837
rect -750 6817 -730 6837
rect -710 6817 -690 6837
rect -2140 6775 -2120 6795
rect -2100 6775 -2080 6795
rect -2060 6775 -2040 6795
rect -2020 6775 -2000 6795
rect -390 6735 -370 6755
rect -350 6735 -330 6755
rect -310 6735 -290 6755
rect -270 6735 -250 6755
rect -230 6735 -210 6755
rect -190 6735 -170 6755
rect -150 6735 -130 6755
rect -110 6735 -90 6755
rect -70 6735 -50 6755
rect -30 6735 -10 6755
rect 10 6735 30 6755
rect 50 6735 70 6755
rect 90 6735 110 6755
rect 130 6735 150 6755
rect 170 6735 190 6755
rect 210 6735 230 6755
rect 250 6735 270 6755
rect 290 6735 310 6755
rect 330 6735 350 6755
rect 370 6735 390 6755
rect -2140 6695 -2120 6715
rect -2100 6695 -2080 6715
rect -2060 6695 -2040 6715
rect -2020 6695 -2000 6715
rect -1470 6653 -1450 6673
rect -1430 6653 -1410 6673
rect -1390 6653 -1370 6673
rect -1350 6653 -1330 6673
rect -1310 6653 -1290 6673
rect -1270 6653 -1250 6673
rect -1230 6653 -1210 6673
rect -1190 6653 -1170 6673
rect -1150 6653 -1130 6673
rect -1110 6653 -1090 6673
rect -1070 6653 -1050 6673
rect -1030 6653 -1010 6673
rect -990 6653 -970 6673
rect -950 6653 -930 6673
rect -910 6653 -890 6673
rect -870 6653 -850 6673
rect -830 6653 -810 6673
rect -790 6653 -770 6673
rect -750 6653 -730 6673
rect -710 6653 -690 6673
rect -2140 6615 -2120 6635
rect -2100 6615 -2080 6635
rect -2060 6615 -2040 6635
rect -2020 6615 -2000 6635
rect -390 6571 -370 6591
rect -350 6571 -330 6591
rect -310 6571 -290 6591
rect -270 6571 -250 6591
rect -230 6571 -210 6591
rect -190 6571 -170 6591
rect -150 6571 -130 6591
rect -110 6571 -90 6591
rect -70 6571 -50 6591
rect -30 6571 -10 6591
rect 10 6571 30 6591
rect 50 6571 70 6591
rect 90 6571 110 6591
rect 130 6571 150 6591
rect 170 6571 190 6591
rect 210 6571 230 6591
rect 250 6571 270 6591
rect 290 6571 310 6591
rect 330 6571 350 6591
rect 370 6571 390 6591
rect -2140 6530 -2120 6550
rect -2100 6530 -2080 6550
rect -2060 6530 -2040 6550
rect -2020 6530 -2000 6550
rect -1470 6489 -1450 6509
rect -1430 6489 -1410 6509
rect -1390 6489 -1370 6509
rect -1350 6489 -1330 6509
rect -1310 6489 -1290 6509
rect -1270 6489 -1250 6509
rect -1230 6489 -1210 6509
rect -1190 6489 -1170 6509
rect -1150 6489 -1130 6509
rect -1110 6489 -1090 6509
rect -1070 6489 -1050 6509
rect -1030 6489 -1010 6509
rect -990 6489 -970 6509
rect -950 6489 -930 6509
rect -910 6489 -890 6509
rect -870 6489 -850 6509
rect -830 6489 -810 6509
rect -790 6489 -770 6509
rect -750 6489 -730 6509
rect -710 6489 -690 6509
rect -2140 6450 -2120 6470
rect -2100 6450 -2080 6470
rect -2060 6450 -2040 6470
rect -2020 6450 -2000 6470
rect -390 6407 -370 6427
rect -350 6407 -330 6427
rect -310 6407 -290 6427
rect -270 6407 -250 6427
rect -230 6407 -210 6427
rect -190 6407 -170 6427
rect -150 6407 -130 6427
rect -110 6407 -90 6427
rect -70 6407 -50 6427
rect -30 6407 -10 6427
rect 10 6407 30 6427
rect 50 6407 70 6427
rect 90 6407 110 6427
rect 130 6407 150 6427
rect 170 6407 190 6427
rect 210 6407 230 6427
rect 250 6407 270 6427
rect 290 6407 310 6427
rect 330 6407 350 6427
rect 370 6407 390 6427
rect -2140 6370 -2120 6390
rect -2100 6370 -2080 6390
rect -2060 6370 -2040 6390
rect -2020 6370 -2000 6390
rect -1470 6325 -1450 6345
rect -1430 6325 -1410 6345
rect -1390 6325 -1370 6345
rect -1350 6325 -1330 6345
rect -1310 6325 -1290 6345
rect -1270 6325 -1250 6345
rect -1230 6325 -1210 6345
rect -1190 6325 -1170 6345
rect -1150 6325 -1130 6345
rect -1110 6325 -1090 6345
rect -1070 6325 -1050 6345
rect -1030 6325 -1010 6345
rect -990 6325 -970 6345
rect -950 6325 -930 6345
rect -910 6325 -890 6345
rect -870 6325 -850 6345
rect -830 6325 -810 6345
rect -790 6325 -770 6345
rect -750 6325 -730 6345
rect -710 6325 -690 6345
rect -1470 6285 -1450 6305
rect -1430 6285 -1410 6305
rect -1390 6285 -1370 6305
rect -1350 6285 -1330 6305
rect -1310 6285 -1290 6305
rect -1270 6285 -1250 6305
rect -1230 6285 -1210 6305
rect -1190 6285 -1170 6305
rect -1150 6285 -1130 6305
rect -1110 6285 -1090 6305
rect -1070 6285 -1050 6305
rect -1030 6285 -1010 6305
rect -990 6285 -970 6305
rect -950 6285 -930 6305
rect -910 6285 -890 6305
rect -870 6285 -850 6305
rect -830 6285 -810 6305
rect -790 6285 -770 6305
rect -750 6285 -730 6305
rect -710 6285 -690 6305
rect -5530 6065 -5510 6085
rect -5490 6065 -5470 6085
rect -5450 6065 -5430 6085
rect -5410 6065 -5390 6085
rect -5370 6065 -5350 6085
rect -5330 6065 -5310 6085
rect -5290 6065 -5270 6085
rect -5250 6065 -5230 6085
rect -5210 6065 -5190 6085
rect -5170 6065 -5150 6085
rect -5130 6065 -5110 6085
rect -5090 6065 -5070 6085
rect -5050 6065 -5030 6085
rect -5010 6065 -4990 6085
rect -4970 6065 -4950 6085
rect -4930 6065 -4910 6085
rect -4890 6065 -4870 6085
rect -4850 6065 -4830 6085
rect -4810 6065 -4790 6085
rect -4770 6065 -4750 6085
rect -5530 6025 -5510 6045
rect -5490 6025 -5470 6045
rect -5450 6025 -5430 6045
rect -5410 6025 -5390 6045
rect -5370 6025 -5350 6045
rect -5330 6025 -5310 6045
rect -5290 6025 -5270 6045
rect -5250 6025 -5230 6045
rect -5210 6025 -5190 6045
rect -5170 6025 -5150 6045
rect -5130 6025 -5110 6045
rect -5090 6025 -5070 6045
rect -5050 6025 -5030 6045
rect -5010 6025 -4990 6045
rect -4970 6025 -4950 6045
rect -4930 6025 -4910 6045
rect -4890 6025 -4870 6045
rect -4850 6025 -4830 6045
rect -4810 6025 -4790 6045
rect -4770 6025 -4750 6045
rect -390 6065 -370 6085
rect -350 6065 -330 6085
rect -310 6065 -290 6085
rect -270 6065 -250 6085
rect -230 6065 -210 6085
rect -190 6065 -170 6085
rect -150 6065 -130 6085
rect -110 6065 -90 6085
rect -70 6065 -50 6085
rect -30 6065 -10 6085
rect 10 6065 30 6085
rect 50 6065 70 6085
rect 90 6065 110 6085
rect 130 6065 150 6085
rect 170 6065 190 6085
rect 210 6065 230 6085
rect 250 6065 270 6085
rect 290 6065 310 6085
rect 330 6065 350 6085
rect 370 6065 390 6085
rect -390 6025 -370 6045
rect -350 6025 -330 6045
rect -310 6025 -290 6045
rect -270 6025 -250 6045
rect -230 6025 -210 6045
rect -190 6025 -170 6045
rect -150 6025 -130 6045
rect -110 6025 -90 6045
rect -70 6025 -50 6045
rect -30 6025 -10 6045
rect 10 6025 30 6045
rect 50 6025 70 6045
rect 90 6025 110 6045
rect 130 6025 150 6045
rect 170 6025 190 6045
rect 210 6025 230 6045
rect 250 6025 270 6045
rect 290 6025 310 6045
rect 330 6025 350 6045
rect 370 6025 390 6045
rect -3070 5975 -3050 6000
rect -3030 5975 -3010 6000
rect -2990 5975 -2970 6000
rect -2950 5975 -2930 6000
rect -2210 5975 -2190 6000
rect -2170 5975 -2150 6000
rect -2130 5975 -2110 6000
rect -2090 5975 -2070 6000
rect -4450 5930 -4430 5950
rect -4410 5930 -4390 5950
rect -4370 5930 -4350 5950
rect -4330 5930 -4310 5950
rect -4290 5930 -4270 5950
rect -4250 5930 -4230 5950
rect -4210 5930 -4190 5950
rect -4170 5930 -4150 5950
rect -4130 5930 -4110 5950
rect -4090 5930 -4070 5950
rect -4050 5930 -4030 5950
rect -4010 5930 -3990 5950
rect -3970 5930 -3950 5950
rect -3930 5930 -3910 5950
rect -3890 5930 -3870 5950
rect -3850 5930 -3830 5950
rect -3810 5930 -3790 5950
rect -3770 5930 -3750 5950
rect -3730 5930 -3710 5950
rect -3690 5930 -3670 5950
rect -1470 5930 -1450 5950
rect -1430 5930 -1410 5950
rect -1390 5930 -1370 5950
rect -1350 5930 -1330 5950
rect -1310 5930 -1290 5950
rect -1270 5930 -1250 5950
rect -1230 5930 -1210 5950
rect -1190 5930 -1170 5950
rect -1150 5930 -1130 5950
rect -1110 5930 -1090 5950
rect -1070 5930 -1050 5950
rect -1030 5930 -1010 5950
rect -990 5930 -970 5950
rect -950 5930 -930 5950
rect -910 5930 -890 5950
rect -870 5930 -850 5950
rect -830 5930 -810 5950
rect -790 5930 -770 5950
rect -750 5930 -730 5950
rect -710 5930 -690 5950
rect -3070 5880 -3050 5905
rect -3030 5880 -3010 5905
rect -2990 5880 -2970 5905
rect -2950 5880 -2930 5905
rect -2210 5880 -2190 5905
rect -2170 5880 -2150 5905
rect -2130 5880 -2110 5905
rect -2090 5880 -2070 5905
rect -5530 5835 -5510 5855
rect -5490 5835 -5470 5855
rect -5450 5835 -5430 5855
rect -5410 5835 -5390 5855
rect -5370 5835 -5350 5855
rect -5330 5835 -5310 5855
rect -5290 5835 -5270 5855
rect -5250 5835 -5230 5855
rect -5210 5835 -5190 5855
rect -5170 5835 -5150 5855
rect -5130 5835 -5110 5855
rect -5090 5835 -5070 5855
rect -5050 5835 -5030 5855
rect -5010 5835 -4990 5855
rect -4970 5835 -4950 5855
rect -4930 5835 -4910 5855
rect -4890 5835 -4870 5855
rect -4850 5835 -4830 5855
rect -4810 5835 -4790 5855
rect -4770 5835 -4750 5855
rect -390 5835 -370 5855
rect -350 5835 -330 5855
rect -310 5835 -290 5855
rect -270 5835 -250 5855
rect -230 5835 -210 5855
rect -190 5835 -170 5855
rect -150 5835 -130 5855
rect -110 5835 -90 5855
rect -70 5835 -50 5855
rect -30 5835 -10 5855
rect 10 5835 30 5855
rect 50 5835 70 5855
rect 90 5835 110 5855
rect 130 5835 150 5855
rect 170 5835 190 5855
rect 210 5835 230 5855
rect 250 5835 270 5855
rect 290 5835 310 5855
rect 330 5835 350 5855
rect 370 5835 390 5855
rect -3070 5785 -3050 5810
rect -3030 5785 -3010 5810
rect -2990 5785 -2970 5810
rect -2950 5785 -2930 5810
rect -2210 5785 -2190 5810
rect -2170 5785 -2150 5810
rect -2130 5785 -2110 5810
rect -2090 5785 -2070 5810
rect -4450 5740 -4430 5760
rect -4410 5740 -4390 5760
rect -4370 5740 -4350 5760
rect -4330 5740 -4310 5760
rect -4290 5740 -4270 5760
rect -4250 5740 -4230 5760
rect -4210 5740 -4190 5760
rect -4170 5740 -4150 5760
rect -4130 5740 -4110 5760
rect -4090 5740 -4070 5760
rect -4050 5740 -4030 5760
rect -4010 5740 -3990 5760
rect -3970 5740 -3950 5760
rect -3930 5740 -3910 5760
rect -3890 5740 -3870 5760
rect -3850 5740 -3830 5760
rect -3810 5740 -3790 5760
rect -3770 5740 -3750 5760
rect -3730 5740 -3710 5760
rect -3690 5740 -3670 5760
rect -1470 5740 -1450 5760
rect -1430 5740 -1410 5760
rect -1390 5740 -1370 5760
rect -1350 5740 -1330 5760
rect -1310 5740 -1290 5760
rect -1270 5740 -1250 5760
rect -1230 5740 -1210 5760
rect -1190 5740 -1170 5760
rect -1150 5740 -1130 5760
rect -1110 5740 -1090 5760
rect -1070 5740 -1050 5760
rect -1030 5740 -1010 5760
rect -990 5740 -970 5760
rect -950 5740 -930 5760
rect -910 5740 -890 5760
rect -870 5740 -850 5760
rect -830 5740 -810 5760
rect -790 5740 -770 5760
rect -750 5740 -730 5760
rect -710 5740 -690 5760
rect -3070 5690 -3050 5715
rect -3030 5690 -3010 5715
rect -2990 5690 -2970 5715
rect -2950 5690 -2930 5715
rect -2210 5690 -2190 5715
rect -2170 5690 -2150 5715
rect -2130 5690 -2110 5715
rect -2090 5690 -2070 5715
rect -5530 5645 -5510 5665
rect -5490 5645 -5470 5665
rect -5450 5645 -5430 5665
rect -5410 5645 -5390 5665
rect -5370 5645 -5350 5665
rect -5330 5645 -5310 5665
rect -5290 5645 -5270 5665
rect -5250 5645 -5230 5665
rect -5210 5645 -5190 5665
rect -5170 5645 -5150 5665
rect -5130 5645 -5110 5665
rect -5090 5645 -5070 5665
rect -5050 5645 -5030 5665
rect -5010 5645 -4990 5665
rect -4970 5645 -4950 5665
rect -4930 5645 -4910 5665
rect -4890 5645 -4870 5665
rect -4850 5645 -4830 5665
rect -4810 5645 -4790 5665
rect -4770 5645 -4750 5665
rect -390 5645 -370 5665
rect -350 5645 -330 5665
rect -310 5645 -290 5665
rect -270 5645 -250 5665
rect -230 5645 -210 5665
rect -190 5645 -170 5665
rect -150 5645 -130 5665
rect -110 5645 -90 5665
rect -70 5645 -50 5665
rect -30 5645 -10 5665
rect 10 5645 30 5665
rect 50 5645 70 5665
rect 90 5645 110 5665
rect 130 5645 150 5665
rect 170 5645 190 5665
rect 210 5645 230 5665
rect 250 5645 270 5665
rect 290 5645 310 5665
rect 330 5645 350 5665
rect 370 5645 390 5665
rect -3070 5595 -3050 5620
rect -3030 5595 -3010 5620
rect -2990 5595 -2970 5620
rect -2950 5595 -2930 5620
rect -2210 5595 -2190 5620
rect -2170 5595 -2150 5620
rect -2130 5595 -2110 5620
rect -2090 5595 -2070 5620
rect -4450 5550 -4430 5570
rect -4410 5550 -4390 5570
rect -4370 5550 -4350 5570
rect -4330 5550 -4310 5570
rect -4290 5550 -4270 5570
rect -4250 5550 -4230 5570
rect -4210 5550 -4190 5570
rect -4170 5550 -4150 5570
rect -4130 5550 -4110 5570
rect -4090 5550 -4070 5570
rect -4050 5550 -4030 5570
rect -4010 5550 -3990 5570
rect -3970 5550 -3950 5570
rect -3930 5550 -3910 5570
rect -3890 5550 -3870 5570
rect -3850 5550 -3830 5570
rect -3810 5550 -3790 5570
rect -3770 5550 -3750 5570
rect -3730 5550 -3710 5570
rect -3690 5550 -3670 5570
rect -1470 5550 -1450 5570
rect -1430 5550 -1410 5570
rect -1390 5550 -1370 5570
rect -1350 5550 -1330 5570
rect -1310 5550 -1290 5570
rect -1270 5550 -1250 5570
rect -1230 5550 -1210 5570
rect -1190 5550 -1170 5570
rect -1150 5550 -1130 5570
rect -1110 5550 -1090 5570
rect -1070 5550 -1050 5570
rect -1030 5550 -1010 5570
rect -990 5550 -970 5570
rect -950 5550 -930 5570
rect -910 5550 -890 5570
rect -870 5550 -850 5570
rect -830 5550 -810 5570
rect -790 5550 -770 5570
rect -750 5550 -730 5570
rect -710 5550 -690 5570
rect -3070 5500 -3050 5525
rect -3030 5500 -3010 5525
rect -2990 5500 -2970 5525
rect -2950 5500 -2930 5525
rect -2210 5500 -2190 5525
rect -2170 5500 -2150 5525
rect -2130 5500 -2110 5525
rect -2090 5500 -2070 5525
rect -5530 5455 -5510 5475
rect -5490 5455 -5470 5475
rect -5450 5455 -5430 5475
rect -5410 5455 -5390 5475
rect -5370 5455 -5350 5475
rect -5330 5455 -5310 5475
rect -5290 5455 -5270 5475
rect -5250 5455 -5230 5475
rect -5210 5455 -5190 5475
rect -5170 5455 -5150 5475
rect -5130 5455 -5110 5475
rect -5090 5455 -5070 5475
rect -5050 5455 -5030 5475
rect -5010 5455 -4990 5475
rect -4970 5455 -4950 5475
rect -4930 5455 -4910 5475
rect -4890 5455 -4870 5475
rect -4850 5455 -4830 5475
rect -4810 5455 -4790 5475
rect -4770 5455 -4750 5475
rect -390 5455 -370 5475
rect -350 5455 -330 5475
rect -310 5455 -290 5475
rect -270 5455 -250 5475
rect -230 5455 -210 5475
rect -190 5455 -170 5475
rect -150 5455 -130 5475
rect -110 5455 -90 5475
rect -70 5455 -50 5475
rect -30 5455 -10 5475
rect 10 5455 30 5475
rect 50 5455 70 5475
rect 90 5455 110 5475
rect 130 5455 150 5475
rect 170 5455 190 5475
rect 210 5455 230 5475
rect 250 5455 270 5475
rect 290 5455 310 5475
rect 330 5455 350 5475
rect 370 5455 390 5475
rect -3070 5405 -3050 5430
rect -3030 5405 -3010 5430
rect -2990 5405 -2970 5430
rect -2950 5405 -2930 5430
rect -2210 5405 -2190 5430
rect -2170 5405 -2150 5430
rect -2130 5405 -2110 5430
rect -2090 5405 -2070 5430
rect -4450 5360 -4430 5380
rect -4410 5360 -4390 5380
rect -4370 5360 -4350 5380
rect -4330 5360 -4310 5380
rect -4290 5360 -4270 5380
rect -4250 5360 -4230 5380
rect -4210 5360 -4190 5380
rect -4170 5360 -4150 5380
rect -4130 5360 -4110 5380
rect -4090 5360 -4070 5380
rect -4050 5360 -4030 5380
rect -4010 5360 -3990 5380
rect -3970 5360 -3950 5380
rect -3930 5360 -3910 5380
rect -3890 5360 -3870 5380
rect -3850 5360 -3830 5380
rect -3810 5360 -3790 5380
rect -3770 5360 -3750 5380
rect -3730 5360 -3710 5380
rect -3690 5360 -3670 5380
rect -1470 5360 -1450 5380
rect -1430 5360 -1410 5380
rect -1390 5360 -1370 5380
rect -1350 5360 -1330 5380
rect -1310 5360 -1290 5380
rect -1270 5360 -1250 5380
rect -1230 5360 -1210 5380
rect -1190 5360 -1170 5380
rect -1150 5360 -1130 5380
rect -1110 5360 -1090 5380
rect -1070 5360 -1050 5380
rect -1030 5360 -1010 5380
rect -990 5360 -970 5380
rect -950 5360 -930 5380
rect -910 5360 -890 5380
rect -870 5360 -850 5380
rect -830 5360 -810 5380
rect -790 5360 -770 5380
rect -750 5360 -730 5380
rect -710 5360 -690 5380
rect -3070 5310 -3050 5335
rect -3030 5310 -3010 5335
rect -2990 5310 -2970 5335
rect -2950 5310 -2930 5335
rect -2210 5310 -2190 5335
rect -2170 5310 -2150 5335
rect -2130 5310 -2110 5335
rect -2090 5310 -2070 5335
rect -5530 5265 -5510 5285
rect -5490 5265 -5470 5285
rect -5450 5265 -5430 5285
rect -5410 5265 -5390 5285
rect -5370 5265 -5350 5285
rect -5330 5265 -5310 5285
rect -5290 5265 -5270 5285
rect -5250 5265 -5230 5285
rect -5210 5265 -5190 5285
rect -5170 5265 -5150 5285
rect -5130 5265 -5110 5285
rect -5090 5265 -5070 5285
rect -5050 5265 -5030 5285
rect -5010 5265 -4990 5285
rect -4970 5265 -4950 5285
rect -4930 5265 -4910 5285
rect -4890 5265 -4870 5285
rect -4850 5265 -4830 5285
rect -4810 5265 -4790 5285
rect -4770 5265 -4750 5285
rect -390 5265 -370 5285
rect -350 5265 -330 5285
rect -310 5265 -290 5285
rect -270 5265 -250 5285
rect -230 5265 -210 5285
rect -190 5265 -170 5285
rect -150 5265 -130 5285
rect -110 5265 -90 5285
rect -70 5265 -50 5285
rect -30 5265 -10 5285
rect 10 5265 30 5285
rect 50 5265 70 5285
rect 90 5265 110 5285
rect 130 5265 150 5285
rect 170 5265 190 5285
rect 210 5265 230 5285
rect 250 5265 270 5285
rect 290 5265 310 5285
rect 330 5265 350 5285
rect 370 5265 390 5285
rect -3070 5215 -3050 5240
rect -3030 5215 -3010 5240
rect -2990 5215 -2970 5240
rect -2950 5215 -2930 5240
rect -2210 5215 -2190 5240
rect -2170 5215 -2150 5240
rect -2130 5215 -2110 5240
rect -2090 5215 -2070 5240
rect -4450 5170 -4430 5190
rect -4410 5170 -4390 5190
rect -4370 5170 -4350 5190
rect -4330 5170 -4310 5190
rect -4290 5170 -4270 5190
rect -4250 5170 -4230 5190
rect -4210 5170 -4190 5190
rect -4170 5170 -4150 5190
rect -4130 5170 -4110 5190
rect -4090 5170 -4070 5190
rect -4050 5170 -4030 5190
rect -4010 5170 -3990 5190
rect -3970 5170 -3950 5190
rect -3930 5170 -3910 5190
rect -3890 5170 -3870 5190
rect -3850 5170 -3830 5190
rect -3810 5170 -3790 5190
rect -3770 5170 -3750 5190
rect -3730 5170 -3710 5190
rect -3690 5170 -3670 5190
rect -1470 5170 -1450 5190
rect -1430 5170 -1410 5190
rect -1390 5170 -1370 5190
rect -1350 5170 -1330 5190
rect -1310 5170 -1290 5190
rect -1270 5170 -1250 5190
rect -1230 5170 -1210 5190
rect -1190 5170 -1170 5190
rect -1150 5170 -1130 5190
rect -1110 5170 -1090 5190
rect -1070 5170 -1050 5190
rect -1030 5170 -1010 5190
rect -990 5170 -970 5190
rect -950 5170 -930 5190
rect -910 5170 -890 5190
rect -870 5170 -850 5190
rect -830 5170 -810 5190
rect -790 5170 -770 5190
rect -750 5170 -730 5190
rect -710 5170 -690 5190
rect -3070 5120 -3050 5145
rect -3030 5120 -3010 5145
rect -2990 5120 -2970 5145
rect -2950 5120 -2930 5145
rect -2210 5120 -2190 5145
rect -2170 5120 -2150 5145
rect -2130 5120 -2110 5145
rect -2090 5120 -2070 5145
rect -5530 5075 -5510 5095
rect -5490 5075 -5470 5095
rect -5450 5075 -5430 5095
rect -5410 5075 -5390 5095
rect -5370 5075 -5350 5095
rect -5330 5075 -5310 5095
rect -5290 5075 -5270 5095
rect -5250 5075 -5230 5095
rect -5210 5075 -5190 5095
rect -5170 5075 -5150 5095
rect -5130 5075 -5110 5095
rect -5090 5075 -5070 5095
rect -5050 5075 -5030 5095
rect -5010 5075 -4990 5095
rect -4970 5075 -4950 5095
rect -4930 5075 -4910 5095
rect -4890 5075 -4870 5095
rect -4850 5075 -4830 5095
rect -4810 5075 -4790 5095
rect -4770 5075 -4750 5095
rect -390 5075 -370 5095
rect -350 5075 -330 5095
rect -310 5075 -290 5095
rect -270 5075 -250 5095
rect -230 5075 -210 5095
rect -190 5075 -170 5095
rect -150 5075 -130 5095
rect -110 5075 -90 5095
rect -70 5075 -50 5095
rect -30 5075 -10 5095
rect 10 5075 30 5095
rect 50 5075 70 5095
rect 90 5075 110 5095
rect 130 5075 150 5095
rect 170 5075 190 5095
rect 210 5075 230 5095
rect 250 5075 270 5095
rect 290 5075 310 5095
rect 330 5075 350 5095
rect 370 5075 390 5095
rect -3070 5025 -3050 5050
rect -3030 5025 -3010 5050
rect -2990 5025 -2970 5050
rect -2950 5025 -2930 5050
rect -2210 5025 -2190 5050
rect -2170 5025 -2150 5050
rect -2130 5025 -2110 5050
rect -2090 5025 -2070 5050
rect -4450 4980 -4430 5000
rect -4410 4980 -4390 5000
rect -4370 4980 -4350 5000
rect -4330 4980 -4310 5000
rect -4290 4980 -4270 5000
rect -4250 4980 -4230 5000
rect -4210 4980 -4190 5000
rect -4170 4980 -4150 5000
rect -4130 4980 -4110 5000
rect -4090 4980 -4070 5000
rect -4050 4980 -4030 5000
rect -4010 4980 -3990 5000
rect -3970 4980 -3950 5000
rect -3930 4980 -3910 5000
rect -3890 4980 -3870 5000
rect -3850 4980 -3830 5000
rect -3810 4980 -3790 5000
rect -3770 4980 -3750 5000
rect -3730 4980 -3710 5000
rect -3690 4980 -3670 5000
rect -1470 4980 -1450 5000
rect -1430 4980 -1410 5000
rect -1390 4980 -1370 5000
rect -1350 4980 -1330 5000
rect -1310 4980 -1290 5000
rect -1270 4980 -1250 5000
rect -1230 4980 -1210 5000
rect -1190 4980 -1170 5000
rect -1150 4980 -1130 5000
rect -1110 4980 -1090 5000
rect -1070 4980 -1050 5000
rect -1030 4980 -1010 5000
rect -990 4980 -970 5000
rect -950 4980 -930 5000
rect -910 4980 -890 5000
rect -870 4980 -850 5000
rect -830 4980 -810 5000
rect -790 4980 -770 5000
rect -750 4980 -730 5000
rect -710 4980 -690 5000
rect -3070 4930 -3050 4955
rect -3030 4930 -3010 4955
rect -2990 4930 -2970 4955
rect -2950 4930 -2930 4955
rect -2210 4930 -2190 4955
rect -2170 4930 -2150 4955
rect -2130 4930 -2110 4955
rect -2090 4930 -2070 4955
rect -5530 4885 -5510 4905
rect -5490 4885 -5470 4905
rect -5450 4885 -5430 4905
rect -5410 4885 -5390 4905
rect -5370 4885 -5350 4905
rect -5330 4885 -5310 4905
rect -5290 4885 -5270 4905
rect -5250 4885 -5230 4905
rect -5210 4885 -5190 4905
rect -5170 4885 -5150 4905
rect -5130 4885 -5110 4905
rect -5090 4885 -5070 4905
rect -5050 4885 -5030 4905
rect -5010 4885 -4990 4905
rect -4970 4885 -4950 4905
rect -4930 4885 -4910 4905
rect -4890 4885 -4870 4905
rect -4850 4885 -4830 4905
rect -4810 4885 -4790 4905
rect -4770 4885 -4750 4905
rect -390 4885 -370 4905
rect -350 4885 -330 4905
rect -310 4885 -290 4905
rect -270 4885 -250 4905
rect -230 4885 -210 4905
rect -190 4885 -170 4905
rect -150 4885 -130 4905
rect -110 4885 -90 4905
rect -70 4885 -50 4905
rect -30 4885 -10 4905
rect 10 4885 30 4905
rect 50 4885 70 4905
rect 90 4885 110 4905
rect 130 4885 150 4905
rect 170 4885 190 4905
rect 210 4885 230 4905
rect 250 4885 270 4905
rect 290 4885 310 4905
rect 330 4885 350 4905
rect 370 4885 390 4905
rect -3070 4835 -3050 4860
rect -3030 4835 -3010 4860
rect -2990 4835 -2970 4860
rect -2950 4835 -2930 4860
rect -2210 4835 -2190 4860
rect -2170 4835 -2150 4860
rect -2130 4835 -2110 4860
rect -2090 4835 -2070 4860
rect -4450 4790 -4430 4810
rect -4410 4790 -4390 4810
rect -4370 4790 -4350 4810
rect -4330 4790 -4310 4810
rect -4290 4790 -4270 4810
rect -4250 4790 -4230 4810
rect -4210 4790 -4190 4810
rect -4170 4790 -4150 4810
rect -4130 4790 -4110 4810
rect -4090 4790 -4070 4810
rect -4050 4790 -4030 4810
rect -4010 4790 -3990 4810
rect -3970 4790 -3950 4810
rect -3930 4790 -3910 4810
rect -3890 4790 -3870 4810
rect -3850 4790 -3830 4810
rect -3810 4790 -3790 4810
rect -3770 4790 -3750 4810
rect -3730 4790 -3710 4810
rect -3690 4790 -3670 4810
rect -1470 4790 -1450 4810
rect -1430 4790 -1410 4810
rect -1390 4790 -1370 4810
rect -1350 4790 -1330 4810
rect -1310 4790 -1290 4810
rect -1270 4790 -1250 4810
rect -1230 4790 -1210 4810
rect -1190 4790 -1170 4810
rect -1150 4790 -1130 4810
rect -1110 4790 -1090 4810
rect -1070 4790 -1050 4810
rect -1030 4790 -1010 4810
rect -990 4790 -970 4810
rect -950 4790 -930 4810
rect -910 4790 -890 4810
rect -870 4790 -850 4810
rect -830 4790 -810 4810
rect -790 4790 -770 4810
rect -750 4790 -730 4810
rect -710 4790 -690 4810
rect -3070 4740 -3050 4765
rect -3030 4740 -3010 4765
rect -2990 4740 -2970 4765
rect -2950 4740 -2930 4765
rect -2210 4740 -2190 4765
rect -2170 4740 -2150 4765
rect -2130 4740 -2110 4765
rect -2090 4740 -2070 4765
rect -5530 4695 -5510 4715
rect -5490 4695 -5470 4715
rect -5450 4695 -5430 4715
rect -5410 4695 -5390 4715
rect -5370 4695 -5350 4715
rect -5330 4695 -5310 4715
rect -5290 4695 -5270 4715
rect -5250 4695 -5230 4715
rect -5210 4695 -5190 4715
rect -5170 4695 -5150 4715
rect -5130 4695 -5110 4715
rect -5090 4695 -5070 4715
rect -5050 4695 -5030 4715
rect -5010 4695 -4990 4715
rect -4970 4695 -4950 4715
rect -4930 4695 -4910 4715
rect -4890 4695 -4870 4715
rect -4850 4695 -4830 4715
rect -4810 4695 -4790 4715
rect -4770 4695 -4750 4715
rect -390 4695 -370 4715
rect -350 4695 -330 4715
rect -310 4695 -290 4715
rect -270 4695 -250 4715
rect -230 4695 -210 4715
rect -190 4695 -170 4715
rect -150 4695 -130 4715
rect -110 4695 -90 4715
rect -70 4695 -50 4715
rect -30 4695 -10 4715
rect 10 4695 30 4715
rect 50 4695 70 4715
rect 90 4695 110 4715
rect 130 4695 150 4715
rect 170 4695 190 4715
rect 210 4695 230 4715
rect 250 4695 270 4715
rect 290 4695 310 4715
rect 330 4695 350 4715
rect 370 4695 390 4715
rect -3070 4645 -3050 4670
rect -3030 4645 -3010 4670
rect -2990 4645 -2970 4670
rect -2950 4645 -2930 4670
rect -2210 4645 -2190 4670
rect -2170 4645 -2150 4670
rect -2130 4645 -2110 4670
rect -2090 4645 -2070 4670
rect -4450 4600 -4430 4620
rect -4410 4600 -4390 4620
rect -4370 4600 -4350 4620
rect -4330 4600 -4310 4620
rect -4290 4600 -4270 4620
rect -4250 4600 -4230 4620
rect -4210 4600 -4190 4620
rect -4170 4600 -4150 4620
rect -4130 4600 -4110 4620
rect -4090 4600 -4070 4620
rect -4050 4600 -4030 4620
rect -4010 4600 -3990 4620
rect -3970 4600 -3950 4620
rect -3930 4600 -3910 4620
rect -3890 4600 -3870 4620
rect -3850 4600 -3830 4620
rect -3810 4600 -3790 4620
rect -3770 4600 -3750 4620
rect -3730 4600 -3710 4620
rect -3690 4600 -3670 4620
rect -1470 4600 -1450 4620
rect -1430 4600 -1410 4620
rect -1390 4600 -1370 4620
rect -1350 4600 -1330 4620
rect -1310 4600 -1290 4620
rect -1270 4600 -1250 4620
rect -1230 4600 -1210 4620
rect -1190 4600 -1170 4620
rect -1150 4600 -1130 4620
rect -1110 4600 -1090 4620
rect -1070 4600 -1050 4620
rect -1030 4600 -1010 4620
rect -990 4600 -970 4620
rect -950 4600 -930 4620
rect -910 4600 -890 4620
rect -870 4600 -850 4620
rect -830 4600 -810 4620
rect -790 4600 -770 4620
rect -750 4600 -730 4620
rect -710 4600 -690 4620
rect -3070 4550 -3050 4575
rect -3030 4550 -3010 4575
rect -2990 4550 -2970 4575
rect -2950 4550 -2930 4575
rect -2210 4550 -2190 4575
rect -2170 4550 -2150 4575
rect -2130 4550 -2110 4575
rect -2090 4550 -2070 4575
rect -5530 4505 -5510 4525
rect -5490 4505 -5470 4525
rect -5450 4505 -5430 4525
rect -5410 4505 -5390 4525
rect -5370 4505 -5350 4525
rect -5330 4505 -5310 4525
rect -5290 4505 -5270 4525
rect -5250 4505 -5230 4525
rect -5210 4505 -5190 4525
rect -5170 4505 -5150 4525
rect -5130 4505 -5110 4525
rect -5090 4505 -5070 4525
rect -5050 4505 -5030 4525
rect -5010 4505 -4990 4525
rect -4970 4505 -4950 4525
rect -4930 4505 -4910 4525
rect -4890 4505 -4870 4525
rect -4850 4505 -4830 4525
rect -4810 4505 -4790 4525
rect -4770 4505 -4750 4525
rect -390 4505 -370 4525
rect -350 4505 -330 4525
rect -310 4505 -290 4525
rect -270 4505 -250 4525
rect -230 4505 -210 4525
rect -190 4505 -170 4525
rect -150 4505 -130 4525
rect -110 4505 -90 4525
rect -70 4505 -50 4525
rect -30 4505 -10 4525
rect 10 4505 30 4525
rect 50 4505 70 4525
rect 90 4505 110 4525
rect 130 4505 150 4525
rect 170 4505 190 4525
rect 210 4505 230 4525
rect 250 4505 270 4525
rect 290 4505 310 4525
rect 330 4505 350 4525
rect 370 4505 390 4525
rect -3070 4455 -3050 4480
rect -3030 4455 -3010 4480
rect -2990 4455 -2970 4480
rect -2950 4455 -2930 4480
rect -2210 4455 -2190 4480
rect -2170 4455 -2150 4480
rect -2130 4455 -2110 4480
rect -2090 4455 -2070 4480
rect -4450 4410 -4430 4430
rect -4410 4410 -4390 4430
rect -4370 4410 -4350 4430
rect -4330 4410 -4310 4430
rect -4290 4410 -4270 4430
rect -4250 4410 -4230 4430
rect -4210 4410 -4190 4430
rect -4170 4410 -4150 4430
rect -4130 4410 -4110 4430
rect -4090 4410 -4070 4430
rect -4050 4410 -4030 4430
rect -4010 4410 -3990 4430
rect -3970 4410 -3950 4430
rect -3930 4410 -3910 4430
rect -3890 4410 -3870 4430
rect -3850 4410 -3830 4430
rect -3810 4410 -3790 4430
rect -3770 4410 -3750 4430
rect -3730 4410 -3710 4430
rect -3690 4410 -3670 4430
rect -1470 4410 -1450 4430
rect -1430 4410 -1410 4430
rect -1390 4410 -1370 4430
rect -1350 4410 -1330 4430
rect -1310 4410 -1290 4430
rect -1270 4410 -1250 4430
rect -1230 4410 -1210 4430
rect -1190 4410 -1170 4430
rect -1150 4410 -1130 4430
rect -1110 4410 -1090 4430
rect -1070 4410 -1050 4430
rect -1030 4410 -1010 4430
rect -990 4410 -970 4430
rect -950 4410 -930 4430
rect -910 4410 -890 4430
rect -870 4410 -850 4430
rect -830 4410 -810 4430
rect -790 4410 -770 4430
rect -750 4410 -730 4430
rect -710 4410 -690 4430
rect -3070 4360 -3050 4385
rect -3030 4360 -3010 4385
rect -2990 4360 -2970 4385
rect -2950 4360 -2930 4385
rect -2210 4360 -2190 4385
rect -2170 4360 -2150 4385
rect -2130 4360 -2110 4385
rect -2090 4360 -2070 4385
rect -5530 4315 -5510 4335
rect -5490 4315 -5470 4335
rect -5450 4315 -5430 4335
rect -5410 4315 -5390 4335
rect -5370 4315 -5350 4335
rect -5330 4315 -5310 4335
rect -5290 4315 -5270 4335
rect -5250 4315 -5230 4335
rect -5210 4315 -5190 4335
rect -5170 4315 -5150 4335
rect -5130 4315 -5110 4335
rect -5090 4315 -5070 4335
rect -5050 4315 -5030 4335
rect -5010 4315 -4990 4335
rect -4970 4315 -4950 4335
rect -4930 4315 -4910 4335
rect -4890 4315 -4870 4335
rect -4850 4315 -4830 4335
rect -4810 4315 -4790 4335
rect -4770 4315 -4750 4335
rect -390 4315 -370 4335
rect -350 4315 -330 4335
rect -310 4315 -290 4335
rect -270 4315 -250 4335
rect -230 4315 -210 4335
rect -190 4315 -170 4335
rect -150 4315 -130 4335
rect -110 4315 -90 4335
rect -70 4315 -50 4335
rect -30 4315 -10 4335
rect 10 4315 30 4335
rect 50 4315 70 4335
rect 90 4315 110 4335
rect 130 4315 150 4335
rect 170 4315 190 4335
rect 210 4315 230 4335
rect 250 4315 270 4335
rect 290 4315 310 4335
rect 330 4315 350 4335
rect 370 4315 390 4335
rect -3070 4265 -3050 4290
rect -3030 4265 -3010 4290
rect -2990 4265 -2970 4290
rect -2950 4265 -2930 4290
rect -2210 4265 -2190 4290
rect -2170 4265 -2150 4290
rect -2130 4265 -2110 4290
rect -2090 4265 -2070 4290
rect -4450 4220 -4430 4240
rect -4410 4220 -4390 4240
rect -4370 4220 -4350 4240
rect -4330 4220 -4310 4240
rect -4290 4220 -4270 4240
rect -4250 4220 -4230 4240
rect -4210 4220 -4190 4240
rect -4170 4220 -4150 4240
rect -4130 4220 -4110 4240
rect -4090 4220 -4070 4240
rect -4050 4220 -4030 4240
rect -4010 4220 -3990 4240
rect -3970 4220 -3950 4240
rect -3930 4220 -3910 4240
rect -3890 4220 -3870 4240
rect -3850 4220 -3830 4240
rect -3810 4220 -3790 4240
rect -3770 4220 -3750 4240
rect -3730 4220 -3710 4240
rect -3690 4220 -3670 4240
rect -1470 4220 -1450 4240
rect -1430 4220 -1410 4240
rect -1390 4220 -1370 4240
rect -1350 4220 -1330 4240
rect -1310 4220 -1290 4240
rect -1270 4220 -1250 4240
rect -1230 4220 -1210 4240
rect -1190 4220 -1170 4240
rect -1150 4220 -1130 4240
rect -1110 4220 -1090 4240
rect -1070 4220 -1050 4240
rect -1030 4220 -1010 4240
rect -990 4220 -970 4240
rect -950 4220 -930 4240
rect -910 4220 -890 4240
rect -870 4220 -850 4240
rect -830 4220 -810 4240
rect -790 4220 -770 4240
rect -750 4220 -730 4240
rect -710 4220 -690 4240
rect -3070 4170 -3050 4195
rect -3030 4170 -3010 4195
rect -2990 4170 -2970 4195
rect -2950 4170 -2930 4195
rect -2210 4170 -2190 4195
rect -2170 4170 -2150 4195
rect -2130 4170 -2110 4195
rect -2090 4170 -2070 4195
rect -5530 4125 -5510 4145
rect -5490 4125 -5470 4145
rect -5450 4125 -5430 4145
rect -5410 4125 -5390 4145
rect -5370 4125 -5350 4145
rect -5330 4125 -5310 4145
rect -5290 4125 -5270 4145
rect -5250 4125 -5230 4145
rect -5210 4125 -5190 4145
rect -5170 4125 -5150 4145
rect -5130 4125 -5110 4145
rect -5090 4125 -5070 4145
rect -5050 4125 -5030 4145
rect -5010 4125 -4990 4145
rect -4970 4125 -4950 4145
rect -4930 4125 -4910 4145
rect -4890 4125 -4870 4145
rect -4850 4125 -4830 4145
rect -4810 4125 -4790 4145
rect -4770 4125 -4750 4145
rect -390 4125 -370 4145
rect -350 4125 -330 4145
rect -310 4125 -290 4145
rect -270 4125 -250 4145
rect -230 4125 -210 4145
rect -190 4125 -170 4145
rect -150 4125 -130 4145
rect -110 4125 -90 4145
rect -70 4125 -50 4145
rect -30 4125 -10 4145
rect 10 4125 30 4145
rect 50 4125 70 4145
rect 90 4125 110 4145
rect 130 4125 150 4145
rect 170 4125 190 4145
rect 210 4125 230 4145
rect 250 4125 270 4145
rect 290 4125 310 4145
rect 330 4125 350 4145
rect 370 4125 390 4145
rect -3070 4075 -3050 4100
rect -3030 4075 -3010 4100
rect -2990 4075 -2970 4100
rect -2950 4075 -2930 4100
rect -2210 4075 -2190 4100
rect -2170 4075 -2150 4100
rect -2130 4075 -2110 4100
rect -2090 4075 -2070 4100
rect -4450 4030 -4430 4050
rect -4410 4030 -4390 4050
rect -4370 4030 -4350 4050
rect -4330 4030 -4310 4050
rect -4290 4030 -4270 4050
rect -4250 4030 -4230 4050
rect -4210 4030 -4190 4050
rect -4170 4030 -4150 4050
rect -4130 4030 -4110 4050
rect -4090 4030 -4070 4050
rect -4050 4030 -4030 4050
rect -4010 4030 -3990 4050
rect -3970 4030 -3950 4050
rect -3930 4030 -3910 4050
rect -3890 4030 -3870 4050
rect -3850 4030 -3830 4050
rect -3810 4030 -3790 4050
rect -3770 4030 -3750 4050
rect -3730 4030 -3710 4050
rect -3690 4030 -3670 4050
rect -1470 4030 -1450 4050
rect -1430 4030 -1410 4050
rect -1390 4030 -1370 4050
rect -1350 4030 -1330 4050
rect -1310 4030 -1290 4050
rect -1270 4030 -1250 4050
rect -1230 4030 -1210 4050
rect -1190 4030 -1170 4050
rect -1150 4030 -1130 4050
rect -1110 4030 -1090 4050
rect -1070 4030 -1050 4050
rect -1030 4030 -1010 4050
rect -990 4030 -970 4050
rect -950 4030 -930 4050
rect -910 4030 -890 4050
rect -870 4030 -850 4050
rect -830 4030 -810 4050
rect -790 4030 -770 4050
rect -750 4030 -730 4050
rect -710 4030 -690 4050
rect -3070 3980 -3050 4005
rect -3030 3980 -3010 4005
rect -2990 3980 -2970 4005
rect -2950 3980 -2930 4005
rect -2210 3980 -2190 4005
rect -2170 3980 -2150 4005
rect -2130 3980 -2110 4005
rect -2090 3980 -2070 4005
rect -5530 3935 -5510 3955
rect -5490 3935 -5470 3955
rect -5450 3935 -5430 3955
rect -5410 3935 -5390 3955
rect -5370 3935 -5350 3955
rect -5330 3935 -5310 3955
rect -5290 3935 -5270 3955
rect -5250 3935 -5230 3955
rect -5210 3935 -5190 3955
rect -5170 3935 -5150 3955
rect -5130 3935 -5110 3955
rect -5090 3935 -5070 3955
rect -5050 3935 -5030 3955
rect -5010 3935 -4990 3955
rect -4970 3935 -4950 3955
rect -4930 3935 -4910 3955
rect -4890 3935 -4870 3955
rect -4850 3935 -4830 3955
rect -4810 3935 -4790 3955
rect -4770 3935 -4750 3955
rect -390 3935 -370 3955
rect -350 3935 -330 3955
rect -310 3935 -290 3955
rect -270 3935 -250 3955
rect -230 3935 -210 3955
rect -190 3935 -170 3955
rect -150 3935 -130 3955
rect -110 3935 -90 3955
rect -70 3935 -50 3955
rect -30 3935 -10 3955
rect 10 3935 30 3955
rect 50 3935 70 3955
rect 90 3935 110 3955
rect 130 3935 150 3955
rect 170 3935 190 3955
rect 210 3935 230 3955
rect 250 3935 270 3955
rect 290 3935 310 3955
rect 330 3935 350 3955
rect 370 3935 390 3955
rect -3070 3885 -3050 3910
rect -3030 3885 -3010 3910
rect -2990 3885 -2970 3910
rect -2950 3885 -2930 3910
rect -2210 3885 -2190 3910
rect -2170 3885 -2150 3910
rect -2130 3885 -2110 3910
rect -2090 3885 -2070 3910
rect -4450 3840 -4430 3860
rect -4410 3840 -4390 3860
rect -4370 3840 -4350 3860
rect -4330 3840 -4310 3860
rect -4290 3840 -4270 3860
rect -4250 3840 -4230 3860
rect -4210 3840 -4190 3860
rect -4170 3840 -4150 3860
rect -4130 3840 -4110 3860
rect -4090 3840 -4070 3860
rect -4050 3840 -4030 3860
rect -4010 3840 -3990 3860
rect -3970 3840 -3950 3860
rect -3930 3840 -3910 3860
rect -3890 3840 -3870 3860
rect -3850 3840 -3830 3860
rect -3810 3840 -3790 3860
rect -3770 3840 -3750 3860
rect -3730 3840 -3710 3860
rect -3690 3840 -3670 3860
rect -1470 3840 -1450 3860
rect -1430 3840 -1410 3860
rect -1390 3840 -1370 3860
rect -1350 3840 -1330 3860
rect -1310 3840 -1290 3860
rect -1270 3840 -1250 3860
rect -1230 3840 -1210 3860
rect -1190 3840 -1170 3860
rect -1150 3840 -1130 3860
rect -1110 3840 -1090 3860
rect -1070 3840 -1050 3860
rect -1030 3840 -1010 3860
rect -990 3840 -970 3860
rect -950 3840 -930 3860
rect -910 3840 -890 3860
rect -870 3840 -850 3860
rect -830 3840 -810 3860
rect -790 3840 -770 3860
rect -750 3840 -730 3860
rect -710 3840 -690 3860
rect -3070 3790 -3050 3815
rect -3030 3790 -3010 3815
rect -2990 3790 -2970 3815
rect -2950 3790 -2930 3815
rect -2210 3790 -2190 3815
rect -2170 3790 -2150 3815
rect -2130 3790 -2110 3815
rect -2090 3790 -2070 3815
rect -5530 3745 -5510 3765
rect -5490 3745 -5470 3765
rect -5450 3745 -5430 3765
rect -5410 3745 -5390 3765
rect -5370 3745 -5350 3765
rect -5330 3745 -5310 3765
rect -5290 3745 -5270 3765
rect -5250 3745 -5230 3765
rect -5210 3745 -5190 3765
rect -5170 3745 -5150 3765
rect -5130 3745 -5110 3765
rect -5090 3745 -5070 3765
rect -5050 3745 -5030 3765
rect -5010 3745 -4990 3765
rect -4970 3745 -4950 3765
rect -4930 3745 -4910 3765
rect -4890 3745 -4870 3765
rect -4850 3745 -4830 3765
rect -4810 3745 -4790 3765
rect -4770 3745 -4750 3765
rect -390 3745 -370 3765
rect -350 3745 -330 3765
rect -310 3745 -290 3765
rect -270 3745 -250 3765
rect -230 3745 -210 3765
rect -190 3745 -170 3765
rect -150 3745 -130 3765
rect -110 3745 -90 3765
rect -70 3745 -50 3765
rect -30 3745 -10 3765
rect 10 3745 30 3765
rect 50 3745 70 3765
rect 90 3745 110 3765
rect 130 3745 150 3765
rect 170 3745 190 3765
rect 210 3745 230 3765
rect 250 3745 270 3765
rect 290 3745 310 3765
rect 330 3745 350 3765
rect 370 3745 390 3765
rect -3070 3695 -3050 3720
rect -3030 3695 -3010 3720
rect -2990 3695 -2970 3720
rect -2950 3695 -2930 3720
rect -2210 3695 -2190 3720
rect -2170 3695 -2150 3720
rect -2130 3695 -2110 3720
rect -2090 3695 -2070 3720
rect -4450 3650 -4430 3670
rect -4410 3650 -4390 3670
rect -4370 3650 -4350 3670
rect -4330 3650 -4310 3670
rect -4290 3650 -4270 3670
rect -4250 3650 -4230 3670
rect -4210 3650 -4190 3670
rect -4170 3650 -4150 3670
rect -4130 3650 -4110 3670
rect -4090 3650 -4070 3670
rect -4050 3650 -4030 3670
rect -4010 3650 -3990 3670
rect -3970 3650 -3950 3670
rect -3930 3650 -3910 3670
rect -3890 3650 -3870 3670
rect -3850 3650 -3830 3670
rect -3810 3650 -3790 3670
rect -3770 3650 -3750 3670
rect -3730 3650 -3710 3670
rect -3690 3650 -3670 3670
rect -1470 3650 -1450 3670
rect -1430 3650 -1410 3670
rect -1390 3650 -1370 3670
rect -1350 3650 -1330 3670
rect -1310 3650 -1290 3670
rect -1270 3650 -1250 3670
rect -1230 3650 -1210 3670
rect -1190 3650 -1170 3670
rect -1150 3650 -1130 3670
rect -1110 3650 -1090 3670
rect -1070 3650 -1050 3670
rect -1030 3650 -1010 3670
rect -990 3650 -970 3670
rect -950 3650 -930 3670
rect -910 3650 -890 3670
rect -870 3650 -850 3670
rect -830 3650 -810 3670
rect -790 3650 -770 3670
rect -750 3650 -730 3670
rect -710 3650 -690 3670
rect -3070 3600 -3050 3625
rect -3030 3600 -3010 3625
rect -2990 3600 -2970 3625
rect -2950 3600 -2930 3625
rect -2210 3600 -2190 3625
rect -2170 3600 -2150 3625
rect -2130 3600 -2110 3625
rect -2090 3600 -2070 3625
rect -5530 3555 -5510 3575
rect -5490 3555 -5470 3575
rect -5450 3555 -5430 3575
rect -5410 3555 -5390 3575
rect -5370 3555 -5350 3575
rect -5330 3555 -5310 3575
rect -5290 3555 -5270 3575
rect -5250 3555 -5230 3575
rect -5210 3555 -5190 3575
rect -5170 3555 -5150 3575
rect -5130 3555 -5110 3575
rect -5090 3555 -5070 3575
rect -5050 3555 -5030 3575
rect -5010 3555 -4990 3575
rect -4970 3555 -4950 3575
rect -4930 3555 -4910 3575
rect -4890 3555 -4870 3575
rect -4850 3555 -4830 3575
rect -4810 3555 -4790 3575
rect -4770 3555 -4750 3575
rect -5530 3515 -5510 3535
rect -5490 3515 -5470 3535
rect -5450 3515 -5430 3535
rect -5410 3515 -5390 3535
rect -5370 3515 -5350 3535
rect -5330 3515 -5310 3535
rect -5290 3515 -5270 3535
rect -5250 3515 -5230 3535
rect -5210 3515 -5190 3535
rect -5170 3515 -5150 3535
rect -5130 3515 -5110 3535
rect -5090 3515 -5070 3535
rect -5050 3515 -5030 3535
rect -5010 3515 -4990 3535
rect -4970 3515 -4950 3535
rect -4930 3515 -4910 3535
rect -4890 3515 -4870 3535
rect -4850 3515 -4830 3535
rect -4810 3515 -4790 3535
rect -4770 3515 -4750 3535
rect -390 3555 -370 3575
rect -350 3555 -330 3575
rect -310 3555 -290 3575
rect -270 3555 -250 3575
rect -230 3555 -210 3575
rect -190 3555 -170 3575
rect -150 3555 -130 3575
rect -110 3555 -90 3575
rect -70 3555 -50 3575
rect -30 3555 -10 3575
rect 10 3555 30 3575
rect 50 3555 70 3575
rect 90 3555 110 3575
rect 130 3555 150 3575
rect 170 3555 190 3575
rect 210 3555 230 3575
rect 250 3555 270 3575
rect 290 3555 310 3575
rect 330 3555 350 3575
rect 370 3555 390 3575
rect -390 3515 -370 3535
rect -350 3515 -330 3535
rect -310 3515 -290 3535
rect -270 3515 -250 3535
rect -230 3515 -210 3535
rect -190 3515 -170 3535
rect -150 3515 -130 3535
rect -110 3515 -90 3535
rect -70 3515 -50 3535
rect -30 3515 -10 3535
rect 10 3515 30 3535
rect 50 3515 70 3535
rect 90 3515 110 3535
rect 130 3515 150 3535
rect 170 3515 190 3535
rect 210 3515 230 3535
rect 250 3515 270 3535
rect 290 3515 310 3535
rect 330 3515 350 3535
rect 370 3515 390 3535
<< metal1 >>
rect -5540 8605 -4740 8650
rect -400 8605 400 8650
rect -5540 8585 -5510 8605
rect -5490 8585 -5470 8605
rect -5450 8585 -5430 8605
rect -5410 8585 -5390 8605
rect -5370 8585 -5350 8605
rect -5330 8585 -5310 8605
rect -5290 8585 -5270 8605
rect -5250 8585 -5230 8605
rect -5210 8585 -5190 8605
rect -5170 8585 -5150 8605
rect -5130 8585 -5110 8605
rect -5090 8585 -5070 8605
rect -5050 8585 -5030 8605
rect -5010 8585 -4990 8605
rect -4970 8585 -4950 8605
rect -4930 8585 -4910 8605
rect -4890 8585 -4870 8605
rect -4850 8585 -4830 8605
rect -4810 8585 -4790 8605
rect -4770 8585 -4740 8605
rect -4460 8585 -3660 8605
rect -1480 8585 -680 8605
rect -400 8585 -370 8605
rect -350 8585 -330 8605
rect -310 8585 -290 8605
rect -270 8585 -250 8605
rect -230 8585 -210 8605
rect -190 8585 -170 8605
rect -150 8585 -130 8605
rect -110 8585 -90 8605
rect -70 8585 -50 8605
rect -30 8585 -10 8605
rect 10 8585 30 8605
rect 50 8585 70 8605
rect 90 8585 110 8605
rect 130 8585 150 8605
rect 170 8585 190 8605
rect 210 8585 230 8605
rect 250 8585 270 8605
rect 290 8585 310 8605
rect 330 8585 350 8605
rect 370 8585 400 8605
rect -5540 8395 -4740 8585
rect -5540 8375 -5530 8395
rect -5510 8375 -5490 8395
rect -5470 8375 -5450 8395
rect -5430 8375 -5410 8395
rect -5390 8375 -5370 8395
rect -5350 8375 -5330 8395
rect -5310 8375 -5290 8395
rect -5270 8375 -5250 8395
rect -5230 8375 -5210 8395
rect -5190 8375 -5170 8395
rect -5150 8375 -5130 8395
rect -5110 8375 -5090 8395
rect -5070 8375 -5050 8395
rect -5030 8375 -5010 8395
rect -4990 8375 -4970 8395
rect -4950 8375 -4930 8395
rect -4910 8375 -4890 8395
rect -4870 8375 -4850 8395
rect -4830 8375 -4810 8395
rect -4790 8375 -4770 8395
rect -4750 8375 -4740 8395
rect -5540 8231 -4740 8375
rect -5540 8211 -5530 8231
rect -5510 8211 -5490 8231
rect -5470 8211 -5450 8231
rect -5430 8211 -5410 8231
rect -5390 8211 -5370 8231
rect -5350 8211 -5330 8231
rect -5310 8211 -5290 8231
rect -5270 8211 -5250 8231
rect -5230 8211 -5210 8231
rect -5190 8211 -5170 8231
rect -5150 8211 -5130 8231
rect -5110 8211 -5090 8231
rect -5070 8211 -5050 8231
rect -5030 8211 -5010 8231
rect -4990 8211 -4970 8231
rect -4950 8211 -4930 8231
rect -4910 8211 -4890 8231
rect -4870 8211 -4850 8231
rect -4830 8211 -4810 8231
rect -4790 8211 -4770 8231
rect -4750 8211 -4740 8231
rect -5540 8067 -4740 8211
rect -5540 8047 -5530 8067
rect -5510 8047 -5490 8067
rect -5470 8047 -5450 8067
rect -5430 8047 -5410 8067
rect -5390 8047 -5370 8067
rect -5350 8047 -5330 8067
rect -5310 8047 -5290 8067
rect -5270 8047 -5250 8067
rect -5230 8047 -5210 8067
rect -5190 8047 -5170 8067
rect -5150 8047 -5130 8067
rect -5110 8047 -5090 8067
rect -5070 8047 -5050 8067
rect -5030 8047 -5010 8067
rect -4990 8047 -4970 8067
rect -4950 8047 -4930 8067
rect -4910 8047 -4890 8067
rect -4870 8047 -4850 8067
rect -4830 8047 -4810 8067
rect -4790 8047 -4770 8067
rect -4750 8047 -4740 8067
rect -5540 7903 -4740 8047
rect -5540 7883 -5530 7903
rect -5510 7883 -5490 7903
rect -5470 7883 -5450 7903
rect -5430 7883 -5410 7903
rect -5390 7883 -5370 7903
rect -5350 7883 -5330 7903
rect -5310 7883 -5290 7903
rect -5270 7883 -5250 7903
rect -5230 7883 -5210 7903
rect -5190 7883 -5170 7903
rect -5150 7883 -5130 7903
rect -5110 7883 -5090 7903
rect -5070 7883 -5050 7903
rect -5030 7883 -5010 7903
rect -4990 7883 -4970 7903
rect -4950 7883 -4930 7903
rect -4910 7883 -4890 7903
rect -4870 7883 -4850 7903
rect -4830 7883 -4810 7903
rect -4790 7883 -4770 7903
rect -4750 7883 -4740 7903
rect -5540 7739 -4740 7883
rect -5540 7719 -5530 7739
rect -5510 7719 -5490 7739
rect -5470 7719 -5450 7739
rect -5430 7719 -5410 7739
rect -5390 7719 -5370 7739
rect -5350 7719 -5330 7739
rect -5310 7719 -5290 7739
rect -5270 7719 -5250 7739
rect -5230 7719 -5210 7739
rect -5190 7719 -5170 7739
rect -5150 7719 -5130 7739
rect -5110 7719 -5090 7739
rect -5070 7719 -5050 7739
rect -5030 7719 -5010 7739
rect -4990 7719 -4970 7739
rect -4950 7719 -4930 7739
rect -4910 7719 -4890 7739
rect -4870 7719 -4850 7739
rect -4830 7719 -4810 7739
rect -4790 7719 -4770 7739
rect -4750 7719 -4740 7739
rect -5540 7575 -4740 7719
rect -5540 7555 -5530 7575
rect -5510 7555 -5490 7575
rect -5470 7555 -5450 7575
rect -5430 7555 -5410 7575
rect -5390 7555 -5370 7575
rect -5350 7555 -5330 7575
rect -5310 7555 -5290 7575
rect -5270 7555 -5250 7575
rect -5230 7555 -5210 7575
rect -5190 7555 -5170 7575
rect -5150 7555 -5130 7575
rect -5110 7555 -5090 7575
rect -5070 7555 -5050 7575
rect -5030 7555 -5010 7575
rect -4990 7555 -4970 7575
rect -4950 7555 -4930 7575
rect -4910 7555 -4890 7575
rect -4870 7555 -4850 7575
rect -4830 7555 -4810 7575
rect -4790 7555 -4770 7575
rect -4750 7555 -4740 7575
rect -5540 7411 -4740 7555
rect -5540 7391 -5530 7411
rect -5510 7391 -5490 7411
rect -5470 7391 -5450 7411
rect -5430 7391 -5410 7411
rect -5390 7391 -5370 7411
rect -5350 7391 -5330 7411
rect -5310 7391 -5290 7411
rect -5270 7391 -5250 7411
rect -5230 7391 -5210 7411
rect -5190 7391 -5170 7411
rect -5150 7391 -5130 7411
rect -5110 7391 -5090 7411
rect -5070 7391 -5050 7411
rect -5030 7391 -5010 7411
rect -4990 7391 -4970 7411
rect -4950 7391 -4930 7411
rect -4910 7391 -4890 7411
rect -4870 7391 -4850 7411
rect -4830 7391 -4810 7411
rect -4790 7391 -4770 7411
rect -4750 7391 -4740 7411
rect -5540 7247 -4740 7391
rect -5540 7227 -5530 7247
rect -5510 7227 -5490 7247
rect -5470 7227 -5450 7247
rect -5430 7227 -5410 7247
rect -5390 7227 -5370 7247
rect -5350 7227 -5330 7247
rect -5310 7227 -5290 7247
rect -5270 7227 -5250 7247
rect -5230 7227 -5210 7247
rect -5190 7227 -5170 7247
rect -5150 7227 -5130 7247
rect -5110 7227 -5090 7247
rect -5070 7227 -5050 7247
rect -5030 7227 -5010 7247
rect -4990 7227 -4970 7247
rect -4950 7227 -4930 7247
rect -4910 7227 -4890 7247
rect -4870 7227 -4850 7247
rect -4830 7227 -4810 7247
rect -4790 7227 -4770 7247
rect -4750 7227 -4740 7247
rect -5540 7083 -4740 7227
rect -5540 7063 -5530 7083
rect -5510 7063 -5490 7083
rect -5470 7063 -5450 7083
rect -5430 7063 -5410 7083
rect -5390 7063 -5370 7083
rect -5350 7063 -5330 7083
rect -5310 7063 -5290 7083
rect -5270 7063 -5250 7083
rect -5230 7063 -5210 7083
rect -5190 7063 -5170 7083
rect -5150 7063 -5130 7083
rect -5110 7063 -5090 7083
rect -5070 7063 -5050 7083
rect -5030 7063 -5010 7083
rect -4990 7063 -4970 7083
rect -4950 7063 -4930 7083
rect -4910 7063 -4890 7083
rect -4870 7063 -4850 7083
rect -4830 7063 -4810 7083
rect -4790 7063 -4770 7083
rect -4750 7063 -4740 7083
rect -5540 6919 -4740 7063
rect -5540 6899 -5530 6919
rect -5510 6899 -5490 6919
rect -5470 6899 -5450 6919
rect -5430 6899 -5410 6919
rect -5390 6899 -5370 6919
rect -5350 6899 -5330 6919
rect -5310 6899 -5290 6919
rect -5270 6899 -5250 6919
rect -5230 6899 -5210 6919
rect -5190 6899 -5170 6919
rect -5150 6899 -5130 6919
rect -5110 6899 -5090 6919
rect -5070 6899 -5050 6919
rect -5030 6899 -5010 6919
rect -4990 6899 -4970 6919
rect -4950 6899 -4930 6919
rect -4910 6899 -4890 6919
rect -4870 6899 -4850 6919
rect -4830 6899 -4810 6919
rect -4790 6899 -4770 6919
rect -4750 6899 -4740 6919
rect -5540 6755 -4740 6899
rect -5540 6735 -5530 6755
rect -5510 6735 -5490 6755
rect -5470 6735 -5450 6755
rect -5430 6735 -5410 6755
rect -5390 6735 -5370 6755
rect -5350 6735 -5330 6755
rect -5310 6735 -5290 6755
rect -5270 6735 -5250 6755
rect -5230 6735 -5210 6755
rect -5190 6735 -5170 6755
rect -5150 6735 -5130 6755
rect -5110 6735 -5090 6755
rect -5070 6735 -5050 6755
rect -5030 6735 -5010 6755
rect -4990 6735 -4970 6755
rect -4950 6735 -4930 6755
rect -4910 6735 -4890 6755
rect -4870 6735 -4850 6755
rect -4830 6735 -4810 6755
rect -4790 6735 -4770 6755
rect -4750 6735 -4740 6755
rect -5540 6591 -4740 6735
rect -5540 6571 -5530 6591
rect -5510 6571 -5490 6591
rect -5470 6571 -5450 6591
rect -5430 6571 -5410 6591
rect -5390 6571 -5370 6591
rect -5350 6571 -5330 6591
rect -5310 6571 -5290 6591
rect -5270 6571 -5250 6591
rect -5230 6571 -5210 6591
rect -5190 6571 -5170 6591
rect -5150 6571 -5130 6591
rect -5110 6571 -5090 6591
rect -5070 6571 -5050 6591
rect -5030 6571 -5010 6591
rect -4990 6571 -4970 6591
rect -4950 6571 -4930 6591
rect -4910 6571 -4890 6591
rect -4870 6571 -4850 6591
rect -4830 6571 -4810 6591
rect -4790 6571 -4770 6591
rect -4750 6571 -4740 6591
rect -5540 6427 -4740 6571
rect -5540 6407 -5530 6427
rect -5510 6407 -5490 6427
rect -5470 6407 -5450 6427
rect -5430 6407 -5410 6427
rect -5390 6407 -5370 6427
rect -5350 6407 -5330 6427
rect -5310 6407 -5290 6427
rect -5270 6407 -5250 6427
rect -5230 6407 -5210 6427
rect -5190 6407 -5170 6427
rect -5150 6407 -5130 6427
rect -5110 6407 -5090 6427
rect -5070 6407 -5050 6427
rect -5030 6407 -5010 6427
rect -4990 6407 -4970 6427
rect -4950 6407 -4930 6427
rect -4910 6407 -4890 6427
rect -4870 6407 -4850 6427
rect -4830 6407 -4810 6427
rect -4790 6407 -4770 6427
rect -4750 6407 -4740 6427
rect -5540 6275 -4740 6407
rect -4460 8520 -3660 8530
rect -4460 8500 -4450 8520
rect -4430 8500 -4410 8520
rect -4390 8500 -4370 8520
rect -4350 8500 -4330 8520
rect -4310 8500 -4290 8520
rect -4270 8500 -4250 8520
rect -4230 8500 -4210 8520
rect -4190 8500 -4170 8520
rect -4150 8500 -4130 8520
rect -4110 8500 -4090 8520
rect -4070 8500 -4050 8520
rect -4030 8500 -4010 8520
rect -3990 8500 -3970 8520
rect -3950 8500 -3930 8520
rect -3910 8500 -3890 8520
rect -3870 8500 -3850 8520
rect -3830 8500 -3810 8520
rect -3790 8500 -3770 8520
rect -3750 8500 -3730 8520
rect -3710 8500 -3690 8520
rect -3670 8500 -3660 8520
rect -4460 8477 -3660 8500
rect -4460 8457 -4450 8477
rect -4430 8457 -4410 8477
rect -4390 8457 -4370 8477
rect -4350 8457 -4330 8477
rect -4310 8457 -4290 8477
rect -4270 8457 -4250 8477
rect -4230 8457 -4210 8477
rect -4190 8457 -4170 8477
rect -4150 8457 -4130 8477
rect -4110 8457 -4090 8477
rect -4070 8457 -4050 8477
rect -4030 8457 -4010 8477
rect -3990 8457 -3970 8477
rect -3950 8457 -3930 8477
rect -3910 8457 -3890 8477
rect -3870 8457 -3850 8477
rect -3830 8457 -3810 8477
rect -3790 8457 -3770 8477
rect -3750 8457 -3730 8477
rect -3710 8457 -3690 8477
rect -3670 8457 -3660 8477
rect -4460 8313 -3660 8457
rect -1480 8520 -680 8530
rect -1480 8500 -1470 8520
rect -1450 8500 -1430 8520
rect -1410 8500 -1390 8520
rect -1370 8500 -1350 8520
rect -1330 8500 -1310 8520
rect -1290 8500 -1270 8520
rect -1250 8500 -1230 8520
rect -1210 8500 -1190 8520
rect -1170 8500 -1150 8520
rect -1130 8500 -1110 8520
rect -1090 8500 -1070 8520
rect -1050 8500 -1030 8520
rect -1010 8500 -990 8520
rect -970 8500 -950 8520
rect -930 8500 -910 8520
rect -890 8500 -870 8520
rect -850 8500 -830 8520
rect -810 8500 -790 8520
rect -770 8500 -750 8520
rect -730 8500 -710 8520
rect -690 8500 -680 8520
rect -1480 8477 -680 8500
rect -1480 8457 -1470 8477
rect -1450 8457 -1430 8477
rect -1410 8457 -1390 8477
rect -1370 8457 -1350 8477
rect -1330 8457 -1310 8477
rect -1290 8457 -1270 8477
rect -1250 8457 -1230 8477
rect -1210 8457 -1190 8477
rect -1170 8457 -1150 8477
rect -1130 8457 -1110 8477
rect -1090 8457 -1070 8477
rect -1050 8457 -1030 8477
rect -1010 8457 -990 8477
rect -970 8457 -950 8477
rect -930 8457 -910 8477
rect -890 8457 -870 8477
rect -850 8457 -830 8477
rect -810 8457 -790 8477
rect -770 8457 -750 8477
rect -730 8457 -710 8477
rect -690 8457 -680 8477
rect -4460 8293 -4450 8313
rect -4430 8293 -4410 8313
rect -4390 8293 -4370 8313
rect -4350 8293 -4330 8313
rect -4310 8293 -4290 8313
rect -4270 8293 -4250 8313
rect -4230 8293 -4210 8313
rect -4190 8293 -4170 8313
rect -4150 8293 -4130 8313
rect -4110 8293 -4090 8313
rect -4070 8293 -4050 8313
rect -4030 8293 -4010 8313
rect -3990 8293 -3970 8313
rect -3950 8293 -3930 8313
rect -3910 8293 -3890 8313
rect -3870 8293 -3850 8313
rect -3830 8293 -3810 8313
rect -3790 8293 -3770 8313
rect -3750 8293 -3730 8313
rect -3710 8293 -3690 8313
rect -3670 8293 -3660 8313
rect -4460 8149 -3660 8293
rect -4460 8129 -4450 8149
rect -4430 8129 -4410 8149
rect -4390 8129 -4370 8149
rect -4350 8129 -4330 8149
rect -4310 8129 -4290 8149
rect -4270 8129 -4250 8149
rect -4230 8129 -4210 8149
rect -4190 8129 -4170 8149
rect -4150 8129 -4130 8149
rect -4110 8129 -4090 8149
rect -4070 8129 -4050 8149
rect -4030 8129 -4010 8149
rect -3990 8129 -3970 8149
rect -3950 8129 -3930 8149
rect -3910 8129 -3890 8149
rect -3870 8129 -3850 8149
rect -3830 8129 -3810 8149
rect -3790 8129 -3770 8149
rect -3750 8129 -3730 8149
rect -3710 8129 -3690 8149
rect -3670 8129 -3660 8149
rect -4460 7985 -3660 8129
rect -4460 7965 -4450 7985
rect -4430 7965 -4410 7985
rect -4390 7965 -4370 7985
rect -4350 7965 -4330 7985
rect -4310 7965 -4290 7985
rect -4270 7965 -4250 7985
rect -4230 7965 -4210 7985
rect -4190 7965 -4170 7985
rect -4150 7965 -4130 7985
rect -4110 7965 -4090 7985
rect -4070 7965 -4050 7985
rect -4030 7965 -4010 7985
rect -3990 7965 -3970 7985
rect -3950 7965 -3930 7985
rect -3910 7965 -3890 7985
rect -3870 7965 -3850 7985
rect -3830 7965 -3810 7985
rect -3790 7965 -3770 7985
rect -3750 7965 -3730 7985
rect -3710 7965 -3690 7985
rect -3670 7965 -3660 7985
rect -4460 7821 -3660 7965
rect -4460 7801 -4450 7821
rect -4430 7801 -4410 7821
rect -4390 7801 -4370 7821
rect -4350 7801 -4330 7821
rect -4310 7801 -4290 7821
rect -4270 7801 -4250 7821
rect -4230 7801 -4210 7821
rect -4190 7801 -4170 7821
rect -4150 7801 -4130 7821
rect -4110 7801 -4090 7821
rect -4070 7801 -4050 7821
rect -4030 7801 -4010 7821
rect -3990 7801 -3970 7821
rect -3950 7801 -3930 7821
rect -3910 7801 -3890 7821
rect -3870 7801 -3850 7821
rect -3830 7801 -3810 7821
rect -3790 7801 -3770 7821
rect -3750 7801 -3730 7821
rect -3710 7801 -3690 7821
rect -3670 7801 -3660 7821
rect -4460 7657 -3660 7801
rect -4460 7637 -4450 7657
rect -4430 7637 -4410 7657
rect -4390 7637 -4370 7657
rect -4350 7637 -4330 7657
rect -4310 7637 -4290 7657
rect -4270 7637 -4250 7657
rect -4230 7637 -4210 7657
rect -4190 7637 -4170 7657
rect -4150 7637 -4130 7657
rect -4110 7637 -4090 7657
rect -4070 7637 -4050 7657
rect -4030 7637 -4010 7657
rect -3990 7637 -3970 7657
rect -3950 7637 -3930 7657
rect -3910 7637 -3890 7657
rect -3870 7637 -3850 7657
rect -3830 7637 -3810 7657
rect -3790 7637 -3770 7657
rect -3750 7637 -3730 7657
rect -3710 7637 -3690 7657
rect -3670 7637 -3660 7657
rect -4460 7493 -3660 7637
rect -4460 7473 -4450 7493
rect -4430 7473 -4410 7493
rect -4390 7473 -4370 7493
rect -4350 7473 -4330 7493
rect -4310 7473 -4290 7493
rect -4270 7473 -4250 7493
rect -4230 7473 -4210 7493
rect -4190 7473 -4170 7493
rect -4150 7473 -4130 7493
rect -4110 7473 -4090 7493
rect -4070 7473 -4050 7493
rect -4030 7473 -4010 7493
rect -3990 7473 -3970 7493
rect -3950 7473 -3930 7493
rect -3910 7473 -3890 7493
rect -3870 7473 -3850 7493
rect -3830 7473 -3810 7493
rect -3790 7473 -3770 7493
rect -3750 7473 -3730 7493
rect -3710 7473 -3690 7493
rect -3670 7473 -3660 7493
rect -4460 7329 -3660 7473
rect -4460 7309 -4450 7329
rect -4430 7309 -4410 7329
rect -4390 7309 -4370 7329
rect -4350 7309 -4330 7329
rect -4310 7309 -4290 7329
rect -4270 7309 -4250 7329
rect -4230 7309 -4210 7329
rect -4190 7309 -4170 7329
rect -4150 7309 -4130 7329
rect -4110 7309 -4090 7329
rect -4070 7309 -4050 7329
rect -4030 7309 -4010 7329
rect -3990 7309 -3970 7329
rect -3950 7309 -3930 7329
rect -3910 7309 -3890 7329
rect -3870 7309 -3850 7329
rect -3830 7309 -3810 7329
rect -3790 7309 -3770 7329
rect -3750 7309 -3730 7329
rect -3710 7309 -3690 7329
rect -3670 7309 -3660 7329
rect -4460 7165 -3660 7309
rect -4460 7145 -4450 7165
rect -4430 7145 -4410 7165
rect -4390 7145 -4370 7165
rect -4350 7145 -4330 7165
rect -4310 7145 -4290 7165
rect -4270 7145 -4250 7165
rect -4230 7145 -4210 7165
rect -4190 7145 -4170 7165
rect -4150 7145 -4130 7165
rect -4110 7145 -4090 7165
rect -4070 7145 -4050 7165
rect -4030 7145 -4010 7165
rect -3990 7145 -3970 7165
rect -3950 7145 -3930 7165
rect -3910 7145 -3890 7165
rect -3870 7145 -3850 7165
rect -3830 7145 -3810 7165
rect -3790 7145 -3770 7165
rect -3750 7145 -3730 7165
rect -3710 7145 -3690 7165
rect -3670 7145 -3660 7165
rect -4460 7001 -3660 7145
rect -4460 6981 -4450 7001
rect -4430 6981 -4410 7001
rect -4390 6981 -4370 7001
rect -4350 6981 -4330 7001
rect -4310 6981 -4290 7001
rect -4270 6981 -4250 7001
rect -4230 6981 -4210 7001
rect -4190 6981 -4170 7001
rect -4150 6981 -4130 7001
rect -4110 6981 -4090 7001
rect -4070 6981 -4050 7001
rect -4030 6981 -4010 7001
rect -3990 6981 -3970 7001
rect -3950 6981 -3930 7001
rect -3910 6981 -3890 7001
rect -3870 6981 -3850 7001
rect -3830 6981 -3810 7001
rect -3790 6981 -3770 7001
rect -3750 6981 -3730 7001
rect -3710 6981 -3690 7001
rect -3670 6981 -3660 7001
rect -4460 6837 -3660 6981
rect -4460 6817 -4450 6837
rect -4430 6817 -4410 6837
rect -4390 6817 -4370 6837
rect -4350 6817 -4330 6837
rect -4310 6817 -4290 6837
rect -4270 6817 -4250 6837
rect -4230 6817 -4210 6837
rect -4190 6817 -4170 6837
rect -4150 6817 -4130 6837
rect -4110 6817 -4090 6837
rect -4070 6817 -4050 6837
rect -4030 6817 -4010 6837
rect -3990 6817 -3970 6837
rect -3950 6817 -3930 6837
rect -3910 6817 -3890 6837
rect -3870 6817 -3850 6837
rect -3830 6817 -3810 6837
rect -3790 6817 -3770 6837
rect -3750 6817 -3730 6837
rect -3710 6817 -3690 6837
rect -3670 6817 -3660 6837
rect -4460 6673 -3660 6817
rect -4460 6653 -4450 6673
rect -4430 6653 -4410 6673
rect -4390 6653 -4370 6673
rect -4350 6653 -4330 6673
rect -4310 6653 -4290 6673
rect -4270 6653 -4250 6673
rect -4230 6653 -4210 6673
rect -4190 6653 -4170 6673
rect -4150 6653 -4130 6673
rect -4110 6653 -4090 6673
rect -4070 6653 -4050 6673
rect -4030 6653 -4010 6673
rect -3990 6653 -3970 6673
rect -3950 6653 -3930 6673
rect -3910 6653 -3890 6673
rect -3870 6653 -3850 6673
rect -3830 6653 -3810 6673
rect -3790 6653 -3770 6673
rect -3750 6653 -3730 6673
rect -3710 6653 -3690 6673
rect -3670 6653 -3660 6673
rect -4460 6509 -3660 6653
rect -4460 6489 -4450 6509
rect -4430 6489 -4410 6509
rect -4390 6489 -4370 6509
rect -4350 6489 -4330 6509
rect -4310 6489 -4290 6509
rect -4270 6489 -4250 6509
rect -4230 6489 -4210 6509
rect -4190 6489 -4170 6509
rect -4150 6489 -4130 6509
rect -4110 6489 -4090 6509
rect -4070 6489 -4050 6509
rect -4030 6489 -4010 6509
rect -3990 6489 -3970 6509
rect -3950 6489 -3930 6509
rect -3910 6489 -3890 6509
rect -3870 6489 -3850 6509
rect -3830 6489 -3810 6509
rect -3790 6489 -3770 6509
rect -3750 6489 -3730 6509
rect -3710 6489 -3690 6509
rect -3670 6489 -3660 6509
rect -4460 6345 -3660 6489
rect -3155 8435 -2990 8445
rect -3155 8415 -3140 8435
rect -3120 8415 -3100 8435
rect -3080 8415 -3060 8435
rect -3040 8415 -3020 8435
rect -3000 8415 -2990 8435
rect -3155 8355 -2990 8415
rect -3155 8335 -3140 8355
rect -3120 8335 -3100 8355
rect -3080 8335 -3060 8355
rect -3040 8335 -3020 8355
rect -3000 8335 -2990 8355
rect -3155 8270 -2990 8335
rect -3155 8250 -3140 8270
rect -3120 8250 -3100 8270
rect -3080 8250 -3060 8270
rect -3040 8250 -3020 8270
rect -3000 8250 -2990 8270
rect -3155 8190 -2990 8250
rect -3155 8170 -3140 8190
rect -3120 8170 -3100 8190
rect -3080 8170 -3060 8190
rect -3040 8170 -3020 8190
rect -3000 8170 -2990 8190
rect -3155 8110 -2990 8170
rect -3155 8090 -3140 8110
rect -3120 8090 -3100 8110
rect -3080 8090 -3060 8110
rect -3040 8090 -3020 8110
rect -3000 8090 -2990 8110
rect -3155 8025 -2990 8090
rect -3155 8005 -3140 8025
rect -3120 8005 -3100 8025
rect -3080 8005 -3060 8025
rect -3040 8005 -3020 8025
rect -3000 8005 -2990 8025
rect -3155 7945 -2990 8005
rect -3155 7925 -3140 7945
rect -3120 7925 -3100 7945
rect -3080 7925 -3060 7945
rect -3040 7925 -3020 7945
rect -3000 7925 -2990 7945
rect -3155 7860 -2990 7925
rect -3155 7840 -3140 7860
rect -3120 7840 -3100 7860
rect -3080 7840 -3060 7860
rect -3040 7840 -3020 7860
rect -3000 7840 -2990 7860
rect -3155 7780 -2990 7840
rect -3155 7760 -3140 7780
rect -3120 7760 -3100 7780
rect -3080 7760 -3060 7780
rect -3040 7760 -3020 7780
rect -3000 7760 -2990 7780
rect -3155 7700 -2990 7760
rect -3155 7680 -3140 7700
rect -3120 7680 -3100 7700
rect -3080 7680 -3060 7700
rect -3040 7680 -3020 7700
rect -3000 7680 -2990 7700
rect -3155 7615 -2990 7680
rect -3155 7595 -3140 7615
rect -3120 7595 -3100 7615
rect -3080 7595 -3060 7615
rect -3040 7595 -3020 7615
rect -3000 7595 -2990 7615
rect -3155 7535 -2990 7595
rect -3155 7515 -3140 7535
rect -3120 7515 -3100 7535
rect -3080 7515 -3060 7535
rect -3040 7515 -3020 7535
rect -3000 7515 -2990 7535
rect -3155 7450 -2990 7515
rect -3155 7430 -3140 7450
rect -3120 7430 -3100 7450
rect -3080 7430 -3060 7450
rect -3040 7430 -3020 7450
rect -3000 7430 -2990 7450
rect -3155 7370 -2990 7430
rect -3155 7350 -3140 7370
rect -3120 7350 -3100 7370
rect -3080 7350 -3060 7370
rect -3040 7350 -3020 7370
rect -3000 7350 -2990 7370
rect -3155 7290 -2990 7350
rect -3155 7270 -3140 7290
rect -3120 7270 -3100 7290
rect -3080 7270 -3060 7290
rect -3040 7270 -3020 7290
rect -3000 7270 -2990 7290
rect -3155 7205 -2990 7270
rect -3155 7185 -3140 7205
rect -3120 7185 -3100 7205
rect -3080 7185 -3060 7205
rect -3040 7185 -3020 7205
rect -3000 7185 -2990 7205
rect -3155 7125 -2990 7185
rect -3155 7105 -3140 7125
rect -3120 7105 -3100 7125
rect -3080 7105 -3060 7125
rect -3040 7105 -3020 7125
rect -3000 7105 -2990 7125
rect -3155 7040 -2990 7105
rect -3155 7020 -3140 7040
rect -3120 7020 -3100 7040
rect -3080 7020 -3060 7040
rect -3040 7020 -3020 7040
rect -3000 7020 -2990 7040
rect -3155 6960 -2990 7020
rect -3155 6940 -3140 6960
rect -3120 6940 -3100 6960
rect -3080 6940 -3060 6960
rect -3040 6940 -3020 6960
rect -3000 6940 -2990 6960
rect -3155 6880 -2990 6940
rect -3155 6860 -3140 6880
rect -3120 6860 -3100 6880
rect -3080 6860 -3060 6880
rect -3040 6860 -3020 6880
rect -3000 6860 -2990 6880
rect -3155 6795 -2990 6860
rect -3155 6775 -3140 6795
rect -3120 6775 -3100 6795
rect -3080 6775 -3060 6795
rect -3040 6775 -3020 6795
rect -3000 6775 -2990 6795
rect -3155 6715 -2990 6775
rect -3155 6695 -3140 6715
rect -3120 6695 -3100 6715
rect -3080 6695 -3060 6715
rect -3040 6695 -3020 6715
rect -3000 6695 -2990 6715
rect -3155 6635 -2990 6695
rect -3155 6615 -3140 6635
rect -3120 6615 -3100 6635
rect -3080 6615 -3060 6635
rect -3040 6615 -3020 6635
rect -3000 6615 -2990 6635
rect -3155 6550 -2990 6615
rect -3155 6530 -3140 6550
rect -3120 6530 -3100 6550
rect -3080 6530 -3060 6550
rect -3040 6530 -3020 6550
rect -3000 6530 -2990 6550
rect -3155 6470 -2990 6530
rect -3155 6450 -3140 6470
rect -3120 6450 -3100 6470
rect -3080 6450 -3060 6470
rect -3040 6450 -3020 6470
rect -3000 6450 -2990 6470
rect -3155 6390 -2990 6450
rect -3155 6370 -3140 6390
rect -3120 6370 -3100 6390
rect -3080 6370 -3060 6390
rect -3040 6370 -3020 6390
rect -3000 6370 -2990 6390
rect -3155 6360 -2990 6370
rect -2150 8435 -1985 8445
rect -2150 8415 -2140 8435
rect -2120 8415 -2100 8435
rect -2080 8415 -2060 8435
rect -2040 8415 -2020 8435
rect -2000 8415 -1985 8435
rect -2150 8355 -1985 8415
rect -2150 8335 -2140 8355
rect -2120 8335 -2100 8355
rect -2080 8335 -2060 8355
rect -2040 8335 -2020 8355
rect -2000 8335 -1985 8355
rect -2150 8270 -1985 8335
rect -2150 8250 -2140 8270
rect -2120 8250 -2100 8270
rect -2080 8250 -2060 8270
rect -2040 8250 -2020 8270
rect -2000 8250 -1985 8270
rect -2150 8190 -1985 8250
rect -2150 8170 -2140 8190
rect -2120 8170 -2100 8190
rect -2080 8170 -2060 8190
rect -2040 8170 -2020 8190
rect -2000 8170 -1985 8190
rect -2150 8110 -1985 8170
rect -2150 8090 -2140 8110
rect -2120 8090 -2100 8110
rect -2080 8090 -2060 8110
rect -2040 8090 -2020 8110
rect -2000 8090 -1985 8110
rect -2150 8025 -1985 8090
rect -2150 8005 -2140 8025
rect -2120 8005 -2100 8025
rect -2080 8005 -2060 8025
rect -2040 8005 -2020 8025
rect -2000 8005 -1985 8025
rect -2150 7945 -1985 8005
rect -2150 7925 -2140 7945
rect -2120 7925 -2100 7945
rect -2080 7925 -2060 7945
rect -2040 7925 -2020 7945
rect -2000 7925 -1985 7945
rect -2150 7860 -1985 7925
rect -2150 7840 -2140 7860
rect -2120 7840 -2100 7860
rect -2080 7840 -2060 7860
rect -2040 7840 -2020 7860
rect -2000 7840 -1985 7860
rect -2150 7780 -1985 7840
rect -2150 7760 -2140 7780
rect -2120 7760 -2100 7780
rect -2080 7760 -2060 7780
rect -2040 7760 -2020 7780
rect -2000 7760 -1985 7780
rect -2150 7700 -1985 7760
rect -2150 7680 -2140 7700
rect -2120 7680 -2100 7700
rect -2080 7680 -2060 7700
rect -2040 7680 -2020 7700
rect -2000 7680 -1985 7700
rect -2150 7615 -1985 7680
rect -2150 7595 -2140 7615
rect -2120 7595 -2100 7615
rect -2080 7595 -2060 7615
rect -2040 7595 -2020 7615
rect -2000 7595 -1985 7615
rect -2150 7535 -1985 7595
rect -2150 7515 -2140 7535
rect -2120 7515 -2100 7535
rect -2080 7515 -2060 7535
rect -2040 7515 -2020 7535
rect -2000 7515 -1985 7535
rect -2150 7450 -1985 7515
rect -2150 7430 -2140 7450
rect -2120 7430 -2100 7450
rect -2080 7430 -2060 7450
rect -2040 7430 -2020 7450
rect -2000 7430 -1985 7450
rect -2150 7370 -1985 7430
rect -2150 7350 -2140 7370
rect -2120 7350 -2100 7370
rect -2080 7350 -2060 7370
rect -2040 7350 -2020 7370
rect -2000 7350 -1985 7370
rect -2150 7290 -1985 7350
rect -2150 7270 -2140 7290
rect -2120 7270 -2100 7290
rect -2080 7270 -2060 7290
rect -2040 7270 -2020 7290
rect -2000 7270 -1985 7290
rect -2150 7205 -1985 7270
rect -2150 7185 -2140 7205
rect -2120 7185 -2100 7205
rect -2080 7185 -2060 7205
rect -2040 7185 -2020 7205
rect -2000 7185 -1985 7205
rect -2150 7125 -1985 7185
rect -2150 7105 -2140 7125
rect -2120 7105 -2100 7125
rect -2080 7105 -2060 7125
rect -2040 7105 -2020 7125
rect -2000 7105 -1985 7125
rect -2150 7040 -1985 7105
rect -2150 7020 -2140 7040
rect -2120 7020 -2100 7040
rect -2080 7020 -2060 7040
rect -2040 7020 -2020 7040
rect -2000 7020 -1985 7040
rect -2150 6960 -1985 7020
rect -2150 6940 -2140 6960
rect -2120 6940 -2100 6960
rect -2080 6940 -2060 6960
rect -2040 6940 -2020 6960
rect -2000 6940 -1985 6960
rect -2150 6880 -1985 6940
rect -2150 6860 -2140 6880
rect -2120 6860 -2100 6880
rect -2080 6860 -2060 6880
rect -2040 6860 -2020 6880
rect -2000 6860 -1985 6880
rect -2150 6795 -1985 6860
rect -2150 6775 -2140 6795
rect -2120 6775 -2100 6795
rect -2080 6775 -2060 6795
rect -2040 6775 -2020 6795
rect -2000 6775 -1985 6795
rect -2150 6715 -1985 6775
rect -2150 6695 -2140 6715
rect -2120 6695 -2100 6715
rect -2080 6695 -2060 6715
rect -2040 6695 -2020 6715
rect -2000 6695 -1985 6715
rect -2150 6635 -1985 6695
rect -2150 6615 -2140 6635
rect -2120 6615 -2100 6635
rect -2080 6615 -2060 6635
rect -2040 6615 -2020 6635
rect -2000 6615 -1985 6635
rect -2150 6550 -1985 6615
rect -2150 6530 -2140 6550
rect -2120 6530 -2100 6550
rect -2080 6530 -2060 6550
rect -2040 6530 -2020 6550
rect -2000 6530 -1985 6550
rect -2150 6470 -1985 6530
rect -2150 6450 -2140 6470
rect -2120 6450 -2100 6470
rect -2080 6450 -2060 6470
rect -2040 6450 -2020 6470
rect -2000 6450 -1985 6470
rect -2150 6390 -1985 6450
rect -2150 6370 -2140 6390
rect -2120 6370 -2100 6390
rect -2080 6370 -2060 6390
rect -2040 6370 -2020 6390
rect -2000 6370 -1985 6390
rect -2150 6360 -1985 6370
rect -1480 8313 -680 8457
rect -1480 8293 -1470 8313
rect -1450 8293 -1430 8313
rect -1410 8293 -1390 8313
rect -1370 8293 -1350 8313
rect -1330 8293 -1310 8313
rect -1290 8293 -1270 8313
rect -1250 8293 -1230 8313
rect -1210 8293 -1190 8313
rect -1170 8293 -1150 8313
rect -1130 8293 -1110 8313
rect -1090 8293 -1070 8313
rect -1050 8293 -1030 8313
rect -1010 8293 -990 8313
rect -970 8293 -950 8313
rect -930 8293 -910 8313
rect -890 8293 -870 8313
rect -850 8293 -830 8313
rect -810 8293 -790 8313
rect -770 8293 -750 8313
rect -730 8293 -710 8313
rect -690 8293 -680 8313
rect -1480 8149 -680 8293
rect -1480 8129 -1470 8149
rect -1450 8129 -1430 8149
rect -1410 8129 -1390 8149
rect -1370 8129 -1350 8149
rect -1330 8129 -1310 8149
rect -1290 8129 -1270 8149
rect -1250 8129 -1230 8149
rect -1210 8129 -1190 8149
rect -1170 8129 -1150 8149
rect -1130 8129 -1110 8149
rect -1090 8129 -1070 8149
rect -1050 8129 -1030 8149
rect -1010 8129 -990 8149
rect -970 8129 -950 8149
rect -930 8129 -910 8149
rect -890 8129 -870 8149
rect -850 8129 -830 8149
rect -810 8129 -790 8149
rect -770 8129 -750 8149
rect -730 8129 -710 8149
rect -690 8129 -680 8149
rect -1480 7985 -680 8129
rect -1480 7965 -1470 7985
rect -1450 7965 -1430 7985
rect -1410 7965 -1390 7985
rect -1370 7965 -1350 7985
rect -1330 7965 -1310 7985
rect -1290 7965 -1270 7985
rect -1250 7965 -1230 7985
rect -1210 7965 -1190 7985
rect -1170 7965 -1150 7985
rect -1130 7965 -1110 7985
rect -1090 7965 -1070 7985
rect -1050 7965 -1030 7985
rect -1010 7965 -990 7985
rect -970 7965 -950 7985
rect -930 7965 -910 7985
rect -890 7965 -870 7985
rect -850 7965 -830 7985
rect -810 7965 -790 7985
rect -770 7965 -750 7985
rect -730 7965 -710 7985
rect -690 7965 -680 7985
rect -1480 7821 -680 7965
rect -1480 7801 -1470 7821
rect -1450 7801 -1430 7821
rect -1410 7801 -1390 7821
rect -1370 7801 -1350 7821
rect -1330 7801 -1310 7821
rect -1290 7801 -1270 7821
rect -1250 7801 -1230 7821
rect -1210 7801 -1190 7821
rect -1170 7801 -1150 7821
rect -1130 7801 -1110 7821
rect -1090 7801 -1070 7821
rect -1050 7801 -1030 7821
rect -1010 7801 -990 7821
rect -970 7801 -950 7821
rect -930 7801 -910 7821
rect -890 7801 -870 7821
rect -850 7801 -830 7821
rect -810 7801 -790 7821
rect -770 7801 -750 7821
rect -730 7801 -710 7821
rect -690 7801 -680 7821
rect -1480 7657 -680 7801
rect -1480 7637 -1470 7657
rect -1450 7637 -1430 7657
rect -1410 7637 -1390 7657
rect -1370 7637 -1350 7657
rect -1330 7637 -1310 7657
rect -1290 7637 -1270 7657
rect -1250 7637 -1230 7657
rect -1210 7637 -1190 7657
rect -1170 7637 -1150 7657
rect -1130 7637 -1110 7657
rect -1090 7637 -1070 7657
rect -1050 7637 -1030 7657
rect -1010 7637 -990 7657
rect -970 7637 -950 7657
rect -930 7637 -910 7657
rect -890 7637 -870 7657
rect -850 7637 -830 7657
rect -810 7637 -790 7657
rect -770 7637 -750 7657
rect -730 7637 -710 7657
rect -690 7637 -680 7657
rect -1480 7493 -680 7637
rect -1480 7473 -1470 7493
rect -1450 7473 -1430 7493
rect -1410 7473 -1390 7493
rect -1370 7473 -1350 7493
rect -1330 7473 -1310 7493
rect -1290 7473 -1270 7493
rect -1250 7473 -1230 7493
rect -1210 7473 -1190 7493
rect -1170 7473 -1150 7493
rect -1130 7473 -1110 7493
rect -1090 7473 -1070 7493
rect -1050 7473 -1030 7493
rect -1010 7473 -990 7493
rect -970 7473 -950 7493
rect -930 7473 -910 7493
rect -890 7473 -870 7493
rect -850 7473 -830 7493
rect -810 7473 -790 7493
rect -770 7473 -750 7493
rect -730 7473 -710 7493
rect -690 7473 -680 7493
rect -1480 7329 -680 7473
rect -1480 7309 -1470 7329
rect -1450 7309 -1430 7329
rect -1410 7309 -1390 7329
rect -1370 7309 -1350 7329
rect -1330 7309 -1310 7329
rect -1290 7309 -1270 7329
rect -1250 7309 -1230 7329
rect -1210 7309 -1190 7329
rect -1170 7309 -1150 7329
rect -1130 7309 -1110 7329
rect -1090 7309 -1070 7329
rect -1050 7309 -1030 7329
rect -1010 7309 -990 7329
rect -970 7309 -950 7329
rect -930 7309 -910 7329
rect -890 7309 -870 7329
rect -850 7309 -830 7329
rect -810 7309 -790 7329
rect -770 7309 -750 7329
rect -730 7309 -710 7329
rect -690 7309 -680 7329
rect -1480 7165 -680 7309
rect -1480 7145 -1470 7165
rect -1450 7145 -1430 7165
rect -1410 7145 -1390 7165
rect -1370 7145 -1350 7165
rect -1330 7145 -1310 7165
rect -1290 7145 -1270 7165
rect -1250 7145 -1230 7165
rect -1210 7145 -1190 7165
rect -1170 7145 -1150 7165
rect -1130 7145 -1110 7165
rect -1090 7145 -1070 7165
rect -1050 7145 -1030 7165
rect -1010 7145 -990 7165
rect -970 7145 -950 7165
rect -930 7145 -910 7165
rect -890 7145 -870 7165
rect -850 7145 -830 7165
rect -810 7145 -790 7165
rect -770 7145 -750 7165
rect -730 7145 -710 7165
rect -690 7145 -680 7165
rect -1480 7001 -680 7145
rect -1480 6981 -1470 7001
rect -1450 6981 -1430 7001
rect -1410 6981 -1390 7001
rect -1370 6981 -1350 7001
rect -1330 6981 -1310 7001
rect -1290 6981 -1270 7001
rect -1250 6981 -1230 7001
rect -1210 6981 -1190 7001
rect -1170 6981 -1150 7001
rect -1130 6981 -1110 7001
rect -1090 6981 -1070 7001
rect -1050 6981 -1030 7001
rect -1010 6981 -990 7001
rect -970 6981 -950 7001
rect -930 6981 -910 7001
rect -890 6981 -870 7001
rect -850 6981 -830 7001
rect -810 6981 -790 7001
rect -770 6981 -750 7001
rect -730 6981 -710 7001
rect -690 6981 -680 7001
rect -1480 6837 -680 6981
rect -1480 6817 -1470 6837
rect -1450 6817 -1430 6837
rect -1410 6817 -1390 6837
rect -1370 6817 -1350 6837
rect -1330 6817 -1310 6837
rect -1290 6817 -1270 6837
rect -1250 6817 -1230 6837
rect -1210 6817 -1190 6837
rect -1170 6817 -1150 6837
rect -1130 6817 -1110 6837
rect -1090 6817 -1070 6837
rect -1050 6817 -1030 6837
rect -1010 6817 -990 6837
rect -970 6817 -950 6837
rect -930 6817 -910 6837
rect -890 6817 -870 6837
rect -850 6817 -830 6837
rect -810 6817 -790 6837
rect -770 6817 -750 6837
rect -730 6817 -710 6837
rect -690 6817 -680 6837
rect -1480 6673 -680 6817
rect -1480 6653 -1470 6673
rect -1450 6653 -1430 6673
rect -1410 6653 -1390 6673
rect -1370 6653 -1350 6673
rect -1330 6653 -1310 6673
rect -1290 6653 -1270 6673
rect -1250 6653 -1230 6673
rect -1210 6653 -1190 6673
rect -1170 6653 -1150 6673
rect -1130 6653 -1110 6673
rect -1090 6653 -1070 6673
rect -1050 6653 -1030 6673
rect -1010 6653 -990 6673
rect -970 6653 -950 6673
rect -930 6653 -910 6673
rect -890 6653 -870 6673
rect -850 6653 -830 6673
rect -810 6653 -790 6673
rect -770 6653 -750 6673
rect -730 6653 -710 6673
rect -690 6653 -680 6673
rect -1480 6509 -680 6653
rect -1480 6489 -1470 6509
rect -1450 6489 -1430 6509
rect -1410 6489 -1390 6509
rect -1370 6489 -1350 6509
rect -1330 6489 -1310 6509
rect -1290 6489 -1270 6509
rect -1250 6489 -1230 6509
rect -1210 6489 -1190 6509
rect -1170 6489 -1150 6509
rect -1130 6489 -1110 6509
rect -1090 6489 -1070 6509
rect -1050 6489 -1030 6509
rect -1010 6489 -990 6509
rect -970 6489 -950 6509
rect -930 6489 -910 6509
rect -890 6489 -870 6509
rect -850 6489 -830 6509
rect -810 6489 -790 6509
rect -770 6489 -750 6509
rect -730 6489 -710 6509
rect -690 6489 -680 6509
rect -4460 6325 -4450 6345
rect -4430 6325 -4410 6345
rect -4390 6325 -4370 6345
rect -4350 6325 -4330 6345
rect -4310 6325 -4290 6345
rect -4270 6325 -4250 6345
rect -4230 6325 -4210 6345
rect -4190 6325 -4170 6345
rect -4150 6325 -4130 6345
rect -4110 6325 -4090 6345
rect -4070 6325 -4050 6345
rect -4030 6325 -4010 6345
rect -3990 6325 -3970 6345
rect -3950 6325 -3930 6345
rect -3910 6325 -3890 6345
rect -3870 6325 -3850 6345
rect -3830 6325 -3810 6345
rect -3790 6325 -3770 6345
rect -3750 6325 -3730 6345
rect -3710 6325 -3690 6345
rect -3670 6325 -3660 6345
rect -4460 6305 -3660 6325
rect -4460 6285 -4450 6305
rect -4430 6285 -4410 6305
rect -4390 6285 -4370 6305
rect -4350 6285 -4330 6305
rect -4310 6285 -4290 6305
rect -4270 6285 -4250 6305
rect -4230 6285 -4210 6305
rect -4190 6285 -4170 6305
rect -4150 6285 -4130 6305
rect -4110 6285 -4090 6305
rect -4070 6285 -4050 6305
rect -4030 6285 -4010 6305
rect -3990 6285 -3970 6305
rect -3950 6285 -3930 6305
rect -3910 6285 -3890 6305
rect -3870 6285 -3850 6305
rect -3830 6285 -3810 6305
rect -3790 6285 -3770 6305
rect -3750 6285 -3730 6305
rect -3710 6285 -3690 6305
rect -3670 6285 -3660 6305
rect -5540 6085 -4740 6095
rect -5540 6065 -5530 6085
rect -5510 6065 -5490 6085
rect -5470 6065 -5450 6085
rect -5430 6065 -5410 6085
rect -5390 6065 -5370 6085
rect -5350 6065 -5330 6085
rect -5310 6065 -5290 6085
rect -5270 6065 -5250 6085
rect -5230 6065 -5210 6085
rect -5190 6065 -5170 6085
rect -5150 6065 -5130 6085
rect -5110 6065 -5090 6085
rect -5070 6065 -5050 6085
rect -5030 6065 -5010 6085
rect -4990 6065 -4970 6085
rect -4950 6065 -4930 6085
rect -4910 6065 -4890 6085
rect -4870 6065 -4850 6085
rect -4830 6065 -4810 6085
rect -4790 6065 -4770 6085
rect -4750 6065 -4740 6085
rect -5540 6045 -4740 6065
rect -5540 6025 -5530 6045
rect -5510 6025 -5490 6045
rect -5470 6025 -5450 6045
rect -5430 6025 -5410 6045
rect -5390 6025 -5370 6045
rect -5350 6025 -5330 6045
rect -5310 6025 -5290 6045
rect -5270 6025 -5250 6045
rect -5230 6025 -5210 6045
rect -5190 6025 -5170 6045
rect -5150 6025 -5130 6045
rect -5110 6025 -5090 6045
rect -5070 6025 -5050 6045
rect -5030 6025 -5010 6045
rect -4990 6025 -4970 6045
rect -4950 6025 -4930 6045
rect -4910 6025 -4890 6045
rect -4870 6025 -4850 6045
rect -4830 6025 -4810 6045
rect -4790 6025 -4770 6045
rect -4750 6025 -4740 6045
rect -5540 5855 -4740 6025
rect -5540 5835 -5530 5855
rect -5510 5835 -5490 5855
rect -5470 5835 -5450 5855
rect -5430 5835 -5410 5855
rect -5390 5835 -5370 5855
rect -5350 5835 -5330 5855
rect -5310 5835 -5290 5855
rect -5270 5835 -5250 5855
rect -5230 5835 -5210 5855
rect -5190 5835 -5170 5855
rect -5150 5835 -5130 5855
rect -5110 5835 -5090 5855
rect -5070 5835 -5050 5855
rect -5030 5835 -5010 5855
rect -4990 5835 -4970 5855
rect -4950 5835 -4930 5855
rect -4910 5835 -4890 5855
rect -4870 5835 -4850 5855
rect -4830 5835 -4810 5855
rect -4790 5835 -4770 5855
rect -4750 5835 -4740 5855
rect -5540 5665 -4740 5835
rect -5540 5645 -5530 5665
rect -5510 5645 -5490 5665
rect -5470 5645 -5450 5665
rect -5430 5645 -5410 5665
rect -5390 5645 -5370 5665
rect -5350 5645 -5330 5665
rect -5310 5645 -5290 5665
rect -5270 5645 -5250 5665
rect -5230 5645 -5210 5665
rect -5190 5645 -5170 5665
rect -5150 5645 -5130 5665
rect -5110 5645 -5090 5665
rect -5070 5645 -5050 5665
rect -5030 5645 -5010 5665
rect -4990 5645 -4970 5665
rect -4950 5645 -4930 5665
rect -4910 5645 -4890 5665
rect -4870 5645 -4850 5665
rect -4830 5645 -4810 5665
rect -4790 5645 -4770 5665
rect -4750 5645 -4740 5665
rect -5540 5475 -4740 5645
rect -5540 5455 -5530 5475
rect -5510 5455 -5490 5475
rect -5470 5455 -5450 5475
rect -5430 5455 -5410 5475
rect -5390 5455 -5370 5475
rect -5350 5455 -5330 5475
rect -5310 5455 -5290 5475
rect -5270 5455 -5250 5475
rect -5230 5455 -5210 5475
rect -5190 5455 -5170 5475
rect -5150 5455 -5130 5475
rect -5110 5455 -5090 5475
rect -5070 5455 -5050 5475
rect -5030 5455 -5010 5475
rect -4990 5455 -4970 5475
rect -4950 5455 -4930 5475
rect -4910 5455 -4890 5475
rect -4870 5455 -4850 5475
rect -4830 5455 -4810 5475
rect -4790 5455 -4770 5475
rect -4750 5455 -4740 5475
rect -5540 5285 -4740 5455
rect -5540 5265 -5530 5285
rect -5510 5265 -5490 5285
rect -5470 5265 -5450 5285
rect -5430 5265 -5410 5285
rect -5390 5265 -5370 5285
rect -5350 5265 -5330 5285
rect -5310 5265 -5290 5285
rect -5270 5265 -5250 5285
rect -5230 5265 -5210 5285
rect -5190 5265 -5170 5285
rect -5150 5265 -5130 5285
rect -5110 5265 -5090 5285
rect -5070 5265 -5050 5285
rect -5030 5265 -5010 5285
rect -4990 5265 -4970 5285
rect -4950 5265 -4930 5285
rect -4910 5265 -4890 5285
rect -4870 5265 -4850 5285
rect -4830 5265 -4810 5285
rect -4790 5265 -4770 5285
rect -4750 5265 -4740 5285
rect -5540 5095 -4740 5265
rect -5540 5075 -5530 5095
rect -5510 5075 -5490 5095
rect -5470 5075 -5450 5095
rect -5430 5075 -5410 5095
rect -5390 5075 -5370 5095
rect -5350 5075 -5330 5095
rect -5310 5075 -5290 5095
rect -5270 5075 -5250 5095
rect -5230 5075 -5210 5095
rect -5190 5075 -5170 5095
rect -5150 5075 -5130 5095
rect -5110 5075 -5090 5095
rect -5070 5075 -5050 5095
rect -5030 5075 -5010 5095
rect -4990 5075 -4970 5095
rect -4950 5075 -4930 5095
rect -4910 5075 -4890 5095
rect -4870 5075 -4850 5095
rect -4830 5075 -4810 5095
rect -4790 5075 -4770 5095
rect -4750 5075 -4740 5095
rect -5540 4905 -4740 5075
rect -5540 4885 -5530 4905
rect -5510 4885 -5490 4905
rect -5470 4885 -5450 4905
rect -5430 4885 -5410 4905
rect -5390 4885 -5370 4905
rect -5350 4885 -5330 4905
rect -5310 4885 -5290 4905
rect -5270 4885 -5250 4905
rect -5230 4885 -5210 4905
rect -5190 4885 -5170 4905
rect -5150 4885 -5130 4905
rect -5110 4885 -5090 4905
rect -5070 4885 -5050 4905
rect -5030 4885 -5010 4905
rect -4990 4885 -4970 4905
rect -4950 4885 -4930 4905
rect -4910 4885 -4890 4905
rect -4870 4885 -4850 4905
rect -4830 4885 -4810 4905
rect -4790 4885 -4770 4905
rect -4750 4885 -4740 4905
rect -5540 4715 -4740 4885
rect -5540 4695 -5530 4715
rect -5510 4695 -5490 4715
rect -5470 4695 -5450 4715
rect -5430 4695 -5410 4715
rect -5390 4695 -5370 4715
rect -5350 4695 -5330 4715
rect -5310 4695 -5290 4715
rect -5270 4695 -5250 4715
rect -5230 4695 -5210 4715
rect -5190 4695 -5170 4715
rect -5150 4695 -5130 4715
rect -5110 4695 -5090 4715
rect -5070 4695 -5050 4715
rect -5030 4695 -5010 4715
rect -4990 4695 -4970 4715
rect -4950 4695 -4930 4715
rect -4910 4695 -4890 4715
rect -4870 4695 -4850 4715
rect -4830 4695 -4810 4715
rect -4790 4695 -4770 4715
rect -4750 4695 -4740 4715
rect -5540 4525 -4740 4695
rect -5540 4505 -5530 4525
rect -5510 4505 -5490 4525
rect -5470 4505 -5450 4525
rect -5430 4505 -5410 4525
rect -5390 4505 -5370 4525
rect -5350 4505 -5330 4525
rect -5310 4505 -5290 4525
rect -5270 4505 -5250 4525
rect -5230 4505 -5210 4525
rect -5190 4505 -5170 4525
rect -5150 4505 -5130 4525
rect -5110 4505 -5090 4525
rect -5070 4505 -5050 4525
rect -5030 4505 -5010 4525
rect -4990 4505 -4970 4525
rect -4950 4505 -4930 4525
rect -4910 4505 -4890 4525
rect -4870 4505 -4850 4525
rect -4830 4505 -4810 4525
rect -4790 4505 -4770 4525
rect -4750 4505 -4740 4525
rect -5540 4335 -4740 4505
rect -5540 4315 -5530 4335
rect -5510 4315 -5490 4335
rect -5470 4315 -5450 4335
rect -5430 4315 -5410 4335
rect -5390 4315 -5370 4335
rect -5350 4315 -5330 4335
rect -5310 4315 -5290 4335
rect -5270 4315 -5250 4335
rect -5230 4315 -5210 4335
rect -5190 4315 -5170 4335
rect -5150 4315 -5130 4335
rect -5110 4315 -5090 4335
rect -5070 4315 -5050 4335
rect -5030 4315 -5010 4335
rect -4990 4315 -4970 4335
rect -4950 4315 -4930 4335
rect -4910 4315 -4890 4335
rect -4870 4315 -4850 4335
rect -4830 4315 -4810 4335
rect -4790 4315 -4770 4335
rect -4750 4315 -4740 4335
rect -5540 4145 -4740 4315
rect -5540 4125 -5530 4145
rect -5510 4125 -5490 4145
rect -5470 4125 -5450 4145
rect -5430 4125 -5410 4145
rect -5390 4125 -5370 4145
rect -5350 4125 -5330 4145
rect -5310 4125 -5290 4145
rect -5270 4125 -5250 4145
rect -5230 4125 -5210 4145
rect -5190 4125 -5170 4145
rect -5150 4125 -5130 4145
rect -5110 4125 -5090 4145
rect -5070 4125 -5050 4145
rect -5030 4125 -5010 4145
rect -4990 4125 -4970 4145
rect -4950 4125 -4930 4145
rect -4910 4125 -4890 4145
rect -4870 4125 -4850 4145
rect -4830 4125 -4810 4145
rect -4790 4125 -4770 4145
rect -4750 4125 -4740 4145
rect -5540 3955 -4740 4125
rect -5540 3935 -5530 3955
rect -5510 3935 -5490 3955
rect -5470 3935 -5450 3955
rect -5430 3935 -5410 3955
rect -5390 3935 -5370 3955
rect -5350 3935 -5330 3955
rect -5310 3935 -5290 3955
rect -5270 3935 -5250 3955
rect -5230 3935 -5210 3955
rect -5190 3935 -5170 3955
rect -5150 3935 -5130 3955
rect -5110 3935 -5090 3955
rect -5070 3935 -5050 3955
rect -5030 3935 -5010 3955
rect -4990 3935 -4970 3955
rect -4950 3935 -4930 3955
rect -4910 3935 -4890 3955
rect -4870 3935 -4850 3955
rect -4830 3935 -4810 3955
rect -4790 3935 -4770 3955
rect -4750 3935 -4740 3955
rect -5540 3765 -4740 3935
rect -5540 3745 -5530 3765
rect -5510 3745 -5490 3765
rect -5470 3745 -5450 3765
rect -5430 3745 -5410 3765
rect -5390 3745 -5370 3765
rect -5350 3745 -5330 3765
rect -5310 3745 -5290 3765
rect -5270 3745 -5250 3765
rect -5230 3745 -5210 3765
rect -5190 3745 -5170 3765
rect -5150 3745 -5130 3765
rect -5110 3745 -5090 3765
rect -5070 3745 -5050 3765
rect -5030 3745 -5010 3765
rect -4990 3745 -4970 3765
rect -4950 3745 -4930 3765
rect -4910 3745 -4890 3765
rect -4870 3745 -4850 3765
rect -4830 3745 -4810 3765
rect -4790 3745 -4770 3765
rect -4750 3745 -4740 3765
rect -5540 3575 -4740 3745
rect -4460 5950 -3660 6285
rect -1480 6345 -680 6489
rect -1480 6325 -1470 6345
rect -1450 6325 -1430 6345
rect -1410 6325 -1390 6345
rect -1370 6325 -1350 6345
rect -1330 6325 -1310 6345
rect -1290 6325 -1270 6345
rect -1250 6325 -1230 6345
rect -1210 6325 -1190 6345
rect -1170 6325 -1150 6345
rect -1130 6325 -1110 6345
rect -1090 6325 -1070 6345
rect -1050 6325 -1030 6345
rect -1010 6325 -990 6345
rect -970 6325 -950 6345
rect -930 6325 -910 6345
rect -890 6325 -870 6345
rect -850 6325 -830 6345
rect -810 6325 -790 6345
rect -770 6325 -750 6345
rect -730 6325 -710 6345
rect -690 6325 -680 6345
rect -1480 6305 -680 6325
rect -1480 6285 -1470 6305
rect -1450 6285 -1430 6305
rect -1410 6285 -1390 6305
rect -1370 6285 -1350 6305
rect -1330 6285 -1310 6305
rect -1290 6285 -1270 6305
rect -1250 6285 -1230 6305
rect -1210 6285 -1190 6305
rect -1170 6285 -1150 6305
rect -1130 6285 -1110 6305
rect -1090 6285 -1070 6305
rect -1050 6285 -1030 6305
rect -1010 6285 -990 6305
rect -970 6285 -950 6305
rect -930 6285 -910 6305
rect -890 6285 -870 6305
rect -850 6285 -830 6305
rect -810 6285 -790 6305
rect -770 6285 -750 6305
rect -730 6285 -710 6305
rect -690 6285 -680 6305
rect -4460 5930 -4450 5950
rect -4430 5930 -4410 5950
rect -4390 5930 -4370 5950
rect -4350 5930 -4330 5950
rect -4310 5930 -4290 5950
rect -4270 5930 -4250 5950
rect -4230 5930 -4210 5950
rect -4190 5930 -4170 5950
rect -4150 5930 -4130 5950
rect -4110 5930 -4090 5950
rect -4070 5930 -4050 5950
rect -4030 5930 -4010 5950
rect -3990 5930 -3970 5950
rect -3950 5930 -3930 5950
rect -3910 5930 -3890 5950
rect -3870 5930 -3850 5950
rect -3830 5930 -3810 5950
rect -3790 5930 -3770 5950
rect -3750 5930 -3730 5950
rect -3710 5930 -3690 5950
rect -3670 5930 -3660 5950
rect -4460 5760 -3660 5930
rect -4460 5740 -4450 5760
rect -4430 5740 -4410 5760
rect -4390 5740 -4370 5760
rect -4350 5740 -4330 5760
rect -4310 5740 -4290 5760
rect -4270 5740 -4250 5760
rect -4230 5740 -4210 5760
rect -4190 5740 -4170 5760
rect -4150 5740 -4130 5760
rect -4110 5740 -4090 5760
rect -4070 5740 -4050 5760
rect -4030 5740 -4010 5760
rect -3990 5740 -3970 5760
rect -3950 5740 -3930 5760
rect -3910 5740 -3890 5760
rect -3870 5740 -3850 5760
rect -3830 5740 -3810 5760
rect -3790 5740 -3770 5760
rect -3750 5740 -3730 5760
rect -3710 5740 -3690 5760
rect -3670 5740 -3660 5760
rect -4460 5570 -3660 5740
rect -4460 5550 -4450 5570
rect -4430 5550 -4410 5570
rect -4390 5550 -4370 5570
rect -4350 5550 -4330 5570
rect -4310 5550 -4290 5570
rect -4270 5550 -4250 5570
rect -4230 5550 -4210 5570
rect -4190 5550 -4170 5570
rect -4150 5550 -4130 5570
rect -4110 5550 -4090 5570
rect -4070 5550 -4050 5570
rect -4030 5550 -4010 5570
rect -3990 5550 -3970 5570
rect -3950 5550 -3930 5570
rect -3910 5550 -3890 5570
rect -3870 5550 -3850 5570
rect -3830 5550 -3810 5570
rect -3790 5550 -3770 5570
rect -3750 5550 -3730 5570
rect -3710 5550 -3690 5570
rect -3670 5550 -3660 5570
rect -4460 5380 -3660 5550
rect -4460 5360 -4450 5380
rect -4430 5360 -4410 5380
rect -4390 5360 -4370 5380
rect -4350 5360 -4330 5380
rect -4310 5360 -4290 5380
rect -4270 5360 -4250 5380
rect -4230 5360 -4210 5380
rect -4190 5360 -4170 5380
rect -4150 5360 -4130 5380
rect -4110 5360 -4090 5380
rect -4070 5360 -4050 5380
rect -4030 5360 -4010 5380
rect -3990 5360 -3970 5380
rect -3950 5360 -3930 5380
rect -3910 5360 -3890 5380
rect -3870 5360 -3850 5380
rect -3830 5360 -3810 5380
rect -3790 5360 -3770 5380
rect -3750 5360 -3730 5380
rect -3710 5360 -3690 5380
rect -3670 5360 -3660 5380
rect -4460 5190 -3660 5360
rect -4460 5170 -4450 5190
rect -4430 5170 -4410 5190
rect -4390 5170 -4370 5190
rect -4350 5170 -4330 5190
rect -4310 5170 -4290 5190
rect -4270 5170 -4250 5190
rect -4230 5170 -4210 5190
rect -4190 5170 -4170 5190
rect -4150 5170 -4130 5190
rect -4110 5170 -4090 5190
rect -4070 5170 -4050 5190
rect -4030 5170 -4010 5190
rect -3990 5170 -3970 5190
rect -3950 5170 -3930 5190
rect -3910 5170 -3890 5190
rect -3870 5170 -3850 5190
rect -3830 5170 -3810 5190
rect -3790 5170 -3770 5190
rect -3750 5170 -3730 5190
rect -3710 5170 -3690 5190
rect -3670 5170 -3660 5190
rect -4460 5000 -3660 5170
rect -4460 4980 -4450 5000
rect -4430 4980 -4410 5000
rect -4390 4980 -4370 5000
rect -4350 4980 -4330 5000
rect -4310 4980 -4290 5000
rect -4270 4980 -4250 5000
rect -4230 4980 -4210 5000
rect -4190 4980 -4170 5000
rect -4150 4980 -4130 5000
rect -4110 4980 -4090 5000
rect -4070 4980 -4050 5000
rect -4030 4980 -4010 5000
rect -3990 4980 -3970 5000
rect -3950 4980 -3930 5000
rect -3910 4980 -3890 5000
rect -3870 4980 -3850 5000
rect -3830 4980 -3810 5000
rect -3790 4980 -3770 5000
rect -3750 4980 -3730 5000
rect -3710 4980 -3690 5000
rect -3670 4980 -3660 5000
rect -4460 4810 -3660 4980
rect -4460 4790 -4450 4810
rect -4430 4790 -4410 4810
rect -4390 4790 -4370 4810
rect -4350 4790 -4330 4810
rect -4310 4790 -4290 4810
rect -4270 4790 -4250 4810
rect -4230 4790 -4210 4810
rect -4190 4790 -4170 4810
rect -4150 4790 -4130 4810
rect -4110 4790 -4090 4810
rect -4070 4790 -4050 4810
rect -4030 4790 -4010 4810
rect -3990 4790 -3970 4810
rect -3950 4790 -3930 4810
rect -3910 4790 -3890 4810
rect -3870 4790 -3850 4810
rect -3830 4790 -3810 4810
rect -3790 4790 -3770 4810
rect -3750 4790 -3730 4810
rect -3710 4790 -3690 4810
rect -3670 4790 -3660 4810
rect -4460 4620 -3660 4790
rect -4460 4600 -4450 4620
rect -4430 4600 -4410 4620
rect -4390 4600 -4370 4620
rect -4350 4600 -4330 4620
rect -4310 4600 -4290 4620
rect -4270 4600 -4250 4620
rect -4230 4600 -4210 4620
rect -4190 4600 -4170 4620
rect -4150 4600 -4130 4620
rect -4110 4600 -4090 4620
rect -4070 4600 -4050 4620
rect -4030 4600 -4010 4620
rect -3990 4600 -3970 4620
rect -3950 4600 -3930 4620
rect -3910 4600 -3890 4620
rect -3870 4600 -3850 4620
rect -3830 4600 -3810 4620
rect -3790 4600 -3770 4620
rect -3750 4600 -3730 4620
rect -3710 4600 -3690 4620
rect -3670 4600 -3660 4620
rect -4460 4430 -3660 4600
rect -4460 4410 -4450 4430
rect -4430 4410 -4410 4430
rect -4390 4410 -4370 4430
rect -4350 4410 -4330 4430
rect -4310 4410 -4290 4430
rect -4270 4410 -4250 4430
rect -4230 4410 -4210 4430
rect -4190 4410 -4170 4430
rect -4150 4410 -4130 4430
rect -4110 4410 -4090 4430
rect -4070 4410 -4050 4430
rect -4030 4410 -4010 4430
rect -3990 4410 -3970 4430
rect -3950 4410 -3930 4430
rect -3910 4410 -3890 4430
rect -3870 4410 -3850 4430
rect -3830 4410 -3810 4430
rect -3790 4410 -3770 4430
rect -3750 4410 -3730 4430
rect -3710 4410 -3690 4430
rect -3670 4410 -3660 4430
rect -4460 4240 -3660 4410
rect -4460 4220 -4450 4240
rect -4430 4220 -4410 4240
rect -4390 4220 -4370 4240
rect -4350 4220 -4330 4240
rect -4310 4220 -4290 4240
rect -4270 4220 -4250 4240
rect -4230 4220 -4210 4240
rect -4190 4220 -4170 4240
rect -4150 4220 -4130 4240
rect -4110 4220 -4090 4240
rect -4070 4220 -4050 4240
rect -4030 4220 -4010 4240
rect -3990 4220 -3970 4240
rect -3950 4220 -3930 4240
rect -3910 4220 -3890 4240
rect -3870 4220 -3850 4240
rect -3830 4220 -3810 4240
rect -3790 4220 -3770 4240
rect -3750 4220 -3730 4240
rect -3710 4220 -3690 4240
rect -3670 4220 -3660 4240
rect -4460 4050 -3660 4220
rect -4460 4030 -4450 4050
rect -4430 4030 -4410 4050
rect -4390 4030 -4370 4050
rect -4350 4030 -4330 4050
rect -4310 4030 -4290 4050
rect -4270 4030 -4250 4050
rect -4230 4030 -4210 4050
rect -4190 4030 -4170 4050
rect -4150 4030 -4130 4050
rect -4110 4030 -4090 4050
rect -4070 4030 -4050 4050
rect -4030 4030 -4010 4050
rect -3990 4030 -3970 4050
rect -3950 4030 -3930 4050
rect -3910 4030 -3890 4050
rect -3870 4030 -3850 4050
rect -3830 4030 -3810 4050
rect -3790 4030 -3770 4050
rect -3750 4030 -3730 4050
rect -3710 4030 -3690 4050
rect -3670 4030 -3660 4050
rect -4460 3860 -3660 4030
rect -4460 3840 -4450 3860
rect -4430 3840 -4410 3860
rect -4390 3840 -4370 3860
rect -4350 3840 -4330 3860
rect -4310 3840 -4290 3860
rect -4270 3840 -4250 3860
rect -4230 3840 -4210 3860
rect -4190 3840 -4170 3860
rect -4150 3840 -4130 3860
rect -4110 3840 -4090 3860
rect -4070 3840 -4050 3860
rect -4030 3840 -4010 3860
rect -3990 3840 -3970 3860
rect -3950 3840 -3930 3860
rect -3910 3840 -3890 3860
rect -3870 3840 -3850 3860
rect -3830 3840 -3810 3860
rect -3790 3840 -3770 3860
rect -3750 3840 -3730 3860
rect -3710 3840 -3690 3860
rect -3670 3840 -3660 3860
rect -4460 3670 -3660 3840
rect -4460 3650 -4450 3670
rect -4430 3650 -4410 3670
rect -4390 3650 -4370 3670
rect -4350 3650 -4330 3670
rect -4310 3650 -4290 3670
rect -4270 3650 -4250 3670
rect -4230 3650 -4210 3670
rect -4190 3650 -4170 3670
rect -4150 3650 -4130 3670
rect -4110 3650 -4090 3670
rect -4070 3650 -4050 3670
rect -4030 3650 -4010 3670
rect -3990 3650 -3970 3670
rect -3950 3650 -3930 3670
rect -3910 3650 -3890 3670
rect -3870 3650 -3850 3670
rect -3830 3650 -3810 3670
rect -3790 3650 -3770 3670
rect -3750 3650 -3730 3670
rect -3710 3650 -3690 3670
rect -3670 3650 -3660 3670
rect -4460 3640 -3660 3650
rect -3075 6010 -2935 6060
rect -3075 6000 -2920 6010
rect -3075 5975 -3070 6000
rect -3050 5975 -3030 6000
rect -3010 5975 -2990 6000
rect -2970 5975 -2950 6000
rect -2930 5975 -2920 6000
rect -3075 5905 -2920 5975
rect -3075 5880 -3070 5905
rect -3050 5880 -3030 5905
rect -3010 5880 -2990 5905
rect -2970 5880 -2950 5905
rect -2930 5880 -2920 5905
rect -3075 5810 -2920 5880
rect -3075 5785 -3070 5810
rect -3050 5785 -3030 5810
rect -3010 5785 -2990 5810
rect -2970 5785 -2950 5810
rect -2930 5785 -2920 5810
rect -3075 5715 -2920 5785
rect -3075 5690 -3070 5715
rect -3050 5690 -3030 5715
rect -3010 5690 -2990 5715
rect -2970 5690 -2950 5715
rect -2930 5690 -2920 5715
rect -3075 5620 -2920 5690
rect -3075 5595 -3070 5620
rect -3050 5595 -3030 5620
rect -3010 5595 -2990 5620
rect -2970 5595 -2950 5620
rect -2930 5595 -2920 5620
rect -3075 5525 -2920 5595
rect -3075 5500 -3070 5525
rect -3050 5500 -3030 5525
rect -3010 5500 -2990 5525
rect -2970 5500 -2950 5525
rect -2930 5500 -2920 5525
rect -3075 5430 -2920 5500
rect -3075 5405 -3070 5430
rect -3050 5405 -3030 5430
rect -3010 5405 -2990 5430
rect -2970 5405 -2950 5430
rect -2930 5405 -2920 5430
rect -3075 5335 -2920 5405
rect -3075 5310 -3070 5335
rect -3050 5310 -3030 5335
rect -3010 5310 -2990 5335
rect -2970 5310 -2950 5335
rect -2930 5310 -2920 5335
rect -3075 5240 -2920 5310
rect -3075 5215 -3070 5240
rect -3050 5215 -3030 5240
rect -3010 5215 -2990 5240
rect -2970 5215 -2950 5240
rect -2930 5215 -2920 5240
rect -3075 5145 -2920 5215
rect -3075 5120 -3070 5145
rect -3050 5120 -3030 5145
rect -3010 5120 -2990 5145
rect -2970 5120 -2950 5145
rect -2930 5120 -2920 5145
rect -3075 5050 -2920 5120
rect -3075 5025 -3070 5050
rect -3050 5025 -3030 5050
rect -3010 5025 -2990 5050
rect -2970 5025 -2950 5050
rect -2930 5025 -2920 5050
rect -3075 4955 -2920 5025
rect -3075 4930 -3070 4955
rect -3050 4930 -3030 4955
rect -3010 4930 -2990 4955
rect -2970 4930 -2950 4955
rect -2930 4930 -2920 4955
rect -3075 4860 -2920 4930
rect -3075 4835 -3070 4860
rect -3050 4835 -3030 4860
rect -3010 4835 -2990 4860
rect -2970 4835 -2950 4860
rect -2930 4835 -2920 4860
rect -3075 4765 -2920 4835
rect -3075 4740 -3070 4765
rect -3050 4740 -3030 4765
rect -3010 4740 -2990 4765
rect -2970 4740 -2950 4765
rect -2930 4740 -2920 4765
rect -3075 4670 -2920 4740
rect -3075 4645 -3070 4670
rect -3050 4645 -3030 4670
rect -3010 4645 -2990 4670
rect -2970 4645 -2950 4670
rect -2930 4645 -2920 4670
rect -3075 4575 -2920 4645
rect -3075 4550 -3070 4575
rect -3050 4550 -3030 4575
rect -3010 4550 -2990 4575
rect -2970 4550 -2950 4575
rect -2930 4550 -2920 4575
rect -3075 4480 -2920 4550
rect -3075 4455 -3070 4480
rect -3050 4455 -3030 4480
rect -3010 4455 -2990 4480
rect -2970 4455 -2950 4480
rect -2930 4455 -2920 4480
rect -3075 4385 -2920 4455
rect -3075 4360 -3070 4385
rect -3050 4360 -3030 4385
rect -3010 4360 -2990 4385
rect -2970 4360 -2950 4385
rect -2930 4360 -2920 4385
rect -3075 4290 -2920 4360
rect -3075 4265 -3070 4290
rect -3050 4265 -3030 4290
rect -3010 4265 -2990 4290
rect -2970 4265 -2950 4290
rect -2930 4265 -2920 4290
rect -3075 4195 -2920 4265
rect -3075 4170 -3070 4195
rect -3050 4170 -3030 4195
rect -3010 4170 -2990 4195
rect -2970 4170 -2950 4195
rect -2930 4170 -2920 4195
rect -3075 4100 -2920 4170
rect -3075 4075 -3070 4100
rect -3050 4075 -3030 4100
rect -3010 4075 -2990 4100
rect -2970 4075 -2950 4100
rect -2930 4075 -2920 4100
rect -3075 4005 -2920 4075
rect -3075 3980 -3070 4005
rect -3050 3980 -3030 4005
rect -3010 3980 -2990 4005
rect -2970 3980 -2950 4005
rect -2930 3980 -2920 4005
rect -3075 3910 -2920 3980
rect -3075 3885 -3070 3910
rect -3050 3885 -3030 3910
rect -3010 3885 -2990 3910
rect -2970 3885 -2950 3910
rect -2930 3885 -2920 3910
rect -3075 3815 -2920 3885
rect -3075 3790 -3070 3815
rect -3050 3790 -3030 3815
rect -3010 3790 -2990 3815
rect -2970 3790 -2950 3815
rect -2930 3790 -2920 3815
rect -3075 3720 -2920 3790
rect -3075 3695 -3070 3720
rect -3050 3695 -3030 3720
rect -3010 3695 -2990 3720
rect -2970 3695 -2950 3720
rect -2930 3695 -2920 3720
rect -3075 3625 -2920 3695
rect -3075 3600 -3070 3625
rect -3050 3600 -3030 3625
rect -3010 3600 -2990 3625
rect -2970 3600 -2950 3625
rect -2930 3600 -2920 3625
rect -3075 3590 -2920 3600
rect -2220 6000 -2065 6060
rect -2220 5975 -2210 6000
rect -2190 5975 -2170 6000
rect -2150 5975 -2130 6000
rect -2110 5975 -2090 6000
rect -2070 5975 -2065 6000
rect -2220 5905 -2065 5975
rect -2220 5880 -2210 5905
rect -2190 5880 -2170 5905
rect -2150 5880 -2130 5905
rect -2110 5880 -2090 5905
rect -2070 5880 -2065 5905
rect -2220 5810 -2065 5880
rect -2220 5785 -2210 5810
rect -2190 5785 -2170 5810
rect -2150 5785 -2130 5810
rect -2110 5785 -2090 5810
rect -2070 5785 -2065 5810
rect -2220 5715 -2065 5785
rect -2220 5690 -2210 5715
rect -2190 5690 -2170 5715
rect -2150 5690 -2130 5715
rect -2110 5690 -2090 5715
rect -2070 5690 -2065 5715
rect -2220 5620 -2065 5690
rect -2220 5595 -2210 5620
rect -2190 5595 -2170 5620
rect -2150 5595 -2130 5620
rect -2110 5595 -2090 5620
rect -2070 5595 -2065 5620
rect -2220 5525 -2065 5595
rect -2220 5500 -2210 5525
rect -2190 5500 -2170 5525
rect -2150 5500 -2130 5525
rect -2110 5500 -2090 5525
rect -2070 5500 -2065 5525
rect -2220 5430 -2065 5500
rect -2220 5405 -2210 5430
rect -2190 5405 -2170 5430
rect -2150 5405 -2130 5430
rect -2110 5405 -2090 5430
rect -2070 5405 -2065 5430
rect -2220 5335 -2065 5405
rect -2220 5310 -2210 5335
rect -2190 5310 -2170 5335
rect -2150 5310 -2130 5335
rect -2110 5310 -2090 5335
rect -2070 5310 -2065 5335
rect -2220 5240 -2065 5310
rect -2220 5215 -2210 5240
rect -2190 5215 -2170 5240
rect -2150 5215 -2130 5240
rect -2110 5215 -2090 5240
rect -2070 5215 -2065 5240
rect -2220 5145 -2065 5215
rect -2220 5120 -2210 5145
rect -2190 5120 -2170 5145
rect -2150 5120 -2130 5145
rect -2110 5120 -2090 5145
rect -2070 5120 -2065 5145
rect -2220 5050 -2065 5120
rect -2220 5025 -2210 5050
rect -2190 5025 -2170 5050
rect -2150 5025 -2130 5050
rect -2110 5025 -2090 5050
rect -2070 5025 -2065 5050
rect -2220 4955 -2065 5025
rect -2220 4930 -2210 4955
rect -2190 4930 -2170 4955
rect -2150 4930 -2130 4955
rect -2110 4930 -2090 4955
rect -2070 4930 -2065 4955
rect -2220 4860 -2065 4930
rect -2220 4835 -2210 4860
rect -2190 4835 -2170 4860
rect -2150 4835 -2130 4860
rect -2110 4835 -2090 4860
rect -2070 4835 -2065 4860
rect -2220 4765 -2065 4835
rect -2220 4740 -2210 4765
rect -2190 4740 -2170 4765
rect -2150 4740 -2130 4765
rect -2110 4740 -2090 4765
rect -2070 4740 -2065 4765
rect -2220 4670 -2065 4740
rect -2220 4645 -2210 4670
rect -2190 4645 -2170 4670
rect -2150 4645 -2130 4670
rect -2110 4645 -2090 4670
rect -2070 4645 -2065 4670
rect -2220 4575 -2065 4645
rect -2220 4550 -2210 4575
rect -2190 4550 -2170 4575
rect -2150 4550 -2130 4575
rect -2110 4550 -2090 4575
rect -2070 4550 -2065 4575
rect -2220 4480 -2065 4550
rect -2220 4455 -2210 4480
rect -2190 4455 -2170 4480
rect -2150 4455 -2130 4480
rect -2110 4455 -2090 4480
rect -2070 4455 -2065 4480
rect -2220 4385 -2065 4455
rect -2220 4360 -2210 4385
rect -2190 4360 -2170 4385
rect -2150 4360 -2130 4385
rect -2110 4360 -2090 4385
rect -2070 4360 -2065 4385
rect -2220 4290 -2065 4360
rect -2220 4265 -2210 4290
rect -2190 4265 -2170 4290
rect -2150 4265 -2130 4290
rect -2110 4265 -2090 4290
rect -2070 4265 -2065 4290
rect -2220 4195 -2065 4265
rect -2220 4170 -2210 4195
rect -2190 4170 -2170 4195
rect -2150 4170 -2130 4195
rect -2110 4170 -2090 4195
rect -2070 4170 -2065 4195
rect -2220 4100 -2065 4170
rect -2220 4075 -2210 4100
rect -2190 4075 -2170 4100
rect -2150 4075 -2130 4100
rect -2110 4075 -2090 4100
rect -2070 4075 -2065 4100
rect -2220 4005 -2065 4075
rect -2220 3980 -2210 4005
rect -2190 3980 -2170 4005
rect -2150 3980 -2130 4005
rect -2110 3980 -2090 4005
rect -2070 3980 -2065 4005
rect -2220 3910 -2065 3980
rect -2220 3885 -2210 3910
rect -2190 3885 -2170 3910
rect -2150 3885 -2130 3910
rect -2110 3885 -2090 3910
rect -2070 3885 -2065 3910
rect -2220 3815 -2065 3885
rect -2220 3790 -2210 3815
rect -2190 3790 -2170 3815
rect -2150 3790 -2130 3815
rect -2110 3790 -2090 3815
rect -2070 3790 -2065 3815
rect -2220 3720 -2065 3790
rect -2220 3695 -2210 3720
rect -2190 3695 -2170 3720
rect -2150 3695 -2130 3720
rect -2110 3695 -2090 3720
rect -2070 3695 -2065 3720
rect -2220 3625 -2065 3695
rect -1480 5950 -680 6285
rect -400 8395 400 8585
rect -400 8375 -390 8395
rect -370 8375 -350 8395
rect -330 8375 -310 8395
rect -290 8375 -270 8395
rect -250 8375 -230 8395
rect -210 8375 -190 8395
rect -170 8375 -150 8395
rect -130 8375 -110 8395
rect -90 8375 -70 8395
rect -50 8375 -30 8395
rect -10 8375 10 8395
rect 30 8375 50 8395
rect 70 8375 90 8395
rect 110 8375 130 8395
rect 150 8375 170 8395
rect 190 8375 210 8395
rect 230 8375 250 8395
rect 270 8375 290 8395
rect 310 8375 330 8395
rect 350 8375 370 8395
rect 390 8375 400 8395
rect -400 8231 400 8375
rect -400 8211 -390 8231
rect -370 8211 -350 8231
rect -330 8211 -310 8231
rect -290 8211 -270 8231
rect -250 8211 -230 8231
rect -210 8211 -190 8231
rect -170 8211 -150 8231
rect -130 8211 -110 8231
rect -90 8211 -70 8231
rect -50 8211 -30 8231
rect -10 8211 10 8231
rect 30 8211 50 8231
rect 70 8211 90 8231
rect 110 8211 130 8231
rect 150 8211 170 8231
rect 190 8211 210 8231
rect 230 8211 250 8231
rect 270 8211 290 8231
rect 310 8211 330 8231
rect 350 8211 370 8231
rect 390 8211 400 8231
rect -400 8067 400 8211
rect -400 8047 -390 8067
rect -370 8047 -350 8067
rect -330 8047 -310 8067
rect -290 8047 -270 8067
rect -250 8047 -230 8067
rect -210 8047 -190 8067
rect -170 8047 -150 8067
rect -130 8047 -110 8067
rect -90 8047 -70 8067
rect -50 8047 -30 8067
rect -10 8047 10 8067
rect 30 8047 50 8067
rect 70 8047 90 8067
rect 110 8047 130 8067
rect 150 8047 170 8067
rect 190 8047 210 8067
rect 230 8047 250 8067
rect 270 8047 290 8067
rect 310 8047 330 8067
rect 350 8047 370 8067
rect 390 8047 400 8067
rect -400 7903 400 8047
rect -400 7883 -390 7903
rect -370 7883 -350 7903
rect -330 7883 -310 7903
rect -290 7883 -270 7903
rect -250 7883 -230 7903
rect -210 7883 -190 7903
rect -170 7883 -150 7903
rect -130 7883 -110 7903
rect -90 7883 -70 7903
rect -50 7883 -30 7903
rect -10 7883 10 7903
rect 30 7883 50 7903
rect 70 7883 90 7903
rect 110 7883 130 7903
rect 150 7883 170 7903
rect 190 7883 210 7903
rect 230 7883 250 7903
rect 270 7883 290 7903
rect 310 7883 330 7903
rect 350 7883 370 7903
rect 390 7883 400 7903
rect -400 7739 400 7883
rect -400 7719 -390 7739
rect -370 7719 -350 7739
rect -330 7719 -310 7739
rect -290 7719 -270 7739
rect -250 7719 -230 7739
rect -210 7719 -190 7739
rect -170 7719 -150 7739
rect -130 7719 -110 7739
rect -90 7719 -70 7739
rect -50 7719 -30 7739
rect -10 7719 10 7739
rect 30 7719 50 7739
rect 70 7719 90 7739
rect 110 7719 130 7739
rect 150 7719 170 7739
rect 190 7719 210 7739
rect 230 7719 250 7739
rect 270 7719 290 7739
rect 310 7719 330 7739
rect 350 7719 370 7739
rect 390 7719 400 7739
rect -400 7575 400 7719
rect -400 7555 -390 7575
rect -370 7555 -350 7575
rect -330 7555 -310 7575
rect -290 7555 -270 7575
rect -250 7555 -230 7575
rect -210 7555 -190 7575
rect -170 7555 -150 7575
rect -130 7555 -110 7575
rect -90 7555 -70 7575
rect -50 7555 -30 7575
rect -10 7555 10 7575
rect 30 7555 50 7575
rect 70 7555 90 7575
rect 110 7555 130 7575
rect 150 7555 170 7575
rect 190 7555 210 7575
rect 230 7555 250 7575
rect 270 7555 290 7575
rect 310 7555 330 7575
rect 350 7555 370 7575
rect 390 7555 400 7575
rect -400 7411 400 7555
rect -400 7391 -390 7411
rect -370 7391 -350 7411
rect -330 7391 -310 7411
rect -290 7391 -270 7411
rect -250 7391 -230 7411
rect -210 7391 -190 7411
rect -170 7391 -150 7411
rect -130 7391 -110 7411
rect -90 7391 -70 7411
rect -50 7391 -30 7411
rect -10 7391 10 7411
rect 30 7391 50 7411
rect 70 7391 90 7411
rect 110 7391 130 7411
rect 150 7391 170 7411
rect 190 7391 210 7411
rect 230 7391 250 7411
rect 270 7391 290 7411
rect 310 7391 330 7411
rect 350 7391 370 7411
rect 390 7391 400 7411
rect -400 7247 400 7391
rect -400 7227 -390 7247
rect -370 7227 -350 7247
rect -330 7227 -310 7247
rect -290 7227 -270 7247
rect -250 7227 -230 7247
rect -210 7227 -190 7247
rect -170 7227 -150 7247
rect -130 7227 -110 7247
rect -90 7227 -70 7247
rect -50 7227 -30 7247
rect -10 7227 10 7247
rect 30 7227 50 7247
rect 70 7227 90 7247
rect 110 7227 130 7247
rect 150 7227 170 7247
rect 190 7227 210 7247
rect 230 7227 250 7247
rect 270 7227 290 7247
rect 310 7227 330 7247
rect 350 7227 370 7247
rect 390 7227 400 7247
rect -400 7083 400 7227
rect -400 7063 -390 7083
rect -370 7063 -350 7083
rect -330 7063 -310 7083
rect -290 7063 -270 7083
rect -250 7063 -230 7083
rect -210 7063 -190 7083
rect -170 7063 -150 7083
rect -130 7063 -110 7083
rect -90 7063 -70 7083
rect -50 7063 -30 7083
rect -10 7063 10 7083
rect 30 7063 50 7083
rect 70 7063 90 7083
rect 110 7063 130 7083
rect 150 7063 170 7083
rect 190 7063 210 7083
rect 230 7063 250 7083
rect 270 7063 290 7083
rect 310 7063 330 7083
rect 350 7063 370 7083
rect 390 7063 400 7083
rect -400 6919 400 7063
rect -400 6899 -390 6919
rect -370 6899 -350 6919
rect -330 6899 -310 6919
rect -290 6899 -270 6919
rect -250 6899 -230 6919
rect -210 6899 -190 6919
rect -170 6899 -150 6919
rect -130 6899 -110 6919
rect -90 6899 -70 6919
rect -50 6899 -30 6919
rect -10 6899 10 6919
rect 30 6899 50 6919
rect 70 6899 90 6919
rect 110 6899 130 6919
rect 150 6899 170 6919
rect 190 6899 210 6919
rect 230 6899 250 6919
rect 270 6899 290 6919
rect 310 6899 330 6919
rect 350 6899 370 6919
rect 390 6899 400 6919
rect -400 6755 400 6899
rect -400 6735 -390 6755
rect -370 6735 -350 6755
rect -330 6735 -310 6755
rect -290 6735 -270 6755
rect -250 6735 -230 6755
rect -210 6735 -190 6755
rect -170 6735 -150 6755
rect -130 6735 -110 6755
rect -90 6735 -70 6755
rect -50 6735 -30 6755
rect -10 6735 10 6755
rect 30 6735 50 6755
rect 70 6735 90 6755
rect 110 6735 130 6755
rect 150 6735 170 6755
rect 190 6735 210 6755
rect 230 6735 250 6755
rect 270 6735 290 6755
rect 310 6735 330 6755
rect 350 6735 370 6755
rect 390 6735 400 6755
rect -400 6591 400 6735
rect -400 6571 -390 6591
rect -370 6571 -350 6591
rect -330 6571 -310 6591
rect -290 6571 -270 6591
rect -250 6571 -230 6591
rect -210 6571 -190 6591
rect -170 6571 -150 6591
rect -130 6571 -110 6591
rect -90 6571 -70 6591
rect -50 6571 -30 6591
rect -10 6571 10 6591
rect 30 6571 50 6591
rect 70 6571 90 6591
rect 110 6571 130 6591
rect 150 6571 170 6591
rect 190 6571 210 6591
rect 230 6571 250 6591
rect 270 6571 290 6591
rect 310 6571 330 6591
rect 350 6571 370 6591
rect 390 6571 400 6591
rect -400 6427 400 6571
rect -400 6407 -390 6427
rect -370 6407 -350 6427
rect -330 6407 -310 6427
rect -290 6407 -270 6427
rect -250 6407 -230 6427
rect -210 6407 -190 6427
rect -170 6407 -150 6427
rect -130 6407 -110 6427
rect -90 6407 -70 6427
rect -50 6407 -30 6427
rect -10 6407 10 6427
rect 30 6407 50 6427
rect 70 6407 90 6427
rect 110 6407 130 6427
rect 150 6407 170 6427
rect 190 6407 210 6427
rect 230 6407 250 6427
rect 270 6407 290 6427
rect 310 6407 330 6427
rect 350 6407 370 6427
rect 390 6407 400 6427
rect -400 6275 400 6407
rect -1480 5930 -1470 5950
rect -1450 5930 -1430 5950
rect -1410 5930 -1390 5950
rect -1370 5930 -1350 5950
rect -1330 5930 -1310 5950
rect -1290 5930 -1270 5950
rect -1250 5930 -1230 5950
rect -1210 5930 -1190 5950
rect -1170 5930 -1150 5950
rect -1130 5930 -1110 5950
rect -1090 5930 -1070 5950
rect -1050 5930 -1030 5950
rect -1010 5930 -990 5950
rect -970 5930 -950 5950
rect -930 5930 -910 5950
rect -890 5930 -870 5950
rect -850 5930 -830 5950
rect -810 5930 -790 5950
rect -770 5930 -750 5950
rect -730 5930 -710 5950
rect -690 5930 -680 5950
rect -1480 5760 -680 5930
rect -1480 5740 -1470 5760
rect -1450 5740 -1430 5760
rect -1410 5740 -1390 5760
rect -1370 5740 -1350 5760
rect -1330 5740 -1310 5760
rect -1290 5740 -1270 5760
rect -1250 5740 -1230 5760
rect -1210 5740 -1190 5760
rect -1170 5740 -1150 5760
rect -1130 5740 -1110 5760
rect -1090 5740 -1070 5760
rect -1050 5740 -1030 5760
rect -1010 5740 -990 5760
rect -970 5740 -950 5760
rect -930 5740 -910 5760
rect -890 5740 -870 5760
rect -850 5740 -830 5760
rect -810 5740 -790 5760
rect -770 5740 -750 5760
rect -730 5740 -710 5760
rect -690 5740 -680 5760
rect -1480 5570 -680 5740
rect -1480 5550 -1470 5570
rect -1450 5550 -1430 5570
rect -1410 5550 -1390 5570
rect -1370 5550 -1350 5570
rect -1330 5550 -1310 5570
rect -1290 5550 -1270 5570
rect -1250 5550 -1230 5570
rect -1210 5550 -1190 5570
rect -1170 5550 -1150 5570
rect -1130 5550 -1110 5570
rect -1090 5550 -1070 5570
rect -1050 5550 -1030 5570
rect -1010 5550 -990 5570
rect -970 5550 -950 5570
rect -930 5550 -910 5570
rect -890 5550 -870 5570
rect -850 5550 -830 5570
rect -810 5550 -790 5570
rect -770 5550 -750 5570
rect -730 5550 -710 5570
rect -690 5550 -680 5570
rect -1480 5380 -680 5550
rect -1480 5360 -1470 5380
rect -1450 5360 -1430 5380
rect -1410 5360 -1390 5380
rect -1370 5360 -1350 5380
rect -1330 5360 -1310 5380
rect -1290 5360 -1270 5380
rect -1250 5360 -1230 5380
rect -1210 5360 -1190 5380
rect -1170 5360 -1150 5380
rect -1130 5360 -1110 5380
rect -1090 5360 -1070 5380
rect -1050 5360 -1030 5380
rect -1010 5360 -990 5380
rect -970 5360 -950 5380
rect -930 5360 -910 5380
rect -890 5360 -870 5380
rect -850 5360 -830 5380
rect -810 5360 -790 5380
rect -770 5360 -750 5380
rect -730 5360 -710 5380
rect -690 5360 -680 5380
rect -1480 5190 -680 5360
rect -1480 5170 -1470 5190
rect -1450 5170 -1430 5190
rect -1410 5170 -1390 5190
rect -1370 5170 -1350 5190
rect -1330 5170 -1310 5190
rect -1290 5170 -1270 5190
rect -1250 5170 -1230 5190
rect -1210 5170 -1190 5190
rect -1170 5170 -1150 5190
rect -1130 5170 -1110 5190
rect -1090 5170 -1070 5190
rect -1050 5170 -1030 5190
rect -1010 5170 -990 5190
rect -970 5170 -950 5190
rect -930 5170 -910 5190
rect -890 5170 -870 5190
rect -850 5170 -830 5190
rect -810 5170 -790 5190
rect -770 5170 -750 5190
rect -730 5170 -710 5190
rect -690 5170 -680 5190
rect -1480 5000 -680 5170
rect -1480 4980 -1470 5000
rect -1450 4980 -1430 5000
rect -1410 4980 -1390 5000
rect -1370 4980 -1350 5000
rect -1330 4980 -1310 5000
rect -1290 4980 -1270 5000
rect -1250 4980 -1230 5000
rect -1210 4980 -1190 5000
rect -1170 4980 -1150 5000
rect -1130 4980 -1110 5000
rect -1090 4980 -1070 5000
rect -1050 4980 -1030 5000
rect -1010 4980 -990 5000
rect -970 4980 -950 5000
rect -930 4980 -910 5000
rect -890 4980 -870 5000
rect -850 4980 -830 5000
rect -810 4980 -790 5000
rect -770 4980 -750 5000
rect -730 4980 -710 5000
rect -690 4980 -680 5000
rect -1480 4810 -680 4980
rect -1480 4790 -1470 4810
rect -1450 4790 -1430 4810
rect -1410 4790 -1390 4810
rect -1370 4790 -1350 4810
rect -1330 4790 -1310 4810
rect -1290 4790 -1270 4810
rect -1250 4790 -1230 4810
rect -1210 4790 -1190 4810
rect -1170 4790 -1150 4810
rect -1130 4790 -1110 4810
rect -1090 4790 -1070 4810
rect -1050 4790 -1030 4810
rect -1010 4790 -990 4810
rect -970 4790 -950 4810
rect -930 4790 -910 4810
rect -890 4790 -870 4810
rect -850 4790 -830 4810
rect -810 4790 -790 4810
rect -770 4790 -750 4810
rect -730 4790 -710 4810
rect -690 4790 -680 4810
rect -1480 4620 -680 4790
rect -1480 4600 -1470 4620
rect -1450 4600 -1430 4620
rect -1410 4600 -1390 4620
rect -1370 4600 -1350 4620
rect -1330 4600 -1310 4620
rect -1290 4600 -1270 4620
rect -1250 4600 -1230 4620
rect -1210 4600 -1190 4620
rect -1170 4600 -1150 4620
rect -1130 4600 -1110 4620
rect -1090 4600 -1070 4620
rect -1050 4600 -1030 4620
rect -1010 4600 -990 4620
rect -970 4600 -950 4620
rect -930 4600 -910 4620
rect -890 4600 -870 4620
rect -850 4600 -830 4620
rect -810 4600 -790 4620
rect -770 4600 -750 4620
rect -730 4600 -710 4620
rect -690 4600 -680 4620
rect -1480 4430 -680 4600
rect -1480 4410 -1470 4430
rect -1450 4410 -1430 4430
rect -1410 4410 -1390 4430
rect -1370 4410 -1350 4430
rect -1330 4410 -1310 4430
rect -1290 4410 -1270 4430
rect -1250 4410 -1230 4430
rect -1210 4410 -1190 4430
rect -1170 4410 -1150 4430
rect -1130 4410 -1110 4430
rect -1090 4410 -1070 4430
rect -1050 4410 -1030 4430
rect -1010 4410 -990 4430
rect -970 4410 -950 4430
rect -930 4410 -910 4430
rect -890 4410 -870 4430
rect -850 4410 -830 4430
rect -810 4410 -790 4430
rect -770 4410 -750 4430
rect -730 4410 -710 4430
rect -690 4410 -680 4430
rect -1480 4240 -680 4410
rect -1480 4220 -1470 4240
rect -1450 4220 -1430 4240
rect -1410 4220 -1390 4240
rect -1370 4220 -1350 4240
rect -1330 4220 -1310 4240
rect -1290 4220 -1270 4240
rect -1250 4220 -1230 4240
rect -1210 4220 -1190 4240
rect -1170 4220 -1150 4240
rect -1130 4220 -1110 4240
rect -1090 4220 -1070 4240
rect -1050 4220 -1030 4240
rect -1010 4220 -990 4240
rect -970 4220 -950 4240
rect -930 4220 -910 4240
rect -890 4220 -870 4240
rect -850 4220 -830 4240
rect -810 4220 -790 4240
rect -770 4220 -750 4240
rect -730 4220 -710 4240
rect -690 4220 -680 4240
rect -1480 4050 -680 4220
rect -1480 4030 -1470 4050
rect -1450 4030 -1430 4050
rect -1410 4030 -1390 4050
rect -1370 4030 -1350 4050
rect -1330 4030 -1310 4050
rect -1290 4030 -1270 4050
rect -1250 4030 -1230 4050
rect -1210 4030 -1190 4050
rect -1170 4030 -1150 4050
rect -1130 4030 -1110 4050
rect -1090 4030 -1070 4050
rect -1050 4030 -1030 4050
rect -1010 4030 -990 4050
rect -970 4030 -950 4050
rect -930 4030 -910 4050
rect -890 4030 -870 4050
rect -850 4030 -830 4050
rect -810 4030 -790 4050
rect -770 4030 -750 4050
rect -730 4030 -710 4050
rect -690 4030 -680 4050
rect -1480 3860 -680 4030
rect -1480 3840 -1470 3860
rect -1450 3840 -1430 3860
rect -1410 3840 -1390 3860
rect -1370 3840 -1350 3860
rect -1330 3840 -1310 3860
rect -1290 3840 -1270 3860
rect -1250 3840 -1230 3860
rect -1210 3840 -1190 3860
rect -1170 3840 -1150 3860
rect -1130 3840 -1110 3860
rect -1090 3840 -1070 3860
rect -1050 3840 -1030 3860
rect -1010 3840 -990 3860
rect -970 3840 -950 3860
rect -930 3840 -910 3860
rect -890 3840 -870 3860
rect -850 3840 -830 3860
rect -810 3840 -790 3860
rect -770 3840 -750 3860
rect -730 3840 -710 3860
rect -690 3840 -680 3860
rect -1480 3670 -680 3840
rect -1480 3650 -1470 3670
rect -1450 3650 -1430 3670
rect -1410 3650 -1390 3670
rect -1370 3650 -1350 3670
rect -1330 3650 -1310 3670
rect -1290 3650 -1270 3670
rect -1250 3650 -1230 3670
rect -1210 3650 -1190 3670
rect -1170 3650 -1150 3670
rect -1130 3650 -1110 3670
rect -1090 3650 -1070 3670
rect -1050 3650 -1030 3670
rect -1010 3650 -990 3670
rect -970 3650 -950 3670
rect -930 3650 -910 3670
rect -890 3650 -870 3670
rect -850 3650 -830 3670
rect -810 3650 -790 3670
rect -770 3650 -750 3670
rect -730 3650 -710 3670
rect -690 3650 -680 3670
rect -1480 3640 -680 3650
rect -400 6085 400 6095
rect -400 6065 -390 6085
rect -370 6065 -350 6085
rect -330 6065 -310 6085
rect -290 6065 -270 6085
rect -250 6065 -230 6085
rect -210 6065 -190 6085
rect -170 6065 -150 6085
rect -130 6065 -110 6085
rect -90 6065 -70 6085
rect -50 6065 -30 6085
rect -10 6065 10 6085
rect 30 6065 50 6085
rect 70 6065 90 6085
rect 110 6065 130 6085
rect 150 6065 170 6085
rect 190 6065 210 6085
rect 230 6065 250 6085
rect 270 6065 290 6085
rect 310 6065 330 6085
rect 350 6065 370 6085
rect 390 6065 400 6085
rect -400 6045 400 6065
rect -400 6025 -390 6045
rect -370 6025 -350 6045
rect -330 6025 -310 6045
rect -290 6025 -270 6045
rect -250 6025 -230 6045
rect -210 6025 -190 6045
rect -170 6025 -150 6045
rect -130 6025 -110 6045
rect -90 6025 -70 6045
rect -50 6025 -30 6045
rect -10 6025 10 6045
rect 30 6025 50 6045
rect 70 6025 90 6045
rect 110 6025 130 6045
rect 150 6025 170 6045
rect 190 6025 210 6045
rect 230 6025 250 6045
rect 270 6025 290 6045
rect 310 6025 330 6045
rect 350 6025 370 6045
rect 390 6025 400 6045
rect -400 5855 400 6025
rect -400 5835 -390 5855
rect -370 5835 -350 5855
rect -330 5835 -310 5855
rect -290 5835 -270 5855
rect -250 5835 -230 5855
rect -210 5835 -190 5855
rect -170 5835 -150 5855
rect -130 5835 -110 5855
rect -90 5835 -70 5855
rect -50 5835 -30 5855
rect -10 5835 10 5855
rect 30 5835 50 5855
rect 70 5835 90 5855
rect 110 5835 130 5855
rect 150 5835 170 5855
rect 190 5835 210 5855
rect 230 5835 250 5855
rect 270 5835 290 5855
rect 310 5835 330 5855
rect 350 5835 370 5855
rect 390 5835 400 5855
rect -400 5665 400 5835
rect -400 5645 -390 5665
rect -370 5645 -350 5665
rect -330 5645 -310 5665
rect -290 5645 -270 5665
rect -250 5645 -230 5665
rect -210 5645 -190 5665
rect -170 5645 -150 5665
rect -130 5645 -110 5665
rect -90 5645 -70 5665
rect -50 5645 -30 5665
rect -10 5645 10 5665
rect 30 5645 50 5665
rect 70 5645 90 5665
rect 110 5645 130 5665
rect 150 5645 170 5665
rect 190 5645 210 5665
rect 230 5645 250 5665
rect 270 5645 290 5665
rect 310 5645 330 5665
rect 350 5645 370 5665
rect 390 5645 400 5665
rect -400 5475 400 5645
rect -400 5455 -390 5475
rect -370 5455 -350 5475
rect -330 5455 -310 5475
rect -290 5455 -270 5475
rect -250 5455 -230 5475
rect -210 5455 -190 5475
rect -170 5455 -150 5475
rect -130 5455 -110 5475
rect -90 5455 -70 5475
rect -50 5455 -30 5475
rect -10 5455 10 5475
rect 30 5455 50 5475
rect 70 5455 90 5475
rect 110 5455 130 5475
rect 150 5455 170 5475
rect 190 5455 210 5475
rect 230 5455 250 5475
rect 270 5455 290 5475
rect 310 5455 330 5475
rect 350 5455 370 5475
rect 390 5455 400 5475
rect -400 5285 400 5455
rect -400 5265 -390 5285
rect -370 5265 -350 5285
rect -330 5265 -310 5285
rect -290 5265 -270 5285
rect -250 5265 -230 5285
rect -210 5265 -190 5285
rect -170 5265 -150 5285
rect -130 5265 -110 5285
rect -90 5265 -70 5285
rect -50 5265 -30 5285
rect -10 5265 10 5285
rect 30 5265 50 5285
rect 70 5265 90 5285
rect 110 5265 130 5285
rect 150 5265 170 5285
rect 190 5265 210 5285
rect 230 5265 250 5285
rect 270 5265 290 5285
rect 310 5265 330 5285
rect 350 5265 370 5285
rect 390 5265 400 5285
rect -400 5095 400 5265
rect -400 5075 -390 5095
rect -370 5075 -350 5095
rect -330 5075 -310 5095
rect -290 5075 -270 5095
rect -250 5075 -230 5095
rect -210 5075 -190 5095
rect -170 5075 -150 5095
rect -130 5075 -110 5095
rect -90 5075 -70 5095
rect -50 5075 -30 5095
rect -10 5075 10 5095
rect 30 5075 50 5095
rect 70 5075 90 5095
rect 110 5075 130 5095
rect 150 5075 170 5095
rect 190 5075 210 5095
rect 230 5075 250 5095
rect 270 5075 290 5095
rect 310 5075 330 5095
rect 350 5075 370 5095
rect 390 5075 400 5095
rect -400 4905 400 5075
rect -400 4885 -390 4905
rect -370 4885 -350 4905
rect -330 4885 -310 4905
rect -290 4885 -270 4905
rect -250 4885 -230 4905
rect -210 4885 -190 4905
rect -170 4885 -150 4905
rect -130 4885 -110 4905
rect -90 4885 -70 4905
rect -50 4885 -30 4905
rect -10 4885 10 4905
rect 30 4885 50 4905
rect 70 4885 90 4905
rect 110 4885 130 4905
rect 150 4885 170 4905
rect 190 4885 210 4905
rect 230 4885 250 4905
rect 270 4885 290 4905
rect 310 4885 330 4905
rect 350 4885 370 4905
rect 390 4885 400 4905
rect -400 4715 400 4885
rect -400 4695 -390 4715
rect -370 4695 -350 4715
rect -330 4695 -310 4715
rect -290 4695 -270 4715
rect -250 4695 -230 4715
rect -210 4695 -190 4715
rect -170 4695 -150 4715
rect -130 4695 -110 4715
rect -90 4695 -70 4715
rect -50 4695 -30 4715
rect -10 4695 10 4715
rect 30 4695 50 4715
rect 70 4695 90 4715
rect 110 4695 130 4715
rect 150 4695 170 4715
rect 190 4695 210 4715
rect 230 4695 250 4715
rect 270 4695 290 4715
rect 310 4695 330 4715
rect 350 4695 370 4715
rect 390 4695 400 4715
rect -400 4525 400 4695
rect -400 4505 -390 4525
rect -370 4505 -350 4525
rect -330 4505 -310 4525
rect -290 4505 -270 4525
rect -250 4505 -230 4525
rect -210 4505 -190 4525
rect -170 4505 -150 4525
rect -130 4505 -110 4525
rect -90 4505 -70 4525
rect -50 4505 -30 4525
rect -10 4505 10 4525
rect 30 4505 50 4525
rect 70 4505 90 4525
rect 110 4505 130 4525
rect 150 4505 170 4525
rect 190 4505 210 4525
rect 230 4505 250 4525
rect 270 4505 290 4525
rect 310 4505 330 4525
rect 350 4505 370 4525
rect 390 4505 400 4525
rect -400 4335 400 4505
rect -400 4315 -390 4335
rect -370 4315 -350 4335
rect -330 4315 -310 4335
rect -290 4315 -270 4335
rect -250 4315 -230 4335
rect -210 4315 -190 4335
rect -170 4315 -150 4335
rect -130 4315 -110 4335
rect -90 4315 -70 4335
rect -50 4315 -30 4335
rect -10 4315 10 4335
rect 30 4315 50 4335
rect 70 4315 90 4335
rect 110 4315 130 4335
rect 150 4315 170 4335
rect 190 4315 210 4335
rect 230 4315 250 4335
rect 270 4315 290 4335
rect 310 4315 330 4335
rect 350 4315 370 4335
rect 390 4315 400 4335
rect -400 4145 400 4315
rect -400 4125 -390 4145
rect -370 4125 -350 4145
rect -330 4125 -310 4145
rect -290 4125 -270 4145
rect -250 4125 -230 4145
rect -210 4125 -190 4145
rect -170 4125 -150 4145
rect -130 4125 -110 4145
rect -90 4125 -70 4145
rect -50 4125 -30 4145
rect -10 4125 10 4145
rect 30 4125 50 4145
rect 70 4125 90 4145
rect 110 4125 130 4145
rect 150 4125 170 4145
rect 190 4125 210 4145
rect 230 4125 250 4145
rect 270 4125 290 4145
rect 310 4125 330 4145
rect 350 4125 370 4145
rect 390 4125 400 4145
rect -400 3955 400 4125
rect -400 3935 -390 3955
rect -370 3935 -350 3955
rect -330 3935 -310 3955
rect -290 3935 -270 3955
rect -250 3935 -230 3955
rect -210 3935 -190 3955
rect -170 3935 -150 3955
rect -130 3935 -110 3955
rect -90 3935 -70 3955
rect -50 3935 -30 3955
rect -10 3935 10 3955
rect 30 3935 50 3955
rect 70 3935 90 3955
rect 110 3935 130 3955
rect 150 3935 170 3955
rect 190 3935 210 3955
rect 230 3935 250 3955
rect 270 3935 290 3955
rect 310 3935 330 3955
rect 350 3935 370 3955
rect 390 3935 400 3955
rect -400 3765 400 3935
rect -400 3745 -390 3765
rect -370 3745 -350 3765
rect -330 3745 -310 3765
rect -290 3745 -270 3765
rect -250 3745 -230 3765
rect -210 3745 -190 3765
rect -170 3745 -150 3765
rect -130 3745 -110 3765
rect -90 3745 -70 3765
rect -50 3745 -30 3765
rect -10 3745 10 3765
rect 30 3745 50 3765
rect 70 3745 90 3765
rect 110 3745 130 3765
rect 150 3745 170 3765
rect 190 3745 210 3765
rect 230 3745 250 3765
rect 270 3745 290 3765
rect 310 3745 330 3765
rect 350 3745 370 3765
rect 390 3745 400 3765
rect -2220 3600 -2210 3625
rect -2190 3600 -2170 3625
rect -2150 3600 -2130 3625
rect -2110 3600 -2090 3625
rect -2070 3600 -2065 3625
rect -2220 3590 -2065 3600
rect -5540 3555 -5530 3575
rect -5510 3555 -5490 3575
rect -5470 3555 -5450 3575
rect -5430 3555 -5410 3575
rect -5390 3555 -5370 3575
rect -5350 3555 -5330 3575
rect -5310 3555 -5290 3575
rect -5270 3555 -5250 3575
rect -5230 3555 -5210 3575
rect -5190 3555 -5170 3575
rect -5150 3555 -5130 3575
rect -5110 3555 -5090 3575
rect -5070 3555 -5050 3575
rect -5030 3555 -5010 3575
rect -4990 3555 -4970 3575
rect -4950 3555 -4930 3575
rect -4910 3555 -4890 3575
rect -4870 3555 -4850 3575
rect -4830 3555 -4810 3575
rect -4790 3555 -4770 3575
rect -4750 3555 -4740 3575
rect -5540 3535 -4740 3555
rect -5540 3515 -5530 3535
rect -5510 3515 -5490 3535
rect -5470 3515 -5450 3535
rect -5430 3515 -5410 3535
rect -5390 3515 -5370 3535
rect -5350 3515 -5330 3535
rect -5310 3515 -5290 3535
rect -5270 3515 -5250 3535
rect -5230 3515 -5210 3535
rect -5190 3515 -5170 3535
rect -5150 3515 -5130 3535
rect -5110 3515 -5090 3535
rect -5070 3515 -5050 3535
rect -5030 3515 -5010 3535
rect -4990 3515 -4970 3535
rect -4950 3515 -4930 3535
rect -4910 3515 -4890 3535
rect -4870 3515 -4850 3535
rect -4830 3515 -4810 3535
rect -4790 3515 -4770 3535
rect -4750 3515 -4740 3535
rect -5540 3500 -4740 3515
rect -400 3575 400 3745
rect -400 3555 -390 3575
rect -370 3555 -350 3575
rect -330 3555 -310 3575
rect -290 3555 -270 3575
rect -250 3555 -230 3575
rect -210 3555 -190 3575
rect -170 3555 -150 3575
rect -130 3555 -110 3575
rect -90 3555 -70 3575
rect -50 3555 -30 3575
rect -10 3555 10 3575
rect 30 3555 50 3575
rect 70 3555 90 3575
rect 110 3555 130 3575
rect 150 3555 170 3575
rect 190 3555 210 3575
rect 230 3555 250 3575
rect 270 3555 290 3575
rect 310 3555 330 3575
rect 350 3555 370 3575
rect 390 3555 400 3575
rect -400 3535 400 3555
rect -400 3515 -390 3535
rect -370 3515 -350 3535
rect -330 3515 -310 3535
rect -290 3515 -270 3535
rect -250 3515 -230 3535
rect -210 3515 -190 3535
rect -170 3515 -150 3535
rect -130 3515 -110 3535
rect -90 3515 -70 3535
rect -50 3515 -30 3535
rect -10 3515 10 3535
rect 30 3515 50 3535
rect 70 3515 90 3535
rect 110 3515 130 3535
rect 150 3515 170 3535
rect 190 3515 210 3535
rect 230 3515 250 3535
rect 270 3515 290 3535
rect 310 3515 330 3535
rect 350 3515 370 3535
rect 390 3515 400 3535
rect -400 3500 400 3515
<< labels >>
rlabel metal1 20 3645 20 3645 1 GND
port 9 n
rlabel metal1 -1075 6275 -1075 6275 1 Vout_p
port 5 n
rlabel metal1 -5140 8635 -5140 8635 1 VDD
port 2 n
rlabel metal1 -4075 6275 -4075 6275 1 Vout_n
port 6 n
rlabel metal1 -3005 7425 -3005 7425 1 Vin_n
port 3 n
rlabel metal1 -5135 3650 -5135 3650 1 GND
port 9 n
rlabel metal1 85 8640 85 8640 1 VDD
port 9 n
rlabel metal1 -2935 4805 -2935 4805 1 Vb4
port 10 n
rlabel metal1 -2210 4805 -2210 4805 1 Vb4
port 10 n
rlabel metal1 -2135 7415 -2135 7415 1 Vin_p
port 11 n
<< end >>
