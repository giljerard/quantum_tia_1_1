magic
tech sky130A
timestamp 1640986451
<< metal1 >>
rect -5540 8475 -4740 8650
rect -400 8475 400 8650
rect -3155 7395 -2990 7455
rect -2150 7395 -1985 7455
rect -4460 6170 -3660 6310
rect -1480 6170 -680 6310
rect -3075 6010 -2920 6060
rect -3075 5700 -2935 6010
rect -3075 5595 -2920 5700
rect -3075 3815 -2935 5595
rect -2220 3815 -2065 6060
rect -5540 3630 -4740 3680
rect -400 3630 400 3680
use sf_half  sf_half_1
timestamp 1640983407
transform -1 0 -2990 0 1 6260
box -145 -2760 2855 2430
use sf_half  sf_half_0
timestamp 1640983407
transform 1 0 -2150 0 1 6260
box -145 -2760 2855 2430
<< labels >>
rlabel metal1 20 3645 20 3645 1 GND
port 9 n
rlabel metal1 10 8635 10 8635 1 VDD
port 2 n
rlabel metal1 -2135 7425 -2135 7425 1 Vin_p
port 4 n
rlabel metal1 -1075 6275 -1075 6275 1 Vout_p
port 5 n
rlabel metal1 -5140 8635 -5140 8635 1 VDD
port 2 n
rlabel metal1 -4075 6275 -4075 6275 1 Vout_n
port 6 n
rlabel metal1 -3005 7425 -3005 7425 1 Vin_n
port 3 n
rlabel metal1 -5135 3650 -5135 3650 1 GND
port 9 n
<< end >>
