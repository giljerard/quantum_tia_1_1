magic
tech sky130A
timestamp 1640983407
<< dnwell >>
rect -105 -105 2815 2390
<< nwell >>
rect -145 2285 2855 2430
rect -145 0 0 2285
rect 2710 0 2855 2285
rect -145 -145 2855 0
<< pwell >>
rect 0 0 2710 2285
<< nmos >>
rect 105 -295 2605 -250
rect 105 -390 2605 -345
rect 105 -485 2605 -440
rect 105 -580 2605 -535
rect 105 -675 2605 -630
rect 105 -770 2605 -725
rect 105 -865 2605 -820
rect 105 -960 2605 -915
rect 105 -1055 2605 -1010
rect 105 -1150 2605 -1105
rect 105 -1245 2605 -1200
rect 105 -1340 2605 -1295
rect 105 -1435 2605 -1390
rect 105 -1530 2605 -1485
rect 105 -1625 2605 -1580
rect 105 -1720 2605 -1675
rect 105 -1815 2605 -1770
rect 105 -1910 2605 -1865
rect 105 -2005 2605 -1960
rect 105 -2100 2605 -2055
rect 105 -2195 2605 -2150
rect 105 -2290 2605 -2245
rect 105 -2385 2605 -2340
rect 105 -2480 2605 -2435
rect 105 -2575 2605 -2530
rect 105 -2670 2605 -2625
<< nmoslvt >>
rect 175 2150 2675 2182
rect 175 2068 2675 2100
rect 175 1986 2675 2018
rect 175 1904 2675 1936
rect 175 1822 2675 1854
rect 175 1740 2675 1772
rect 175 1658 2675 1690
rect 175 1576 2675 1608
rect 175 1494 2675 1526
rect 175 1412 2675 1444
rect 175 1330 2675 1362
rect 175 1248 2675 1280
rect 175 1166 2675 1198
rect 175 1084 2675 1116
rect 175 1002 2675 1034
rect 175 920 2675 952
rect 175 838 2675 870
rect 175 756 2675 788
rect 175 674 2675 706
rect 175 592 2675 624
rect 175 510 2675 542
rect 175 428 2675 460
rect 175 346 2675 378
rect 175 264 2675 296
rect 175 182 2675 214
rect 175 100 2675 132
<< ndiff >>
rect 175 2217 2675 2230
rect 175 2197 200 2217
rect 220 2197 240 2217
rect 260 2197 280 2217
rect 300 2197 320 2217
rect 340 2197 360 2217
rect 380 2197 400 2217
rect 420 2197 440 2217
rect 460 2197 480 2217
rect 500 2197 520 2217
rect 540 2197 560 2217
rect 580 2197 600 2217
rect 620 2197 640 2217
rect 660 2197 680 2217
rect 700 2197 720 2217
rect 740 2197 760 2217
rect 780 2197 800 2217
rect 820 2197 840 2217
rect 860 2197 880 2217
rect 900 2197 920 2217
rect 940 2197 960 2217
rect 980 2197 1000 2217
rect 1020 2197 1040 2217
rect 1060 2197 1080 2217
rect 1100 2197 1120 2217
rect 1140 2197 1160 2217
rect 1180 2197 1200 2217
rect 1220 2197 1240 2217
rect 1260 2197 1280 2217
rect 1300 2197 1320 2217
rect 1340 2197 1360 2217
rect 1380 2197 1400 2217
rect 1420 2197 1440 2217
rect 1460 2197 1480 2217
rect 1500 2197 1520 2217
rect 1540 2197 1560 2217
rect 1580 2197 1600 2217
rect 1620 2197 1640 2217
rect 1660 2197 1680 2217
rect 1700 2197 1720 2217
rect 1740 2197 1760 2217
rect 1780 2197 1800 2217
rect 1820 2197 1840 2217
rect 1860 2197 1880 2217
rect 1900 2197 1920 2217
rect 1940 2197 1960 2217
rect 1980 2197 2000 2217
rect 2020 2197 2040 2217
rect 2060 2197 2080 2217
rect 2100 2197 2120 2217
rect 2140 2197 2160 2217
rect 2180 2197 2200 2217
rect 2220 2197 2240 2217
rect 2260 2197 2280 2217
rect 2300 2197 2320 2217
rect 2340 2197 2360 2217
rect 2380 2197 2400 2217
rect 2420 2197 2440 2217
rect 2460 2197 2480 2217
rect 2500 2197 2520 2217
rect 2540 2197 2560 2217
rect 2580 2197 2600 2217
rect 2620 2197 2640 2217
rect 2660 2197 2675 2217
rect 175 2182 2675 2197
rect 175 2135 2675 2150
rect 175 2115 200 2135
rect 220 2115 240 2135
rect 260 2115 280 2135
rect 300 2115 320 2135
rect 340 2115 360 2135
rect 380 2115 400 2135
rect 420 2115 440 2135
rect 460 2115 480 2135
rect 500 2115 520 2135
rect 540 2115 560 2135
rect 580 2115 600 2135
rect 620 2115 640 2135
rect 660 2115 680 2135
rect 700 2115 720 2135
rect 740 2115 760 2135
rect 780 2115 800 2135
rect 820 2115 840 2135
rect 860 2115 880 2135
rect 900 2115 920 2135
rect 940 2115 960 2135
rect 980 2115 1000 2135
rect 1020 2115 1040 2135
rect 1060 2115 1080 2135
rect 1100 2115 1120 2135
rect 1140 2115 1160 2135
rect 1180 2115 1200 2135
rect 1220 2115 1240 2135
rect 1260 2115 1280 2135
rect 1300 2115 1320 2135
rect 1340 2115 1360 2135
rect 1380 2115 1400 2135
rect 1420 2115 1440 2135
rect 1460 2115 1480 2135
rect 1500 2115 1520 2135
rect 1540 2115 1560 2135
rect 1580 2115 1600 2135
rect 1620 2115 1640 2135
rect 1660 2115 1680 2135
rect 1700 2115 1720 2135
rect 1740 2115 1760 2135
rect 1780 2115 1800 2135
rect 1820 2115 1840 2135
rect 1860 2115 1880 2135
rect 1900 2115 1920 2135
rect 1940 2115 1960 2135
rect 1980 2115 2000 2135
rect 2020 2115 2040 2135
rect 2060 2115 2080 2135
rect 2100 2115 2120 2135
rect 2140 2115 2160 2135
rect 2180 2115 2200 2135
rect 2220 2115 2240 2135
rect 2260 2115 2280 2135
rect 2300 2115 2320 2135
rect 2340 2115 2360 2135
rect 2380 2115 2400 2135
rect 2420 2115 2440 2135
rect 2460 2115 2480 2135
rect 2500 2115 2520 2135
rect 2540 2115 2560 2135
rect 2580 2115 2600 2135
rect 2620 2115 2640 2135
rect 2660 2115 2675 2135
rect 175 2100 2675 2115
rect 175 2053 2675 2068
rect 175 2033 200 2053
rect 220 2033 240 2053
rect 260 2033 280 2053
rect 300 2033 320 2053
rect 340 2033 360 2053
rect 380 2033 400 2053
rect 420 2033 440 2053
rect 460 2033 480 2053
rect 500 2033 520 2053
rect 540 2033 560 2053
rect 580 2033 600 2053
rect 620 2033 640 2053
rect 660 2033 680 2053
rect 700 2033 720 2053
rect 740 2033 760 2053
rect 780 2033 800 2053
rect 820 2033 840 2053
rect 860 2033 880 2053
rect 900 2033 920 2053
rect 940 2033 960 2053
rect 980 2033 1000 2053
rect 1020 2033 1040 2053
rect 1060 2033 1080 2053
rect 1100 2033 1120 2053
rect 1140 2033 1160 2053
rect 1180 2033 1200 2053
rect 1220 2033 1240 2053
rect 1260 2033 1280 2053
rect 1300 2033 1320 2053
rect 1340 2033 1360 2053
rect 1380 2033 1400 2053
rect 1420 2033 1440 2053
rect 1460 2033 1480 2053
rect 1500 2033 1520 2053
rect 1540 2033 1560 2053
rect 1580 2033 1600 2053
rect 1620 2033 1640 2053
rect 1660 2033 1680 2053
rect 1700 2033 1720 2053
rect 1740 2033 1760 2053
rect 1780 2033 1800 2053
rect 1820 2033 1840 2053
rect 1860 2033 1880 2053
rect 1900 2033 1920 2053
rect 1940 2033 1960 2053
rect 1980 2033 2000 2053
rect 2020 2033 2040 2053
rect 2060 2033 2080 2053
rect 2100 2033 2120 2053
rect 2140 2033 2160 2053
rect 2180 2033 2200 2053
rect 2220 2033 2240 2053
rect 2260 2033 2280 2053
rect 2300 2033 2320 2053
rect 2340 2033 2360 2053
rect 2380 2033 2400 2053
rect 2420 2033 2440 2053
rect 2460 2033 2480 2053
rect 2500 2033 2520 2053
rect 2540 2033 2560 2053
rect 2580 2033 2600 2053
rect 2620 2033 2640 2053
rect 2660 2033 2675 2053
rect 175 2018 2675 2033
rect 175 1971 2675 1986
rect 175 1951 200 1971
rect 220 1951 240 1971
rect 260 1951 280 1971
rect 300 1951 320 1971
rect 340 1951 360 1971
rect 380 1951 400 1971
rect 420 1951 440 1971
rect 460 1951 480 1971
rect 500 1951 520 1971
rect 540 1951 560 1971
rect 580 1951 600 1971
rect 620 1951 640 1971
rect 660 1951 680 1971
rect 700 1951 720 1971
rect 740 1951 760 1971
rect 780 1951 800 1971
rect 820 1951 840 1971
rect 860 1951 880 1971
rect 900 1951 920 1971
rect 940 1951 960 1971
rect 980 1951 1000 1971
rect 1020 1951 1040 1971
rect 1060 1951 1080 1971
rect 1100 1951 1120 1971
rect 1140 1951 1160 1971
rect 1180 1951 1200 1971
rect 1220 1951 1240 1971
rect 1260 1951 1280 1971
rect 1300 1951 1320 1971
rect 1340 1951 1360 1971
rect 1380 1951 1400 1971
rect 1420 1951 1440 1971
rect 1460 1951 1480 1971
rect 1500 1951 1520 1971
rect 1540 1951 1560 1971
rect 1580 1951 1600 1971
rect 1620 1951 1640 1971
rect 1660 1951 1680 1971
rect 1700 1951 1720 1971
rect 1740 1951 1760 1971
rect 1780 1951 1800 1971
rect 1820 1951 1840 1971
rect 1860 1951 1880 1971
rect 1900 1951 1920 1971
rect 1940 1951 1960 1971
rect 1980 1951 2000 1971
rect 2020 1951 2040 1971
rect 2060 1951 2080 1971
rect 2100 1951 2120 1971
rect 2140 1951 2160 1971
rect 2180 1951 2200 1971
rect 2220 1951 2240 1971
rect 2260 1951 2280 1971
rect 2300 1951 2320 1971
rect 2340 1951 2360 1971
rect 2380 1951 2400 1971
rect 2420 1951 2440 1971
rect 2460 1951 2480 1971
rect 2500 1951 2520 1971
rect 2540 1951 2560 1971
rect 2580 1951 2600 1971
rect 2620 1951 2640 1971
rect 2660 1951 2675 1971
rect 175 1936 2675 1951
rect 175 1889 2675 1904
rect 175 1869 200 1889
rect 220 1869 240 1889
rect 260 1869 280 1889
rect 300 1869 320 1889
rect 340 1869 360 1889
rect 380 1869 400 1889
rect 420 1869 440 1889
rect 460 1869 480 1889
rect 500 1869 520 1889
rect 540 1869 560 1889
rect 580 1869 600 1889
rect 620 1869 640 1889
rect 660 1869 680 1889
rect 700 1869 720 1889
rect 740 1869 760 1889
rect 780 1869 800 1889
rect 820 1869 840 1889
rect 860 1869 880 1889
rect 900 1869 920 1889
rect 940 1869 960 1889
rect 980 1869 1000 1889
rect 1020 1869 1040 1889
rect 1060 1869 1080 1889
rect 1100 1869 1120 1889
rect 1140 1869 1160 1889
rect 1180 1869 1200 1889
rect 1220 1869 1240 1889
rect 1260 1869 1280 1889
rect 1300 1869 1320 1889
rect 1340 1869 1360 1889
rect 1380 1869 1400 1889
rect 1420 1869 1440 1889
rect 1460 1869 1480 1889
rect 1500 1869 1520 1889
rect 1540 1869 1560 1889
rect 1580 1869 1600 1889
rect 1620 1869 1640 1889
rect 1660 1869 1680 1889
rect 1700 1869 1720 1889
rect 1740 1869 1760 1889
rect 1780 1869 1800 1889
rect 1820 1869 1840 1889
rect 1860 1869 1880 1889
rect 1900 1869 1920 1889
rect 1940 1869 1960 1889
rect 1980 1869 2000 1889
rect 2020 1869 2040 1889
rect 2060 1869 2080 1889
rect 2100 1869 2120 1889
rect 2140 1869 2160 1889
rect 2180 1869 2200 1889
rect 2220 1869 2240 1889
rect 2260 1869 2280 1889
rect 2300 1869 2320 1889
rect 2340 1869 2360 1889
rect 2380 1869 2400 1889
rect 2420 1869 2440 1889
rect 2460 1869 2480 1889
rect 2500 1869 2520 1889
rect 2540 1869 2560 1889
rect 2580 1869 2600 1889
rect 2620 1869 2640 1889
rect 2660 1869 2675 1889
rect 175 1854 2675 1869
rect 175 1807 2675 1822
rect 175 1787 200 1807
rect 220 1787 240 1807
rect 260 1787 280 1807
rect 300 1787 320 1807
rect 340 1787 360 1807
rect 380 1787 400 1807
rect 420 1787 440 1807
rect 460 1787 480 1807
rect 500 1787 520 1807
rect 540 1787 560 1807
rect 580 1787 600 1807
rect 620 1787 640 1807
rect 660 1787 680 1807
rect 700 1787 720 1807
rect 740 1787 760 1807
rect 780 1787 800 1807
rect 820 1787 840 1807
rect 860 1787 880 1807
rect 900 1787 920 1807
rect 940 1787 960 1807
rect 980 1787 1000 1807
rect 1020 1787 1040 1807
rect 1060 1787 1080 1807
rect 1100 1787 1120 1807
rect 1140 1787 1160 1807
rect 1180 1787 1200 1807
rect 1220 1787 1240 1807
rect 1260 1787 1280 1807
rect 1300 1787 1320 1807
rect 1340 1787 1360 1807
rect 1380 1787 1400 1807
rect 1420 1787 1440 1807
rect 1460 1787 1480 1807
rect 1500 1787 1520 1807
rect 1540 1787 1560 1807
rect 1580 1787 1600 1807
rect 1620 1787 1640 1807
rect 1660 1787 1680 1807
rect 1700 1787 1720 1807
rect 1740 1787 1760 1807
rect 1780 1787 1800 1807
rect 1820 1787 1840 1807
rect 1860 1787 1880 1807
rect 1900 1787 1920 1807
rect 1940 1787 1960 1807
rect 1980 1787 2000 1807
rect 2020 1787 2040 1807
rect 2060 1787 2080 1807
rect 2100 1787 2120 1807
rect 2140 1787 2160 1807
rect 2180 1787 2200 1807
rect 2220 1787 2240 1807
rect 2260 1787 2280 1807
rect 2300 1787 2320 1807
rect 2340 1787 2360 1807
rect 2380 1787 2400 1807
rect 2420 1787 2440 1807
rect 2460 1787 2480 1807
rect 2500 1787 2520 1807
rect 2540 1787 2560 1807
rect 2580 1787 2600 1807
rect 2620 1787 2640 1807
rect 2660 1787 2675 1807
rect 175 1772 2675 1787
rect 175 1725 2675 1740
rect 175 1705 200 1725
rect 220 1705 240 1725
rect 260 1705 280 1725
rect 300 1705 320 1725
rect 340 1705 360 1725
rect 380 1705 400 1725
rect 420 1705 440 1725
rect 460 1705 480 1725
rect 500 1705 520 1725
rect 540 1705 560 1725
rect 580 1705 600 1725
rect 620 1705 640 1725
rect 660 1705 680 1725
rect 700 1705 720 1725
rect 740 1705 760 1725
rect 780 1705 800 1725
rect 820 1705 840 1725
rect 860 1705 880 1725
rect 900 1705 920 1725
rect 940 1705 960 1725
rect 980 1705 1000 1725
rect 1020 1705 1040 1725
rect 1060 1705 1080 1725
rect 1100 1705 1120 1725
rect 1140 1705 1160 1725
rect 1180 1705 1200 1725
rect 1220 1705 1240 1725
rect 1260 1705 1280 1725
rect 1300 1705 1320 1725
rect 1340 1705 1360 1725
rect 1380 1705 1400 1725
rect 1420 1705 1440 1725
rect 1460 1705 1480 1725
rect 1500 1705 1520 1725
rect 1540 1705 1560 1725
rect 1580 1705 1600 1725
rect 1620 1705 1640 1725
rect 1660 1705 1680 1725
rect 1700 1705 1720 1725
rect 1740 1705 1760 1725
rect 1780 1705 1800 1725
rect 1820 1705 1840 1725
rect 1860 1705 1880 1725
rect 1900 1705 1920 1725
rect 1940 1705 1960 1725
rect 1980 1705 2000 1725
rect 2020 1705 2040 1725
rect 2060 1705 2080 1725
rect 2100 1705 2120 1725
rect 2140 1705 2160 1725
rect 2180 1705 2200 1725
rect 2220 1705 2240 1725
rect 2260 1705 2280 1725
rect 2300 1705 2320 1725
rect 2340 1705 2360 1725
rect 2380 1705 2400 1725
rect 2420 1705 2440 1725
rect 2460 1705 2480 1725
rect 2500 1705 2520 1725
rect 2540 1705 2560 1725
rect 2580 1705 2600 1725
rect 2620 1705 2640 1725
rect 2660 1705 2675 1725
rect 175 1690 2675 1705
rect 175 1643 2675 1658
rect 175 1623 200 1643
rect 220 1623 240 1643
rect 260 1623 280 1643
rect 300 1623 320 1643
rect 340 1623 360 1643
rect 380 1623 400 1643
rect 420 1623 440 1643
rect 460 1623 480 1643
rect 500 1623 520 1643
rect 540 1623 560 1643
rect 580 1623 600 1643
rect 620 1623 640 1643
rect 660 1623 680 1643
rect 700 1623 720 1643
rect 740 1623 760 1643
rect 780 1623 800 1643
rect 820 1623 840 1643
rect 860 1623 880 1643
rect 900 1623 920 1643
rect 940 1623 960 1643
rect 980 1623 1000 1643
rect 1020 1623 1040 1643
rect 1060 1623 1080 1643
rect 1100 1623 1120 1643
rect 1140 1623 1160 1643
rect 1180 1623 1200 1643
rect 1220 1623 1240 1643
rect 1260 1623 1280 1643
rect 1300 1623 1320 1643
rect 1340 1623 1360 1643
rect 1380 1623 1400 1643
rect 1420 1623 1440 1643
rect 1460 1623 1480 1643
rect 1500 1623 1520 1643
rect 1540 1623 1560 1643
rect 1580 1623 1600 1643
rect 1620 1623 1640 1643
rect 1660 1623 1680 1643
rect 1700 1623 1720 1643
rect 1740 1623 1760 1643
rect 1780 1623 1800 1643
rect 1820 1623 1840 1643
rect 1860 1623 1880 1643
rect 1900 1623 1920 1643
rect 1940 1623 1960 1643
rect 1980 1623 2000 1643
rect 2020 1623 2040 1643
rect 2060 1623 2080 1643
rect 2100 1623 2120 1643
rect 2140 1623 2160 1643
rect 2180 1623 2200 1643
rect 2220 1623 2240 1643
rect 2260 1623 2280 1643
rect 2300 1623 2320 1643
rect 2340 1623 2360 1643
rect 2380 1623 2400 1643
rect 2420 1623 2440 1643
rect 2460 1623 2480 1643
rect 2500 1623 2520 1643
rect 2540 1623 2560 1643
rect 2580 1623 2600 1643
rect 2620 1623 2640 1643
rect 2660 1623 2675 1643
rect 175 1608 2675 1623
rect 175 1561 2675 1576
rect 175 1541 200 1561
rect 220 1541 240 1561
rect 260 1541 280 1561
rect 300 1541 320 1561
rect 340 1541 360 1561
rect 380 1541 400 1561
rect 420 1541 440 1561
rect 460 1541 480 1561
rect 500 1541 520 1561
rect 540 1541 560 1561
rect 580 1541 600 1561
rect 620 1541 640 1561
rect 660 1541 680 1561
rect 700 1541 720 1561
rect 740 1541 760 1561
rect 780 1541 800 1561
rect 820 1541 840 1561
rect 860 1541 880 1561
rect 900 1541 920 1561
rect 940 1541 960 1561
rect 980 1541 1000 1561
rect 1020 1541 1040 1561
rect 1060 1541 1080 1561
rect 1100 1541 1120 1561
rect 1140 1541 1160 1561
rect 1180 1541 1200 1561
rect 1220 1541 1240 1561
rect 1260 1541 1280 1561
rect 1300 1541 1320 1561
rect 1340 1541 1360 1561
rect 1380 1541 1400 1561
rect 1420 1541 1440 1561
rect 1460 1541 1480 1561
rect 1500 1541 1520 1561
rect 1540 1541 1560 1561
rect 1580 1541 1600 1561
rect 1620 1541 1640 1561
rect 1660 1541 1680 1561
rect 1700 1541 1720 1561
rect 1740 1541 1760 1561
rect 1780 1541 1800 1561
rect 1820 1541 1840 1561
rect 1860 1541 1880 1561
rect 1900 1541 1920 1561
rect 1940 1541 1960 1561
rect 1980 1541 2000 1561
rect 2020 1541 2040 1561
rect 2060 1541 2080 1561
rect 2100 1541 2120 1561
rect 2140 1541 2160 1561
rect 2180 1541 2200 1561
rect 2220 1541 2240 1561
rect 2260 1541 2280 1561
rect 2300 1541 2320 1561
rect 2340 1541 2360 1561
rect 2380 1541 2400 1561
rect 2420 1541 2440 1561
rect 2460 1541 2480 1561
rect 2500 1541 2520 1561
rect 2540 1541 2560 1561
rect 2580 1541 2600 1561
rect 2620 1541 2640 1561
rect 2660 1541 2675 1561
rect 175 1526 2675 1541
rect 175 1479 2675 1494
rect 175 1459 200 1479
rect 220 1459 240 1479
rect 260 1459 280 1479
rect 300 1459 320 1479
rect 340 1459 360 1479
rect 380 1459 400 1479
rect 420 1459 440 1479
rect 460 1459 480 1479
rect 500 1459 520 1479
rect 540 1459 560 1479
rect 580 1459 600 1479
rect 620 1459 640 1479
rect 660 1459 680 1479
rect 700 1459 720 1479
rect 740 1459 760 1479
rect 780 1459 800 1479
rect 820 1459 840 1479
rect 860 1459 880 1479
rect 900 1459 920 1479
rect 940 1459 960 1479
rect 980 1459 1000 1479
rect 1020 1459 1040 1479
rect 1060 1459 1080 1479
rect 1100 1459 1120 1479
rect 1140 1459 1160 1479
rect 1180 1459 1200 1479
rect 1220 1459 1240 1479
rect 1260 1459 1280 1479
rect 1300 1459 1320 1479
rect 1340 1459 1360 1479
rect 1380 1459 1400 1479
rect 1420 1459 1440 1479
rect 1460 1459 1480 1479
rect 1500 1459 1520 1479
rect 1540 1459 1560 1479
rect 1580 1459 1600 1479
rect 1620 1459 1640 1479
rect 1660 1459 1680 1479
rect 1700 1459 1720 1479
rect 1740 1459 1760 1479
rect 1780 1459 1800 1479
rect 1820 1459 1840 1479
rect 1860 1459 1880 1479
rect 1900 1459 1920 1479
rect 1940 1459 1960 1479
rect 1980 1459 2000 1479
rect 2020 1459 2040 1479
rect 2060 1459 2080 1479
rect 2100 1459 2120 1479
rect 2140 1459 2160 1479
rect 2180 1459 2200 1479
rect 2220 1459 2240 1479
rect 2260 1459 2280 1479
rect 2300 1459 2320 1479
rect 2340 1459 2360 1479
rect 2380 1459 2400 1479
rect 2420 1459 2440 1479
rect 2460 1459 2480 1479
rect 2500 1459 2520 1479
rect 2540 1459 2560 1479
rect 2580 1459 2600 1479
rect 2620 1459 2640 1479
rect 2660 1459 2675 1479
rect 175 1444 2675 1459
rect 175 1397 2675 1412
rect 175 1377 200 1397
rect 220 1377 240 1397
rect 260 1377 280 1397
rect 300 1377 320 1397
rect 340 1377 360 1397
rect 380 1377 400 1397
rect 420 1377 440 1397
rect 460 1377 480 1397
rect 500 1377 520 1397
rect 540 1377 560 1397
rect 580 1377 600 1397
rect 620 1377 640 1397
rect 660 1377 680 1397
rect 700 1377 720 1397
rect 740 1377 760 1397
rect 780 1377 800 1397
rect 820 1377 840 1397
rect 860 1377 880 1397
rect 900 1377 920 1397
rect 940 1377 960 1397
rect 980 1377 1000 1397
rect 1020 1377 1040 1397
rect 1060 1377 1080 1397
rect 1100 1377 1120 1397
rect 1140 1377 1160 1397
rect 1180 1377 1200 1397
rect 1220 1377 1240 1397
rect 1260 1377 1280 1397
rect 1300 1377 1320 1397
rect 1340 1377 1360 1397
rect 1380 1377 1400 1397
rect 1420 1377 1440 1397
rect 1460 1377 1480 1397
rect 1500 1377 1520 1397
rect 1540 1377 1560 1397
rect 1580 1377 1600 1397
rect 1620 1377 1640 1397
rect 1660 1377 1680 1397
rect 1700 1377 1720 1397
rect 1740 1377 1760 1397
rect 1780 1377 1800 1397
rect 1820 1377 1840 1397
rect 1860 1377 1880 1397
rect 1900 1377 1920 1397
rect 1940 1377 1960 1397
rect 1980 1377 2000 1397
rect 2020 1377 2040 1397
rect 2060 1377 2080 1397
rect 2100 1377 2120 1397
rect 2140 1377 2160 1397
rect 2180 1377 2200 1397
rect 2220 1377 2240 1397
rect 2260 1377 2280 1397
rect 2300 1377 2320 1397
rect 2340 1377 2360 1397
rect 2380 1377 2400 1397
rect 2420 1377 2440 1397
rect 2460 1377 2480 1397
rect 2500 1377 2520 1397
rect 2540 1377 2560 1397
rect 2580 1377 2600 1397
rect 2620 1377 2640 1397
rect 2660 1377 2675 1397
rect 175 1362 2675 1377
rect 175 1315 2675 1330
rect 175 1295 200 1315
rect 220 1295 240 1315
rect 260 1295 280 1315
rect 300 1295 320 1315
rect 340 1295 360 1315
rect 380 1295 400 1315
rect 420 1295 440 1315
rect 460 1295 480 1315
rect 500 1295 520 1315
rect 540 1295 560 1315
rect 580 1295 600 1315
rect 620 1295 640 1315
rect 660 1295 680 1315
rect 700 1295 720 1315
rect 740 1295 760 1315
rect 780 1295 800 1315
rect 820 1295 840 1315
rect 860 1295 880 1315
rect 900 1295 920 1315
rect 940 1295 960 1315
rect 980 1295 1000 1315
rect 1020 1295 1040 1315
rect 1060 1295 1080 1315
rect 1100 1295 1120 1315
rect 1140 1295 1160 1315
rect 1180 1295 1200 1315
rect 1220 1295 1240 1315
rect 1260 1295 1280 1315
rect 1300 1295 1320 1315
rect 1340 1295 1360 1315
rect 1380 1295 1400 1315
rect 1420 1295 1440 1315
rect 1460 1295 1480 1315
rect 1500 1295 1520 1315
rect 1540 1295 1560 1315
rect 1580 1295 1600 1315
rect 1620 1295 1640 1315
rect 1660 1295 1680 1315
rect 1700 1295 1720 1315
rect 1740 1295 1760 1315
rect 1780 1295 1800 1315
rect 1820 1295 1840 1315
rect 1860 1295 1880 1315
rect 1900 1295 1920 1315
rect 1940 1295 1960 1315
rect 1980 1295 2000 1315
rect 2020 1295 2040 1315
rect 2060 1295 2080 1315
rect 2100 1295 2120 1315
rect 2140 1295 2160 1315
rect 2180 1295 2200 1315
rect 2220 1295 2240 1315
rect 2260 1295 2280 1315
rect 2300 1295 2320 1315
rect 2340 1295 2360 1315
rect 2380 1295 2400 1315
rect 2420 1295 2440 1315
rect 2460 1295 2480 1315
rect 2500 1295 2520 1315
rect 2540 1295 2560 1315
rect 2580 1295 2600 1315
rect 2620 1295 2640 1315
rect 2660 1295 2675 1315
rect 175 1280 2675 1295
rect 175 1233 2675 1248
rect 175 1213 200 1233
rect 220 1213 240 1233
rect 260 1213 280 1233
rect 300 1213 320 1233
rect 340 1213 360 1233
rect 380 1213 400 1233
rect 420 1213 440 1233
rect 460 1213 480 1233
rect 500 1213 520 1233
rect 540 1213 560 1233
rect 580 1213 600 1233
rect 620 1213 640 1233
rect 660 1213 680 1233
rect 700 1213 720 1233
rect 740 1213 760 1233
rect 780 1213 800 1233
rect 820 1213 840 1233
rect 860 1213 880 1233
rect 900 1213 920 1233
rect 940 1213 960 1233
rect 980 1213 1000 1233
rect 1020 1213 1040 1233
rect 1060 1213 1080 1233
rect 1100 1213 1120 1233
rect 1140 1213 1160 1233
rect 1180 1213 1200 1233
rect 1220 1213 1240 1233
rect 1260 1213 1280 1233
rect 1300 1213 1320 1233
rect 1340 1213 1360 1233
rect 1380 1213 1400 1233
rect 1420 1213 1440 1233
rect 1460 1213 1480 1233
rect 1500 1213 1520 1233
rect 1540 1213 1560 1233
rect 1580 1213 1600 1233
rect 1620 1213 1640 1233
rect 1660 1213 1680 1233
rect 1700 1213 1720 1233
rect 1740 1213 1760 1233
rect 1780 1213 1800 1233
rect 1820 1213 1840 1233
rect 1860 1213 1880 1233
rect 1900 1213 1920 1233
rect 1940 1213 1960 1233
rect 1980 1213 2000 1233
rect 2020 1213 2040 1233
rect 2060 1213 2080 1233
rect 2100 1213 2120 1233
rect 2140 1213 2160 1233
rect 2180 1213 2200 1233
rect 2220 1213 2240 1233
rect 2260 1213 2280 1233
rect 2300 1213 2320 1233
rect 2340 1213 2360 1233
rect 2380 1213 2400 1233
rect 2420 1213 2440 1233
rect 2460 1213 2480 1233
rect 2500 1213 2520 1233
rect 2540 1213 2560 1233
rect 2580 1213 2600 1233
rect 2620 1213 2640 1233
rect 2660 1213 2675 1233
rect 175 1198 2675 1213
rect 175 1151 2675 1166
rect 175 1131 200 1151
rect 220 1131 240 1151
rect 260 1131 280 1151
rect 300 1131 320 1151
rect 340 1131 360 1151
rect 380 1131 400 1151
rect 420 1131 440 1151
rect 460 1131 480 1151
rect 500 1131 520 1151
rect 540 1131 560 1151
rect 580 1131 600 1151
rect 620 1131 640 1151
rect 660 1131 680 1151
rect 700 1131 720 1151
rect 740 1131 760 1151
rect 780 1131 800 1151
rect 820 1131 840 1151
rect 860 1131 880 1151
rect 900 1131 920 1151
rect 940 1131 960 1151
rect 980 1131 1000 1151
rect 1020 1131 1040 1151
rect 1060 1131 1080 1151
rect 1100 1131 1120 1151
rect 1140 1131 1160 1151
rect 1180 1131 1200 1151
rect 1220 1131 1240 1151
rect 1260 1131 1280 1151
rect 1300 1131 1320 1151
rect 1340 1131 1360 1151
rect 1380 1131 1400 1151
rect 1420 1131 1440 1151
rect 1460 1131 1480 1151
rect 1500 1131 1520 1151
rect 1540 1131 1560 1151
rect 1580 1131 1600 1151
rect 1620 1131 1640 1151
rect 1660 1131 1680 1151
rect 1700 1131 1720 1151
rect 1740 1131 1760 1151
rect 1780 1131 1800 1151
rect 1820 1131 1840 1151
rect 1860 1131 1880 1151
rect 1900 1131 1920 1151
rect 1940 1131 1960 1151
rect 1980 1131 2000 1151
rect 2020 1131 2040 1151
rect 2060 1131 2080 1151
rect 2100 1131 2120 1151
rect 2140 1131 2160 1151
rect 2180 1131 2200 1151
rect 2220 1131 2240 1151
rect 2260 1131 2280 1151
rect 2300 1131 2320 1151
rect 2340 1131 2360 1151
rect 2380 1131 2400 1151
rect 2420 1131 2440 1151
rect 2460 1131 2480 1151
rect 2500 1131 2520 1151
rect 2540 1131 2560 1151
rect 2580 1131 2600 1151
rect 2620 1131 2640 1151
rect 2660 1131 2675 1151
rect 175 1116 2675 1131
rect 175 1069 2675 1084
rect 175 1049 200 1069
rect 220 1049 240 1069
rect 260 1049 280 1069
rect 300 1049 320 1069
rect 340 1049 360 1069
rect 380 1049 400 1069
rect 420 1049 440 1069
rect 460 1049 480 1069
rect 500 1049 520 1069
rect 540 1049 560 1069
rect 580 1049 600 1069
rect 620 1049 640 1069
rect 660 1049 680 1069
rect 700 1049 720 1069
rect 740 1049 760 1069
rect 780 1049 800 1069
rect 820 1049 840 1069
rect 860 1049 880 1069
rect 900 1049 920 1069
rect 940 1049 960 1069
rect 980 1049 1000 1069
rect 1020 1049 1040 1069
rect 1060 1049 1080 1069
rect 1100 1049 1120 1069
rect 1140 1049 1160 1069
rect 1180 1049 1200 1069
rect 1220 1049 1240 1069
rect 1260 1049 1280 1069
rect 1300 1049 1320 1069
rect 1340 1049 1360 1069
rect 1380 1049 1400 1069
rect 1420 1049 1440 1069
rect 1460 1049 1480 1069
rect 1500 1049 1520 1069
rect 1540 1049 1560 1069
rect 1580 1049 1600 1069
rect 1620 1049 1640 1069
rect 1660 1049 1680 1069
rect 1700 1049 1720 1069
rect 1740 1049 1760 1069
rect 1780 1049 1800 1069
rect 1820 1049 1840 1069
rect 1860 1049 1880 1069
rect 1900 1049 1920 1069
rect 1940 1049 1960 1069
rect 1980 1049 2000 1069
rect 2020 1049 2040 1069
rect 2060 1049 2080 1069
rect 2100 1049 2120 1069
rect 2140 1049 2160 1069
rect 2180 1049 2200 1069
rect 2220 1049 2240 1069
rect 2260 1049 2280 1069
rect 2300 1049 2320 1069
rect 2340 1049 2360 1069
rect 2380 1049 2400 1069
rect 2420 1049 2440 1069
rect 2460 1049 2480 1069
rect 2500 1049 2520 1069
rect 2540 1049 2560 1069
rect 2580 1049 2600 1069
rect 2620 1049 2640 1069
rect 2660 1049 2675 1069
rect 175 1034 2675 1049
rect 175 987 2675 1002
rect 175 967 200 987
rect 220 967 240 987
rect 260 967 280 987
rect 300 967 320 987
rect 340 967 360 987
rect 380 967 400 987
rect 420 967 440 987
rect 460 967 480 987
rect 500 967 520 987
rect 540 967 560 987
rect 580 967 600 987
rect 620 967 640 987
rect 660 967 680 987
rect 700 967 720 987
rect 740 967 760 987
rect 780 967 800 987
rect 820 967 840 987
rect 860 967 880 987
rect 900 967 920 987
rect 940 967 960 987
rect 980 967 1000 987
rect 1020 967 1040 987
rect 1060 967 1080 987
rect 1100 967 1120 987
rect 1140 967 1160 987
rect 1180 967 1200 987
rect 1220 967 1240 987
rect 1260 967 1280 987
rect 1300 967 1320 987
rect 1340 967 1360 987
rect 1380 967 1400 987
rect 1420 967 1440 987
rect 1460 967 1480 987
rect 1500 967 1520 987
rect 1540 967 1560 987
rect 1580 967 1600 987
rect 1620 967 1640 987
rect 1660 967 1680 987
rect 1700 967 1720 987
rect 1740 967 1760 987
rect 1780 967 1800 987
rect 1820 967 1840 987
rect 1860 967 1880 987
rect 1900 967 1920 987
rect 1940 967 1960 987
rect 1980 967 2000 987
rect 2020 967 2040 987
rect 2060 967 2080 987
rect 2100 967 2120 987
rect 2140 967 2160 987
rect 2180 967 2200 987
rect 2220 967 2240 987
rect 2260 967 2280 987
rect 2300 967 2320 987
rect 2340 967 2360 987
rect 2380 967 2400 987
rect 2420 967 2440 987
rect 2460 967 2480 987
rect 2500 967 2520 987
rect 2540 967 2560 987
rect 2580 967 2600 987
rect 2620 967 2640 987
rect 2660 967 2675 987
rect 175 952 2675 967
rect 175 905 2675 920
rect 175 885 200 905
rect 220 885 240 905
rect 260 885 280 905
rect 300 885 320 905
rect 340 885 360 905
rect 380 885 400 905
rect 420 885 440 905
rect 460 885 480 905
rect 500 885 520 905
rect 540 885 560 905
rect 580 885 600 905
rect 620 885 640 905
rect 660 885 680 905
rect 700 885 720 905
rect 740 885 760 905
rect 780 885 800 905
rect 820 885 840 905
rect 860 885 880 905
rect 900 885 920 905
rect 940 885 960 905
rect 980 885 1000 905
rect 1020 885 1040 905
rect 1060 885 1080 905
rect 1100 885 1120 905
rect 1140 885 1160 905
rect 1180 885 1200 905
rect 1220 885 1240 905
rect 1260 885 1280 905
rect 1300 885 1320 905
rect 1340 885 1360 905
rect 1380 885 1400 905
rect 1420 885 1440 905
rect 1460 885 1480 905
rect 1500 885 1520 905
rect 1540 885 1560 905
rect 1580 885 1600 905
rect 1620 885 1640 905
rect 1660 885 1680 905
rect 1700 885 1720 905
rect 1740 885 1760 905
rect 1780 885 1800 905
rect 1820 885 1840 905
rect 1860 885 1880 905
rect 1900 885 1920 905
rect 1940 885 1960 905
rect 1980 885 2000 905
rect 2020 885 2040 905
rect 2060 885 2080 905
rect 2100 885 2120 905
rect 2140 885 2160 905
rect 2180 885 2200 905
rect 2220 885 2240 905
rect 2260 885 2280 905
rect 2300 885 2320 905
rect 2340 885 2360 905
rect 2380 885 2400 905
rect 2420 885 2440 905
rect 2460 885 2480 905
rect 2500 885 2520 905
rect 2540 885 2560 905
rect 2580 885 2600 905
rect 2620 885 2640 905
rect 2660 885 2675 905
rect 175 870 2675 885
rect 175 823 2675 838
rect 175 803 200 823
rect 220 803 240 823
rect 260 803 280 823
rect 300 803 320 823
rect 340 803 360 823
rect 380 803 400 823
rect 420 803 440 823
rect 460 803 480 823
rect 500 803 520 823
rect 540 803 560 823
rect 580 803 600 823
rect 620 803 640 823
rect 660 803 680 823
rect 700 803 720 823
rect 740 803 760 823
rect 780 803 800 823
rect 820 803 840 823
rect 860 803 880 823
rect 900 803 920 823
rect 940 803 960 823
rect 980 803 1000 823
rect 1020 803 1040 823
rect 1060 803 1080 823
rect 1100 803 1120 823
rect 1140 803 1160 823
rect 1180 803 1200 823
rect 1220 803 1240 823
rect 1260 803 1280 823
rect 1300 803 1320 823
rect 1340 803 1360 823
rect 1380 803 1400 823
rect 1420 803 1440 823
rect 1460 803 1480 823
rect 1500 803 1520 823
rect 1540 803 1560 823
rect 1580 803 1600 823
rect 1620 803 1640 823
rect 1660 803 1680 823
rect 1700 803 1720 823
rect 1740 803 1760 823
rect 1780 803 1800 823
rect 1820 803 1840 823
rect 1860 803 1880 823
rect 1900 803 1920 823
rect 1940 803 1960 823
rect 1980 803 2000 823
rect 2020 803 2040 823
rect 2060 803 2080 823
rect 2100 803 2120 823
rect 2140 803 2160 823
rect 2180 803 2200 823
rect 2220 803 2240 823
rect 2260 803 2280 823
rect 2300 803 2320 823
rect 2340 803 2360 823
rect 2380 803 2400 823
rect 2420 803 2440 823
rect 2460 803 2480 823
rect 2500 803 2520 823
rect 2540 803 2560 823
rect 2580 803 2600 823
rect 2620 803 2640 823
rect 2660 803 2675 823
rect 175 788 2675 803
rect 175 741 2675 756
rect 175 721 200 741
rect 220 721 240 741
rect 260 721 280 741
rect 300 721 320 741
rect 340 721 360 741
rect 380 721 400 741
rect 420 721 440 741
rect 460 721 480 741
rect 500 721 520 741
rect 540 721 560 741
rect 580 721 600 741
rect 620 721 640 741
rect 660 721 680 741
rect 700 721 720 741
rect 740 721 760 741
rect 780 721 800 741
rect 820 721 840 741
rect 860 721 880 741
rect 900 721 920 741
rect 940 721 960 741
rect 980 721 1000 741
rect 1020 721 1040 741
rect 1060 721 1080 741
rect 1100 721 1120 741
rect 1140 721 1160 741
rect 1180 721 1200 741
rect 1220 721 1240 741
rect 1260 721 1280 741
rect 1300 721 1320 741
rect 1340 721 1360 741
rect 1380 721 1400 741
rect 1420 721 1440 741
rect 1460 721 1480 741
rect 1500 721 1520 741
rect 1540 721 1560 741
rect 1580 721 1600 741
rect 1620 721 1640 741
rect 1660 721 1680 741
rect 1700 721 1720 741
rect 1740 721 1760 741
rect 1780 721 1800 741
rect 1820 721 1840 741
rect 1860 721 1880 741
rect 1900 721 1920 741
rect 1940 721 1960 741
rect 1980 721 2000 741
rect 2020 721 2040 741
rect 2060 721 2080 741
rect 2100 721 2120 741
rect 2140 721 2160 741
rect 2180 721 2200 741
rect 2220 721 2240 741
rect 2260 721 2280 741
rect 2300 721 2320 741
rect 2340 721 2360 741
rect 2380 721 2400 741
rect 2420 721 2440 741
rect 2460 721 2480 741
rect 2500 721 2520 741
rect 2540 721 2560 741
rect 2580 721 2600 741
rect 2620 721 2640 741
rect 2660 721 2675 741
rect 175 706 2675 721
rect 175 659 2675 674
rect 175 639 200 659
rect 220 639 240 659
rect 260 639 280 659
rect 300 639 320 659
rect 340 639 360 659
rect 380 639 400 659
rect 420 639 440 659
rect 460 639 480 659
rect 500 639 520 659
rect 540 639 560 659
rect 580 639 600 659
rect 620 639 640 659
rect 660 639 680 659
rect 700 639 720 659
rect 740 639 760 659
rect 780 639 800 659
rect 820 639 840 659
rect 860 639 880 659
rect 900 639 920 659
rect 940 639 960 659
rect 980 639 1000 659
rect 1020 639 1040 659
rect 1060 639 1080 659
rect 1100 639 1120 659
rect 1140 639 1160 659
rect 1180 639 1200 659
rect 1220 639 1240 659
rect 1260 639 1280 659
rect 1300 639 1320 659
rect 1340 639 1360 659
rect 1380 639 1400 659
rect 1420 639 1440 659
rect 1460 639 1480 659
rect 1500 639 1520 659
rect 1540 639 1560 659
rect 1580 639 1600 659
rect 1620 639 1640 659
rect 1660 639 1680 659
rect 1700 639 1720 659
rect 1740 639 1760 659
rect 1780 639 1800 659
rect 1820 639 1840 659
rect 1860 639 1880 659
rect 1900 639 1920 659
rect 1940 639 1960 659
rect 1980 639 2000 659
rect 2020 639 2040 659
rect 2060 639 2080 659
rect 2100 639 2120 659
rect 2140 639 2160 659
rect 2180 639 2200 659
rect 2220 639 2240 659
rect 2260 639 2280 659
rect 2300 639 2320 659
rect 2340 639 2360 659
rect 2380 639 2400 659
rect 2420 639 2440 659
rect 2460 639 2480 659
rect 2500 639 2520 659
rect 2540 639 2560 659
rect 2580 639 2600 659
rect 2620 639 2640 659
rect 2660 639 2675 659
rect 175 624 2675 639
rect 175 577 2675 592
rect 175 557 200 577
rect 220 557 240 577
rect 260 557 280 577
rect 300 557 320 577
rect 340 557 360 577
rect 380 557 400 577
rect 420 557 440 577
rect 460 557 480 577
rect 500 557 520 577
rect 540 557 560 577
rect 580 557 600 577
rect 620 557 640 577
rect 660 557 680 577
rect 700 557 720 577
rect 740 557 760 577
rect 780 557 800 577
rect 820 557 840 577
rect 860 557 880 577
rect 900 557 920 577
rect 940 557 960 577
rect 980 557 1000 577
rect 1020 557 1040 577
rect 1060 557 1080 577
rect 1100 557 1120 577
rect 1140 557 1160 577
rect 1180 557 1200 577
rect 1220 557 1240 577
rect 1260 557 1280 577
rect 1300 557 1320 577
rect 1340 557 1360 577
rect 1380 557 1400 577
rect 1420 557 1440 577
rect 1460 557 1480 577
rect 1500 557 1520 577
rect 1540 557 1560 577
rect 1580 557 1600 577
rect 1620 557 1640 577
rect 1660 557 1680 577
rect 1700 557 1720 577
rect 1740 557 1760 577
rect 1780 557 1800 577
rect 1820 557 1840 577
rect 1860 557 1880 577
rect 1900 557 1920 577
rect 1940 557 1960 577
rect 1980 557 2000 577
rect 2020 557 2040 577
rect 2060 557 2080 577
rect 2100 557 2120 577
rect 2140 557 2160 577
rect 2180 557 2200 577
rect 2220 557 2240 577
rect 2260 557 2280 577
rect 2300 557 2320 577
rect 2340 557 2360 577
rect 2380 557 2400 577
rect 2420 557 2440 577
rect 2460 557 2480 577
rect 2500 557 2520 577
rect 2540 557 2560 577
rect 2580 557 2600 577
rect 2620 557 2640 577
rect 2660 557 2675 577
rect 175 542 2675 557
rect 175 495 2675 510
rect 175 475 200 495
rect 220 475 240 495
rect 260 475 280 495
rect 300 475 320 495
rect 340 475 360 495
rect 380 475 400 495
rect 420 475 440 495
rect 460 475 480 495
rect 500 475 520 495
rect 540 475 560 495
rect 580 475 600 495
rect 620 475 640 495
rect 660 475 680 495
rect 700 475 720 495
rect 740 475 760 495
rect 780 475 800 495
rect 820 475 840 495
rect 860 475 880 495
rect 900 475 920 495
rect 940 475 960 495
rect 980 475 1000 495
rect 1020 475 1040 495
rect 1060 475 1080 495
rect 1100 475 1120 495
rect 1140 475 1160 495
rect 1180 475 1200 495
rect 1220 475 1240 495
rect 1260 475 1280 495
rect 1300 475 1320 495
rect 1340 475 1360 495
rect 1380 475 1400 495
rect 1420 475 1440 495
rect 1460 475 1480 495
rect 1500 475 1520 495
rect 1540 475 1560 495
rect 1580 475 1600 495
rect 1620 475 1640 495
rect 1660 475 1680 495
rect 1700 475 1720 495
rect 1740 475 1760 495
rect 1780 475 1800 495
rect 1820 475 1840 495
rect 1860 475 1880 495
rect 1900 475 1920 495
rect 1940 475 1960 495
rect 1980 475 2000 495
rect 2020 475 2040 495
rect 2060 475 2080 495
rect 2100 475 2120 495
rect 2140 475 2160 495
rect 2180 475 2200 495
rect 2220 475 2240 495
rect 2260 475 2280 495
rect 2300 475 2320 495
rect 2340 475 2360 495
rect 2380 475 2400 495
rect 2420 475 2440 495
rect 2460 475 2480 495
rect 2500 475 2520 495
rect 2540 475 2560 495
rect 2580 475 2600 495
rect 2620 475 2640 495
rect 2660 475 2675 495
rect 175 460 2675 475
rect 175 413 2675 428
rect 175 393 200 413
rect 220 393 240 413
rect 260 393 280 413
rect 300 393 320 413
rect 340 393 360 413
rect 380 393 400 413
rect 420 393 440 413
rect 460 393 480 413
rect 500 393 520 413
rect 540 393 560 413
rect 580 393 600 413
rect 620 393 640 413
rect 660 393 680 413
rect 700 393 720 413
rect 740 393 760 413
rect 780 393 800 413
rect 820 393 840 413
rect 860 393 880 413
rect 900 393 920 413
rect 940 393 960 413
rect 980 393 1000 413
rect 1020 393 1040 413
rect 1060 393 1080 413
rect 1100 393 1120 413
rect 1140 393 1160 413
rect 1180 393 1200 413
rect 1220 393 1240 413
rect 1260 393 1280 413
rect 1300 393 1320 413
rect 1340 393 1360 413
rect 1380 393 1400 413
rect 1420 393 1440 413
rect 1460 393 1480 413
rect 1500 393 1520 413
rect 1540 393 1560 413
rect 1580 393 1600 413
rect 1620 393 1640 413
rect 1660 393 1680 413
rect 1700 393 1720 413
rect 1740 393 1760 413
rect 1780 393 1800 413
rect 1820 393 1840 413
rect 1860 393 1880 413
rect 1900 393 1920 413
rect 1940 393 1960 413
rect 1980 393 2000 413
rect 2020 393 2040 413
rect 2060 393 2080 413
rect 2100 393 2120 413
rect 2140 393 2160 413
rect 2180 393 2200 413
rect 2220 393 2240 413
rect 2260 393 2280 413
rect 2300 393 2320 413
rect 2340 393 2360 413
rect 2380 393 2400 413
rect 2420 393 2440 413
rect 2460 393 2480 413
rect 2500 393 2520 413
rect 2540 393 2560 413
rect 2580 393 2600 413
rect 2620 393 2640 413
rect 2660 393 2675 413
rect 175 378 2675 393
rect 175 331 2675 346
rect 175 311 200 331
rect 220 311 240 331
rect 260 311 280 331
rect 300 311 320 331
rect 340 311 360 331
rect 380 311 400 331
rect 420 311 440 331
rect 460 311 480 331
rect 500 311 520 331
rect 540 311 560 331
rect 580 311 600 331
rect 620 311 640 331
rect 660 311 680 331
rect 700 311 720 331
rect 740 311 760 331
rect 780 311 800 331
rect 820 311 840 331
rect 860 311 880 331
rect 900 311 920 331
rect 940 311 960 331
rect 980 311 1000 331
rect 1020 311 1040 331
rect 1060 311 1080 331
rect 1100 311 1120 331
rect 1140 311 1160 331
rect 1180 311 1200 331
rect 1220 311 1240 331
rect 1260 311 1280 331
rect 1300 311 1320 331
rect 1340 311 1360 331
rect 1380 311 1400 331
rect 1420 311 1440 331
rect 1460 311 1480 331
rect 1500 311 1520 331
rect 1540 311 1560 331
rect 1580 311 1600 331
rect 1620 311 1640 331
rect 1660 311 1680 331
rect 1700 311 1720 331
rect 1740 311 1760 331
rect 1780 311 1800 331
rect 1820 311 1840 331
rect 1860 311 1880 331
rect 1900 311 1920 331
rect 1940 311 1960 331
rect 1980 311 2000 331
rect 2020 311 2040 331
rect 2060 311 2080 331
rect 2100 311 2120 331
rect 2140 311 2160 331
rect 2180 311 2200 331
rect 2220 311 2240 331
rect 2260 311 2280 331
rect 2300 311 2320 331
rect 2340 311 2360 331
rect 2380 311 2400 331
rect 2420 311 2440 331
rect 2460 311 2480 331
rect 2500 311 2520 331
rect 2540 311 2560 331
rect 2580 311 2600 331
rect 2620 311 2640 331
rect 2660 311 2675 331
rect 175 296 2675 311
rect 175 249 2675 264
rect 175 229 200 249
rect 220 229 240 249
rect 260 229 280 249
rect 300 229 320 249
rect 340 229 360 249
rect 380 229 400 249
rect 420 229 440 249
rect 460 229 480 249
rect 500 229 520 249
rect 540 229 560 249
rect 580 229 600 249
rect 620 229 640 249
rect 660 229 680 249
rect 700 229 720 249
rect 740 229 760 249
rect 780 229 800 249
rect 820 229 840 249
rect 860 229 880 249
rect 900 229 920 249
rect 940 229 960 249
rect 980 229 1000 249
rect 1020 229 1040 249
rect 1060 229 1080 249
rect 1100 229 1120 249
rect 1140 229 1160 249
rect 1180 229 1200 249
rect 1220 229 1240 249
rect 1260 229 1280 249
rect 1300 229 1320 249
rect 1340 229 1360 249
rect 1380 229 1400 249
rect 1420 229 1440 249
rect 1460 229 1480 249
rect 1500 229 1520 249
rect 1540 229 1560 249
rect 1580 229 1600 249
rect 1620 229 1640 249
rect 1660 229 1680 249
rect 1700 229 1720 249
rect 1740 229 1760 249
rect 1780 229 1800 249
rect 1820 229 1840 249
rect 1860 229 1880 249
rect 1900 229 1920 249
rect 1940 229 1960 249
rect 1980 229 2000 249
rect 2020 229 2040 249
rect 2060 229 2080 249
rect 2100 229 2120 249
rect 2140 229 2160 249
rect 2180 229 2200 249
rect 2220 229 2240 249
rect 2260 229 2280 249
rect 2300 229 2320 249
rect 2340 229 2360 249
rect 2380 229 2400 249
rect 2420 229 2440 249
rect 2460 229 2480 249
rect 2500 229 2520 249
rect 2540 229 2560 249
rect 2580 229 2600 249
rect 2620 229 2640 249
rect 2660 229 2675 249
rect 175 214 2675 229
rect 175 167 2675 182
rect 175 147 200 167
rect 220 147 240 167
rect 260 147 280 167
rect 300 147 320 167
rect 340 147 360 167
rect 380 147 400 167
rect 420 147 440 167
rect 460 147 480 167
rect 500 147 520 167
rect 540 147 560 167
rect 580 147 600 167
rect 620 147 640 167
rect 660 147 680 167
rect 700 147 720 167
rect 740 147 760 167
rect 780 147 800 167
rect 820 147 840 167
rect 860 147 880 167
rect 900 147 920 167
rect 940 147 960 167
rect 980 147 1000 167
rect 1020 147 1040 167
rect 1060 147 1080 167
rect 1100 147 1120 167
rect 1140 147 1160 167
rect 1180 147 1200 167
rect 1220 147 1240 167
rect 1260 147 1280 167
rect 1300 147 1320 167
rect 1340 147 1360 167
rect 1380 147 1400 167
rect 1420 147 1440 167
rect 1460 147 1480 167
rect 1500 147 1520 167
rect 1540 147 1560 167
rect 1580 147 1600 167
rect 1620 147 1640 167
rect 1660 147 1680 167
rect 1700 147 1720 167
rect 1740 147 1760 167
rect 1780 147 1800 167
rect 1820 147 1840 167
rect 1860 147 1880 167
rect 1900 147 1920 167
rect 1940 147 1960 167
rect 1980 147 2000 167
rect 2020 147 2040 167
rect 2060 147 2080 167
rect 2100 147 2120 167
rect 2140 147 2160 167
rect 2180 147 2200 167
rect 2220 147 2240 167
rect 2260 147 2280 167
rect 2300 147 2320 167
rect 2340 147 2360 167
rect 2380 147 2400 167
rect 2420 147 2440 167
rect 2460 147 2480 167
rect 2500 147 2520 167
rect 2540 147 2560 167
rect 2580 147 2600 167
rect 2620 147 2640 167
rect 2660 147 2675 167
rect 175 132 2675 147
rect 175 85 2675 100
rect 175 65 200 85
rect 220 65 240 85
rect 260 65 280 85
rect 300 65 320 85
rect 340 65 360 85
rect 380 65 400 85
rect 420 65 440 85
rect 460 65 480 85
rect 500 65 520 85
rect 540 65 560 85
rect 580 65 600 85
rect 620 65 640 85
rect 660 65 680 85
rect 700 65 720 85
rect 740 65 760 85
rect 780 65 800 85
rect 820 65 840 85
rect 860 65 880 85
rect 900 65 920 85
rect 940 65 960 85
rect 980 65 1000 85
rect 1020 65 1040 85
rect 1060 65 1080 85
rect 1100 65 1120 85
rect 1140 65 1160 85
rect 1180 65 1200 85
rect 1220 65 1240 85
rect 1260 65 1280 85
rect 1300 65 1320 85
rect 1340 65 1360 85
rect 1380 65 1400 85
rect 1420 65 1440 85
rect 1460 65 1480 85
rect 1500 65 1520 85
rect 1540 65 1560 85
rect 1580 65 1600 85
rect 1620 65 1640 85
rect 1660 65 1680 85
rect 1700 65 1720 85
rect 1740 65 1760 85
rect 1780 65 1800 85
rect 1820 65 1840 85
rect 1860 65 1880 85
rect 1900 65 1920 85
rect 1940 65 1960 85
rect 1980 65 2000 85
rect 2020 65 2040 85
rect 2060 65 2080 85
rect 2100 65 2120 85
rect 2140 65 2160 85
rect 2180 65 2200 85
rect 2220 65 2240 85
rect 2260 65 2280 85
rect 2300 65 2320 85
rect 2340 65 2360 85
rect 2380 65 2400 85
rect 2420 65 2440 85
rect 2460 65 2480 85
rect 2500 65 2520 85
rect 2540 65 2560 85
rect 2580 65 2600 85
rect 2620 65 2640 85
rect 2660 65 2675 85
rect 175 55 2675 65
rect 105 -215 2605 -205
rect 105 -235 120 -215
rect 140 -235 160 -215
rect 180 -235 200 -215
rect 220 -235 240 -215
rect 260 -235 280 -215
rect 300 -235 320 -215
rect 340 -235 360 -215
rect 380 -235 400 -215
rect 420 -235 440 -215
rect 460 -235 480 -215
rect 500 -235 520 -215
rect 540 -235 560 -215
rect 580 -235 600 -215
rect 620 -235 640 -215
rect 660 -235 680 -215
rect 700 -235 720 -215
rect 740 -235 760 -215
rect 780 -235 800 -215
rect 820 -235 840 -215
rect 860 -235 880 -215
rect 900 -235 920 -215
rect 940 -235 960 -215
rect 980 -235 1000 -215
rect 1020 -235 1040 -215
rect 1060 -235 1080 -215
rect 1100 -235 1120 -215
rect 1140 -235 1160 -215
rect 1180 -235 1200 -215
rect 1220 -235 1240 -215
rect 1260 -235 1280 -215
rect 1300 -235 1320 -215
rect 1340 -235 1360 -215
rect 1380 -235 1400 -215
rect 1420 -235 1440 -215
rect 1460 -235 1480 -215
rect 1500 -235 1520 -215
rect 1540 -235 1560 -215
rect 1580 -235 1600 -215
rect 1620 -235 1640 -215
rect 1660 -235 1680 -215
rect 1700 -235 1720 -215
rect 1740 -235 1760 -215
rect 1780 -235 1800 -215
rect 1820 -235 1840 -215
rect 1860 -235 1880 -215
rect 1900 -235 1920 -215
rect 1940 -235 1960 -215
rect 1980 -235 2000 -215
rect 2020 -235 2040 -215
rect 2060 -235 2080 -215
rect 2100 -235 2120 -215
rect 2140 -235 2160 -215
rect 2180 -235 2200 -215
rect 2220 -235 2240 -215
rect 2260 -235 2280 -215
rect 2300 -235 2320 -215
rect 2340 -235 2360 -215
rect 2380 -235 2400 -215
rect 2420 -235 2440 -215
rect 2460 -235 2480 -215
rect 2500 -235 2520 -215
rect 2540 -235 2560 -215
rect 2590 -235 2605 -215
rect 105 -250 2605 -235
rect 105 -310 2605 -295
rect 105 -330 120 -310
rect 140 -330 160 -310
rect 180 -330 200 -310
rect 220 -330 240 -310
rect 260 -330 280 -310
rect 300 -330 320 -310
rect 340 -330 360 -310
rect 380 -330 400 -310
rect 420 -330 440 -310
rect 460 -330 480 -310
rect 500 -330 520 -310
rect 540 -330 560 -310
rect 580 -330 600 -310
rect 620 -330 640 -310
rect 660 -330 680 -310
rect 700 -330 720 -310
rect 740 -330 760 -310
rect 780 -330 800 -310
rect 820 -330 840 -310
rect 860 -330 880 -310
rect 900 -330 920 -310
rect 940 -330 960 -310
rect 980 -330 1000 -310
rect 1020 -330 1040 -310
rect 1060 -330 1080 -310
rect 1100 -330 1120 -310
rect 1140 -330 1160 -310
rect 1180 -330 1200 -310
rect 1220 -330 1240 -310
rect 1260 -330 1280 -310
rect 1300 -330 1320 -310
rect 1340 -330 1360 -310
rect 1380 -330 1400 -310
rect 1420 -330 1440 -310
rect 1460 -330 1480 -310
rect 1500 -330 1520 -310
rect 1540 -330 1560 -310
rect 1580 -330 1600 -310
rect 1620 -330 1640 -310
rect 1660 -330 1680 -310
rect 1700 -330 1720 -310
rect 1740 -330 1760 -310
rect 1780 -330 1800 -310
rect 1820 -330 1840 -310
rect 1860 -330 1880 -310
rect 1900 -330 1920 -310
rect 1940 -330 1960 -310
rect 1980 -330 2000 -310
rect 2020 -330 2040 -310
rect 2060 -330 2080 -310
rect 2100 -330 2120 -310
rect 2140 -330 2160 -310
rect 2180 -330 2200 -310
rect 2220 -330 2240 -310
rect 2260 -330 2280 -310
rect 2300 -330 2320 -310
rect 2340 -330 2360 -310
rect 2380 -330 2400 -310
rect 2420 -330 2440 -310
rect 2460 -330 2480 -310
rect 2500 -330 2520 -310
rect 2540 -330 2560 -310
rect 2590 -330 2605 -310
rect 105 -345 2605 -330
rect 105 -405 2605 -390
rect 105 -425 120 -405
rect 140 -425 160 -405
rect 180 -425 200 -405
rect 220 -425 240 -405
rect 260 -425 280 -405
rect 300 -425 320 -405
rect 340 -425 360 -405
rect 380 -425 400 -405
rect 420 -425 440 -405
rect 460 -425 480 -405
rect 500 -425 520 -405
rect 540 -425 560 -405
rect 580 -425 600 -405
rect 620 -425 640 -405
rect 660 -425 680 -405
rect 700 -425 720 -405
rect 740 -425 760 -405
rect 780 -425 800 -405
rect 820 -425 840 -405
rect 860 -425 880 -405
rect 900 -425 920 -405
rect 940 -425 960 -405
rect 980 -425 1000 -405
rect 1020 -425 1040 -405
rect 1060 -425 1080 -405
rect 1100 -425 1120 -405
rect 1140 -425 1160 -405
rect 1180 -425 1200 -405
rect 1220 -425 1240 -405
rect 1260 -425 1280 -405
rect 1300 -425 1320 -405
rect 1340 -425 1360 -405
rect 1380 -425 1400 -405
rect 1420 -425 1440 -405
rect 1460 -425 1480 -405
rect 1500 -425 1520 -405
rect 1540 -425 1560 -405
rect 1580 -425 1600 -405
rect 1620 -425 1640 -405
rect 1660 -425 1680 -405
rect 1700 -425 1720 -405
rect 1740 -425 1760 -405
rect 1780 -425 1800 -405
rect 1820 -425 1840 -405
rect 1860 -425 1880 -405
rect 1900 -425 1920 -405
rect 1940 -425 1960 -405
rect 1980 -425 2000 -405
rect 2020 -425 2040 -405
rect 2060 -425 2080 -405
rect 2100 -425 2120 -405
rect 2140 -425 2160 -405
rect 2180 -425 2200 -405
rect 2220 -425 2240 -405
rect 2260 -425 2280 -405
rect 2300 -425 2320 -405
rect 2340 -425 2360 -405
rect 2380 -425 2400 -405
rect 2420 -425 2440 -405
rect 2460 -425 2480 -405
rect 2500 -425 2520 -405
rect 2540 -425 2560 -405
rect 2590 -425 2605 -405
rect 105 -440 2605 -425
rect 105 -500 2605 -485
rect 105 -520 120 -500
rect 140 -520 160 -500
rect 180 -520 200 -500
rect 220 -520 240 -500
rect 260 -520 280 -500
rect 300 -520 320 -500
rect 340 -520 360 -500
rect 380 -520 400 -500
rect 420 -520 440 -500
rect 460 -520 480 -500
rect 500 -520 520 -500
rect 540 -520 560 -500
rect 580 -520 600 -500
rect 620 -520 640 -500
rect 660 -520 680 -500
rect 700 -520 720 -500
rect 740 -520 760 -500
rect 780 -520 800 -500
rect 820 -520 840 -500
rect 860 -520 880 -500
rect 900 -520 920 -500
rect 940 -520 960 -500
rect 980 -520 1000 -500
rect 1020 -520 1040 -500
rect 1060 -520 1080 -500
rect 1100 -520 1120 -500
rect 1140 -520 1160 -500
rect 1180 -520 1200 -500
rect 1220 -520 1240 -500
rect 1260 -520 1280 -500
rect 1300 -520 1320 -500
rect 1340 -520 1360 -500
rect 1380 -520 1400 -500
rect 1420 -520 1440 -500
rect 1460 -520 1480 -500
rect 1500 -520 1520 -500
rect 1540 -520 1560 -500
rect 1580 -520 1600 -500
rect 1620 -520 1640 -500
rect 1660 -520 1680 -500
rect 1700 -520 1720 -500
rect 1740 -520 1760 -500
rect 1780 -520 1800 -500
rect 1820 -520 1840 -500
rect 1860 -520 1880 -500
rect 1900 -520 1920 -500
rect 1940 -520 1960 -500
rect 1980 -520 2000 -500
rect 2020 -520 2040 -500
rect 2060 -520 2080 -500
rect 2100 -520 2120 -500
rect 2140 -520 2160 -500
rect 2180 -520 2200 -500
rect 2220 -520 2240 -500
rect 2260 -520 2280 -500
rect 2300 -520 2320 -500
rect 2340 -520 2360 -500
rect 2380 -520 2400 -500
rect 2420 -520 2440 -500
rect 2460 -520 2480 -500
rect 2500 -520 2520 -500
rect 2540 -520 2560 -500
rect 2590 -520 2605 -500
rect 105 -535 2605 -520
rect 105 -595 2605 -580
rect 105 -615 120 -595
rect 140 -615 160 -595
rect 180 -615 200 -595
rect 220 -615 240 -595
rect 260 -615 280 -595
rect 300 -615 320 -595
rect 340 -615 360 -595
rect 380 -615 400 -595
rect 420 -615 440 -595
rect 460 -615 480 -595
rect 500 -615 520 -595
rect 540 -615 560 -595
rect 580 -615 600 -595
rect 620 -615 640 -595
rect 660 -615 680 -595
rect 700 -615 720 -595
rect 740 -615 760 -595
rect 780 -615 800 -595
rect 820 -615 840 -595
rect 860 -615 880 -595
rect 900 -615 920 -595
rect 940 -615 960 -595
rect 980 -615 1000 -595
rect 1020 -615 1040 -595
rect 1060 -615 1080 -595
rect 1100 -615 1120 -595
rect 1140 -615 1160 -595
rect 1180 -615 1200 -595
rect 1220 -615 1240 -595
rect 1260 -615 1280 -595
rect 1300 -615 1320 -595
rect 1340 -615 1360 -595
rect 1380 -615 1400 -595
rect 1420 -615 1440 -595
rect 1460 -615 1480 -595
rect 1500 -615 1520 -595
rect 1540 -615 1560 -595
rect 1580 -615 1600 -595
rect 1620 -615 1640 -595
rect 1660 -615 1680 -595
rect 1700 -615 1720 -595
rect 1740 -615 1760 -595
rect 1780 -615 1800 -595
rect 1820 -615 1840 -595
rect 1860 -615 1880 -595
rect 1900 -615 1920 -595
rect 1940 -615 1960 -595
rect 1980 -615 2000 -595
rect 2020 -615 2040 -595
rect 2060 -615 2080 -595
rect 2100 -615 2120 -595
rect 2140 -615 2160 -595
rect 2180 -615 2200 -595
rect 2220 -615 2240 -595
rect 2260 -615 2280 -595
rect 2300 -615 2320 -595
rect 2340 -615 2360 -595
rect 2380 -615 2400 -595
rect 2420 -615 2440 -595
rect 2460 -615 2480 -595
rect 2500 -615 2520 -595
rect 2540 -615 2560 -595
rect 2590 -615 2605 -595
rect 105 -630 2605 -615
rect 105 -690 2605 -675
rect 105 -710 120 -690
rect 140 -710 160 -690
rect 180 -710 200 -690
rect 220 -710 240 -690
rect 260 -710 280 -690
rect 300 -710 320 -690
rect 340 -710 360 -690
rect 380 -710 400 -690
rect 420 -710 440 -690
rect 460 -710 480 -690
rect 500 -710 520 -690
rect 540 -710 560 -690
rect 580 -710 600 -690
rect 620 -710 640 -690
rect 660 -710 680 -690
rect 700 -710 720 -690
rect 740 -710 760 -690
rect 780 -710 800 -690
rect 820 -710 840 -690
rect 860 -710 880 -690
rect 900 -710 920 -690
rect 940 -710 960 -690
rect 980 -710 1000 -690
rect 1020 -710 1040 -690
rect 1060 -710 1080 -690
rect 1100 -710 1120 -690
rect 1140 -710 1160 -690
rect 1180 -710 1200 -690
rect 1220 -710 1240 -690
rect 1260 -710 1280 -690
rect 1300 -710 1320 -690
rect 1340 -710 1360 -690
rect 1380 -710 1400 -690
rect 1420 -710 1440 -690
rect 1460 -710 1480 -690
rect 1500 -710 1520 -690
rect 1540 -710 1560 -690
rect 1580 -710 1600 -690
rect 1620 -710 1640 -690
rect 1660 -710 1680 -690
rect 1700 -710 1720 -690
rect 1740 -710 1760 -690
rect 1780 -710 1800 -690
rect 1820 -710 1840 -690
rect 1860 -710 1880 -690
rect 1900 -710 1920 -690
rect 1940 -710 1960 -690
rect 1980 -710 2000 -690
rect 2020 -710 2040 -690
rect 2060 -710 2080 -690
rect 2100 -710 2120 -690
rect 2140 -710 2160 -690
rect 2180 -710 2200 -690
rect 2220 -710 2240 -690
rect 2260 -710 2280 -690
rect 2300 -710 2320 -690
rect 2340 -710 2360 -690
rect 2380 -710 2400 -690
rect 2420 -710 2440 -690
rect 2460 -710 2480 -690
rect 2500 -710 2520 -690
rect 2540 -710 2560 -690
rect 2590 -710 2605 -690
rect 105 -725 2605 -710
rect 105 -785 2605 -770
rect 105 -805 120 -785
rect 140 -805 160 -785
rect 180 -805 200 -785
rect 220 -805 240 -785
rect 260 -805 280 -785
rect 300 -805 320 -785
rect 340 -805 360 -785
rect 380 -805 400 -785
rect 420 -805 440 -785
rect 460 -805 480 -785
rect 500 -805 520 -785
rect 540 -805 560 -785
rect 580 -805 600 -785
rect 620 -805 640 -785
rect 660 -805 680 -785
rect 700 -805 720 -785
rect 740 -805 760 -785
rect 780 -805 800 -785
rect 820 -805 840 -785
rect 860 -805 880 -785
rect 900 -805 920 -785
rect 940 -805 960 -785
rect 980 -805 1000 -785
rect 1020 -805 1040 -785
rect 1060 -805 1080 -785
rect 1100 -805 1120 -785
rect 1140 -805 1160 -785
rect 1180 -805 1200 -785
rect 1220 -805 1240 -785
rect 1260 -805 1280 -785
rect 1300 -805 1320 -785
rect 1340 -805 1360 -785
rect 1380 -805 1400 -785
rect 1420 -805 1440 -785
rect 1460 -805 1480 -785
rect 1500 -805 1520 -785
rect 1540 -805 1560 -785
rect 1580 -805 1600 -785
rect 1620 -805 1640 -785
rect 1660 -805 1680 -785
rect 1700 -805 1720 -785
rect 1740 -805 1760 -785
rect 1780 -805 1800 -785
rect 1820 -805 1840 -785
rect 1860 -805 1880 -785
rect 1900 -805 1920 -785
rect 1940 -805 1960 -785
rect 1980 -805 2000 -785
rect 2020 -805 2040 -785
rect 2060 -805 2080 -785
rect 2100 -805 2120 -785
rect 2140 -805 2160 -785
rect 2180 -805 2200 -785
rect 2220 -805 2240 -785
rect 2260 -805 2280 -785
rect 2300 -805 2320 -785
rect 2340 -805 2360 -785
rect 2380 -805 2400 -785
rect 2420 -805 2440 -785
rect 2460 -805 2480 -785
rect 2500 -805 2520 -785
rect 2540 -805 2560 -785
rect 2590 -805 2605 -785
rect 105 -820 2605 -805
rect 105 -880 2605 -865
rect 105 -900 120 -880
rect 140 -900 160 -880
rect 180 -900 200 -880
rect 220 -900 240 -880
rect 260 -900 280 -880
rect 300 -900 320 -880
rect 340 -900 360 -880
rect 380 -900 400 -880
rect 420 -900 440 -880
rect 460 -900 480 -880
rect 500 -900 520 -880
rect 540 -900 560 -880
rect 580 -900 600 -880
rect 620 -900 640 -880
rect 660 -900 680 -880
rect 700 -900 720 -880
rect 740 -900 760 -880
rect 780 -900 800 -880
rect 820 -900 840 -880
rect 860 -900 880 -880
rect 900 -900 920 -880
rect 940 -900 960 -880
rect 980 -900 1000 -880
rect 1020 -900 1040 -880
rect 1060 -900 1080 -880
rect 1100 -900 1120 -880
rect 1140 -900 1160 -880
rect 1180 -900 1200 -880
rect 1220 -900 1240 -880
rect 1260 -900 1280 -880
rect 1300 -900 1320 -880
rect 1340 -900 1360 -880
rect 1380 -900 1400 -880
rect 1420 -900 1440 -880
rect 1460 -900 1480 -880
rect 1500 -900 1520 -880
rect 1540 -900 1560 -880
rect 1580 -900 1600 -880
rect 1620 -900 1640 -880
rect 1660 -900 1680 -880
rect 1700 -900 1720 -880
rect 1740 -900 1760 -880
rect 1780 -900 1800 -880
rect 1820 -900 1840 -880
rect 1860 -900 1880 -880
rect 1900 -900 1920 -880
rect 1940 -900 1960 -880
rect 1980 -900 2000 -880
rect 2020 -900 2040 -880
rect 2060 -900 2080 -880
rect 2100 -900 2120 -880
rect 2140 -900 2160 -880
rect 2180 -900 2200 -880
rect 2220 -900 2240 -880
rect 2260 -900 2280 -880
rect 2300 -900 2320 -880
rect 2340 -900 2360 -880
rect 2380 -900 2400 -880
rect 2420 -900 2440 -880
rect 2460 -900 2480 -880
rect 2500 -900 2520 -880
rect 2540 -900 2560 -880
rect 2590 -900 2605 -880
rect 105 -915 2605 -900
rect 105 -975 2605 -960
rect 105 -995 120 -975
rect 140 -995 160 -975
rect 180 -995 200 -975
rect 220 -995 240 -975
rect 260 -995 280 -975
rect 300 -995 320 -975
rect 340 -995 360 -975
rect 380 -995 400 -975
rect 420 -995 440 -975
rect 460 -995 480 -975
rect 500 -995 520 -975
rect 540 -995 560 -975
rect 580 -995 600 -975
rect 620 -995 640 -975
rect 660 -995 680 -975
rect 700 -995 720 -975
rect 740 -995 760 -975
rect 780 -995 800 -975
rect 820 -995 840 -975
rect 860 -995 880 -975
rect 900 -995 920 -975
rect 940 -995 960 -975
rect 980 -995 1000 -975
rect 1020 -995 1040 -975
rect 1060 -995 1080 -975
rect 1100 -995 1120 -975
rect 1140 -995 1160 -975
rect 1180 -995 1200 -975
rect 1220 -995 1240 -975
rect 1260 -995 1280 -975
rect 1300 -995 1320 -975
rect 1340 -995 1360 -975
rect 1380 -995 1400 -975
rect 1420 -995 1440 -975
rect 1460 -995 1480 -975
rect 1500 -995 1520 -975
rect 1540 -995 1560 -975
rect 1580 -995 1600 -975
rect 1620 -995 1640 -975
rect 1660 -995 1680 -975
rect 1700 -995 1720 -975
rect 1740 -995 1760 -975
rect 1780 -995 1800 -975
rect 1820 -995 1840 -975
rect 1860 -995 1880 -975
rect 1900 -995 1920 -975
rect 1940 -995 1960 -975
rect 1980 -995 2000 -975
rect 2020 -995 2040 -975
rect 2060 -995 2080 -975
rect 2100 -995 2120 -975
rect 2140 -995 2160 -975
rect 2180 -995 2200 -975
rect 2220 -995 2240 -975
rect 2260 -995 2280 -975
rect 2300 -995 2320 -975
rect 2340 -995 2360 -975
rect 2380 -995 2400 -975
rect 2420 -995 2440 -975
rect 2460 -995 2480 -975
rect 2500 -995 2520 -975
rect 2540 -995 2560 -975
rect 2590 -995 2605 -975
rect 105 -1010 2605 -995
rect 105 -1070 2605 -1055
rect 105 -1090 120 -1070
rect 140 -1090 160 -1070
rect 180 -1090 200 -1070
rect 220 -1090 240 -1070
rect 260 -1090 280 -1070
rect 300 -1090 320 -1070
rect 340 -1090 360 -1070
rect 380 -1090 400 -1070
rect 420 -1090 440 -1070
rect 460 -1090 480 -1070
rect 500 -1090 520 -1070
rect 540 -1090 560 -1070
rect 580 -1090 600 -1070
rect 620 -1090 640 -1070
rect 660 -1090 680 -1070
rect 700 -1090 720 -1070
rect 740 -1090 760 -1070
rect 780 -1090 800 -1070
rect 820 -1090 840 -1070
rect 860 -1090 880 -1070
rect 900 -1090 920 -1070
rect 940 -1090 960 -1070
rect 980 -1090 1000 -1070
rect 1020 -1090 1040 -1070
rect 1060 -1090 1080 -1070
rect 1100 -1090 1120 -1070
rect 1140 -1090 1160 -1070
rect 1180 -1090 1200 -1070
rect 1220 -1090 1240 -1070
rect 1260 -1090 1280 -1070
rect 1300 -1090 1320 -1070
rect 1340 -1090 1360 -1070
rect 1380 -1090 1400 -1070
rect 1420 -1090 1440 -1070
rect 1460 -1090 1480 -1070
rect 1500 -1090 1520 -1070
rect 1540 -1090 1560 -1070
rect 1580 -1090 1600 -1070
rect 1620 -1090 1640 -1070
rect 1660 -1090 1680 -1070
rect 1700 -1090 1720 -1070
rect 1740 -1090 1760 -1070
rect 1780 -1090 1800 -1070
rect 1820 -1090 1840 -1070
rect 1860 -1090 1880 -1070
rect 1900 -1090 1920 -1070
rect 1940 -1090 1960 -1070
rect 1980 -1090 2000 -1070
rect 2020 -1090 2040 -1070
rect 2060 -1090 2080 -1070
rect 2100 -1090 2120 -1070
rect 2140 -1090 2160 -1070
rect 2180 -1090 2200 -1070
rect 2220 -1090 2240 -1070
rect 2260 -1090 2280 -1070
rect 2300 -1090 2320 -1070
rect 2340 -1090 2360 -1070
rect 2380 -1090 2400 -1070
rect 2420 -1090 2440 -1070
rect 2460 -1090 2480 -1070
rect 2500 -1090 2520 -1070
rect 2540 -1090 2560 -1070
rect 2590 -1090 2605 -1070
rect 105 -1105 2605 -1090
rect 105 -1165 2605 -1150
rect 105 -1185 120 -1165
rect 140 -1185 160 -1165
rect 180 -1185 200 -1165
rect 220 -1185 240 -1165
rect 260 -1185 280 -1165
rect 300 -1185 320 -1165
rect 340 -1185 360 -1165
rect 380 -1185 400 -1165
rect 420 -1185 440 -1165
rect 460 -1185 480 -1165
rect 500 -1185 520 -1165
rect 540 -1185 560 -1165
rect 580 -1185 600 -1165
rect 620 -1185 640 -1165
rect 660 -1185 680 -1165
rect 700 -1185 720 -1165
rect 740 -1185 760 -1165
rect 780 -1185 800 -1165
rect 820 -1185 840 -1165
rect 860 -1185 880 -1165
rect 900 -1185 920 -1165
rect 940 -1185 960 -1165
rect 980 -1185 1000 -1165
rect 1020 -1185 1040 -1165
rect 1060 -1185 1080 -1165
rect 1100 -1185 1120 -1165
rect 1140 -1185 1160 -1165
rect 1180 -1185 1200 -1165
rect 1220 -1185 1240 -1165
rect 1260 -1185 1280 -1165
rect 1300 -1185 1320 -1165
rect 1340 -1185 1360 -1165
rect 1380 -1185 1400 -1165
rect 1420 -1185 1440 -1165
rect 1460 -1185 1480 -1165
rect 1500 -1185 1520 -1165
rect 1540 -1185 1560 -1165
rect 1580 -1185 1600 -1165
rect 1620 -1185 1640 -1165
rect 1660 -1185 1680 -1165
rect 1700 -1185 1720 -1165
rect 1740 -1185 1760 -1165
rect 1780 -1185 1800 -1165
rect 1820 -1185 1840 -1165
rect 1860 -1185 1880 -1165
rect 1900 -1185 1920 -1165
rect 1940 -1185 1960 -1165
rect 1980 -1185 2000 -1165
rect 2020 -1185 2040 -1165
rect 2060 -1185 2080 -1165
rect 2100 -1185 2120 -1165
rect 2140 -1185 2160 -1165
rect 2180 -1185 2200 -1165
rect 2220 -1185 2240 -1165
rect 2260 -1185 2280 -1165
rect 2300 -1185 2320 -1165
rect 2340 -1185 2360 -1165
rect 2380 -1185 2400 -1165
rect 2420 -1185 2440 -1165
rect 2460 -1185 2480 -1165
rect 2500 -1185 2520 -1165
rect 2540 -1185 2560 -1165
rect 2590 -1185 2605 -1165
rect 105 -1200 2605 -1185
rect 105 -1260 2605 -1245
rect 105 -1280 120 -1260
rect 140 -1280 160 -1260
rect 180 -1280 200 -1260
rect 220 -1280 240 -1260
rect 260 -1280 280 -1260
rect 300 -1280 320 -1260
rect 340 -1280 360 -1260
rect 380 -1280 400 -1260
rect 420 -1280 440 -1260
rect 460 -1280 480 -1260
rect 500 -1280 520 -1260
rect 540 -1280 560 -1260
rect 580 -1280 600 -1260
rect 620 -1280 640 -1260
rect 660 -1280 680 -1260
rect 700 -1280 720 -1260
rect 740 -1280 760 -1260
rect 780 -1280 800 -1260
rect 820 -1280 840 -1260
rect 860 -1280 880 -1260
rect 900 -1280 920 -1260
rect 940 -1280 960 -1260
rect 980 -1280 1000 -1260
rect 1020 -1280 1040 -1260
rect 1060 -1280 1080 -1260
rect 1100 -1280 1120 -1260
rect 1140 -1280 1160 -1260
rect 1180 -1280 1200 -1260
rect 1220 -1280 1240 -1260
rect 1260 -1280 1280 -1260
rect 1300 -1280 1320 -1260
rect 1340 -1280 1360 -1260
rect 1380 -1280 1400 -1260
rect 1420 -1280 1440 -1260
rect 1460 -1280 1480 -1260
rect 1500 -1280 1520 -1260
rect 1540 -1280 1560 -1260
rect 1580 -1280 1600 -1260
rect 1620 -1280 1640 -1260
rect 1660 -1280 1680 -1260
rect 1700 -1280 1720 -1260
rect 1740 -1280 1760 -1260
rect 1780 -1280 1800 -1260
rect 1820 -1280 1840 -1260
rect 1860 -1280 1880 -1260
rect 1900 -1280 1920 -1260
rect 1940 -1280 1960 -1260
rect 1980 -1280 2000 -1260
rect 2020 -1280 2040 -1260
rect 2060 -1280 2080 -1260
rect 2100 -1280 2120 -1260
rect 2140 -1280 2160 -1260
rect 2180 -1280 2200 -1260
rect 2220 -1280 2240 -1260
rect 2260 -1280 2280 -1260
rect 2300 -1280 2320 -1260
rect 2340 -1280 2360 -1260
rect 2380 -1280 2400 -1260
rect 2420 -1280 2440 -1260
rect 2460 -1280 2480 -1260
rect 2500 -1280 2520 -1260
rect 2540 -1280 2560 -1260
rect 2590 -1280 2605 -1260
rect 105 -1295 2605 -1280
rect 105 -1355 2605 -1340
rect 105 -1375 120 -1355
rect 140 -1375 160 -1355
rect 180 -1375 200 -1355
rect 220 -1375 240 -1355
rect 260 -1375 280 -1355
rect 300 -1375 320 -1355
rect 340 -1375 360 -1355
rect 380 -1375 400 -1355
rect 420 -1375 440 -1355
rect 460 -1375 480 -1355
rect 500 -1375 520 -1355
rect 540 -1375 560 -1355
rect 580 -1375 600 -1355
rect 620 -1375 640 -1355
rect 660 -1375 680 -1355
rect 700 -1375 720 -1355
rect 740 -1375 760 -1355
rect 780 -1375 800 -1355
rect 820 -1375 840 -1355
rect 860 -1375 880 -1355
rect 900 -1375 920 -1355
rect 940 -1375 960 -1355
rect 980 -1375 1000 -1355
rect 1020 -1375 1040 -1355
rect 1060 -1375 1080 -1355
rect 1100 -1375 1120 -1355
rect 1140 -1375 1160 -1355
rect 1180 -1375 1200 -1355
rect 1220 -1375 1240 -1355
rect 1260 -1375 1280 -1355
rect 1300 -1375 1320 -1355
rect 1340 -1375 1360 -1355
rect 1380 -1375 1400 -1355
rect 1420 -1375 1440 -1355
rect 1460 -1375 1480 -1355
rect 1500 -1375 1520 -1355
rect 1540 -1375 1560 -1355
rect 1580 -1375 1600 -1355
rect 1620 -1375 1640 -1355
rect 1660 -1375 1680 -1355
rect 1700 -1375 1720 -1355
rect 1740 -1375 1760 -1355
rect 1780 -1375 1800 -1355
rect 1820 -1375 1840 -1355
rect 1860 -1375 1880 -1355
rect 1900 -1375 1920 -1355
rect 1940 -1375 1960 -1355
rect 1980 -1375 2000 -1355
rect 2020 -1375 2040 -1355
rect 2060 -1375 2080 -1355
rect 2100 -1375 2120 -1355
rect 2140 -1375 2160 -1355
rect 2180 -1375 2200 -1355
rect 2220 -1375 2240 -1355
rect 2260 -1375 2280 -1355
rect 2300 -1375 2320 -1355
rect 2340 -1375 2360 -1355
rect 2380 -1375 2400 -1355
rect 2420 -1375 2440 -1355
rect 2460 -1375 2480 -1355
rect 2500 -1375 2520 -1355
rect 2540 -1375 2560 -1355
rect 2590 -1375 2605 -1355
rect 105 -1390 2605 -1375
rect 105 -1450 2605 -1435
rect 105 -1470 120 -1450
rect 140 -1470 160 -1450
rect 180 -1470 200 -1450
rect 220 -1470 240 -1450
rect 260 -1470 280 -1450
rect 300 -1470 320 -1450
rect 340 -1470 360 -1450
rect 380 -1470 400 -1450
rect 420 -1470 440 -1450
rect 460 -1470 480 -1450
rect 500 -1470 520 -1450
rect 540 -1470 560 -1450
rect 580 -1470 600 -1450
rect 620 -1470 640 -1450
rect 660 -1470 680 -1450
rect 700 -1470 720 -1450
rect 740 -1470 760 -1450
rect 780 -1470 800 -1450
rect 820 -1470 840 -1450
rect 860 -1470 880 -1450
rect 900 -1470 920 -1450
rect 940 -1470 960 -1450
rect 980 -1470 1000 -1450
rect 1020 -1470 1040 -1450
rect 1060 -1470 1080 -1450
rect 1100 -1470 1120 -1450
rect 1140 -1470 1160 -1450
rect 1180 -1470 1200 -1450
rect 1220 -1470 1240 -1450
rect 1260 -1470 1280 -1450
rect 1300 -1470 1320 -1450
rect 1340 -1470 1360 -1450
rect 1380 -1470 1400 -1450
rect 1420 -1470 1440 -1450
rect 1460 -1470 1480 -1450
rect 1500 -1470 1520 -1450
rect 1540 -1470 1560 -1450
rect 1580 -1470 1600 -1450
rect 1620 -1470 1640 -1450
rect 1660 -1470 1680 -1450
rect 1700 -1470 1720 -1450
rect 1740 -1470 1760 -1450
rect 1780 -1470 1800 -1450
rect 1820 -1470 1840 -1450
rect 1860 -1470 1880 -1450
rect 1900 -1470 1920 -1450
rect 1940 -1470 1960 -1450
rect 1980 -1470 2000 -1450
rect 2020 -1470 2040 -1450
rect 2060 -1470 2080 -1450
rect 2100 -1470 2120 -1450
rect 2140 -1470 2160 -1450
rect 2180 -1470 2200 -1450
rect 2220 -1470 2240 -1450
rect 2260 -1470 2280 -1450
rect 2300 -1470 2320 -1450
rect 2340 -1470 2360 -1450
rect 2380 -1470 2400 -1450
rect 2420 -1470 2440 -1450
rect 2460 -1470 2480 -1450
rect 2500 -1470 2520 -1450
rect 2540 -1470 2560 -1450
rect 2590 -1470 2605 -1450
rect 105 -1485 2605 -1470
rect 105 -1545 2605 -1530
rect 105 -1565 120 -1545
rect 140 -1565 160 -1545
rect 180 -1565 200 -1545
rect 220 -1565 240 -1545
rect 260 -1565 280 -1545
rect 300 -1565 320 -1545
rect 340 -1565 360 -1545
rect 380 -1565 400 -1545
rect 420 -1565 440 -1545
rect 460 -1565 480 -1545
rect 500 -1565 520 -1545
rect 540 -1565 560 -1545
rect 580 -1565 600 -1545
rect 620 -1565 640 -1545
rect 660 -1565 680 -1545
rect 700 -1565 720 -1545
rect 740 -1565 760 -1545
rect 780 -1565 800 -1545
rect 820 -1565 840 -1545
rect 860 -1565 880 -1545
rect 900 -1565 920 -1545
rect 940 -1565 960 -1545
rect 980 -1565 1000 -1545
rect 1020 -1565 1040 -1545
rect 1060 -1565 1080 -1545
rect 1100 -1565 1120 -1545
rect 1140 -1565 1160 -1545
rect 1180 -1565 1200 -1545
rect 1220 -1565 1240 -1545
rect 1260 -1565 1280 -1545
rect 1300 -1565 1320 -1545
rect 1340 -1565 1360 -1545
rect 1380 -1565 1400 -1545
rect 1420 -1565 1440 -1545
rect 1460 -1565 1480 -1545
rect 1500 -1565 1520 -1545
rect 1540 -1565 1560 -1545
rect 1580 -1565 1600 -1545
rect 1620 -1565 1640 -1545
rect 1660 -1565 1680 -1545
rect 1700 -1565 1720 -1545
rect 1740 -1565 1760 -1545
rect 1780 -1565 1800 -1545
rect 1820 -1565 1840 -1545
rect 1860 -1565 1880 -1545
rect 1900 -1565 1920 -1545
rect 1940 -1565 1960 -1545
rect 1980 -1565 2000 -1545
rect 2020 -1565 2040 -1545
rect 2060 -1565 2080 -1545
rect 2100 -1565 2120 -1545
rect 2140 -1565 2160 -1545
rect 2180 -1565 2200 -1545
rect 2220 -1565 2240 -1545
rect 2260 -1565 2280 -1545
rect 2300 -1565 2320 -1545
rect 2340 -1565 2360 -1545
rect 2380 -1565 2400 -1545
rect 2420 -1565 2440 -1545
rect 2460 -1565 2480 -1545
rect 2500 -1565 2520 -1545
rect 2540 -1565 2560 -1545
rect 2590 -1565 2605 -1545
rect 105 -1580 2605 -1565
rect 105 -1640 2605 -1625
rect 105 -1660 120 -1640
rect 140 -1660 160 -1640
rect 180 -1660 200 -1640
rect 220 -1660 240 -1640
rect 260 -1660 280 -1640
rect 300 -1660 320 -1640
rect 340 -1660 360 -1640
rect 380 -1660 400 -1640
rect 420 -1660 440 -1640
rect 460 -1660 480 -1640
rect 500 -1660 520 -1640
rect 540 -1660 560 -1640
rect 580 -1660 600 -1640
rect 620 -1660 640 -1640
rect 660 -1660 680 -1640
rect 700 -1660 720 -1640
rect 740 -1660 760 -1640
rect 780 -1660 800 -1640
rect 820 -1660 840 -1640
rect 860 -1660 880 -1640
rect 900 -1660 920 -1640
rect 940 -1660 960 -1640
rect 980 -1660 1000 -1640
rect 1020 -1660 1040 -1640
rect 1060 -1660 1080 -1640
rect 1100 -1660 1120 -1640
rect 1140 -1660 1160 -1640
rect 1180 -1660 1200 -1640
rect 1220 -1660 1240 -1640
rect 1260 -1660 1280 -1640
rect 1300 -1660 1320 -1640
rect 1340 -1660 1360 -1640
rect 1380 -1660 1400 -1640
rect 1420 -1660 1440 -1640
rect 1460 -1660 1480 -1640
rect 1500 -1660 1520 -1640
rect 1540 -1660 1560 -1640
rect 1580 -1660 1600 -1640
rect 1620 -1660 1640 -1640
rect 1660 -1660 1680 -1640
rect 1700 -1660 1720 -1640
rect 1740 -1660 1760 -1640
rect 1780 -1660 1800 -1640
rect 1820 -1660 1840 -1640
rect 1860 -1660 1880 -1640
rect 1900 -1660 1920 -1640
rect 1940 -1660 1960 -1640
rect 1980 -1660 2000 -1640
rect 2020 -1660 2040 -1640
rect 2060 -1660 2080 -1640
rect 2100 -1660 2120 -1640
rect 2140 -1660 2160 -1640
rect 2180 -1660 2200 -1640
rect 2220 -1660 2240 -1640
rect 2260 -1660 2280 -1640
rect 2300 -1660 2320 -1640
rect 2340 -1660 2360 -1640
rect 2380 -1660 2400 -1640
rect 2420 -1660 2440 -1640
rect 2460 -1660 2480 -1640
rect 2500 -1660 2520 -1640
rect 2540 -1660 2560 -1640
rect 2590 -1660 2605 -1640
rect 105 -1675 2605 -1660
rect 105 -1735 2605 -1720
rect 105 -1755 120 -1735
rect 140 -1755 160 -1735
rect 180 -1755 200 -1735
rect 220 -1755 240 -1735
rect 260 -1755 280 -1735
rect 300 -1755 320 -1735
rect 340 -1755 360 -1735
rect 380 -1755 400 -1735
rect 420 -1755 440 -1735
rect 460 -1755 480 -1735
rect 500 -1755 520 -1735
rect 540 -1755 560 -1735
rect 580 -1755 600 -1735
rect 620 -1755 640 -1735
rect 660 -1755 680 -1735
rect 700 -1755 720 -1735
rect 740 -1755 760 -1735
rect 780 -1755 800 -1735
rect 820 -1755 840 -1735
rect 860 -1755 880 -1735
rect 900 -1755 920 -1735
rect 940 -1755 960 -1735
rect 980 -1755 1000 -1735
rect 1020 -1755 1040 -1735
rect 1060 -1755 1080 -1735
rect 1100 -1755 1120 -1735
rect 1140 -1755 1160 -1735
rect 1180 -1755 1200 -1735
rect 1220 -1755 1240 -1735
rect 1260 -1755 1280 -1735
rect 1300 -1755 1320 -1735
rect 1340 -1755 1360 -1735
rect 1380 -1755 1400 -1735
rect 1420 -1755 1440 -1735
rect 1460 -1755 1480 -1735
rect 1500 -1755 1520 -1735
rect 1540 -1755 1560 -1735
rect 1580 -1755 1600 -1735
rect 1620 -1755 1640 -1735
rect 1660 -1755 1680 -1735
rect 1700 -1755 1720 -1735
rect 1740 -1755 1760 -1735
rect 1780 -1755 1800 -1735
rect 1820 -1755 1840 -1735
rect 1860 -1755 1880 -1735
rect 1900 -1755 1920 -1735
rect 1940 -1755 1960 -1735
rect 1980 -1755 2000 -1735
rect 2020 -1755 2040 -1735
rect 2060 -1755 2080 -1735
rect 2100 -1755 2120 -1735
rect 2140 -1755 2160 -1735
rect 2180 -1755 2200 -1735
rect 2220 -1755 2240 -1735
rect 2260 -1755 2280 -1735
rect 2300 -1755 2320 -1735
rect 2340 -1755 2360 -1735
rect 2380 -1755 2400 -1735
rect 2420 -1755 2440 -1735
rect 2460 -1755 2480 -1735
rect 2500 -1755 2520 -1735
rect 2540 -1755 2560 -1735
rect 2590 -1755 2605 -1735
rect 105 -1770 2605 -1755
rect 105 -1830 2605 -1815
rect 105 -1850 120 -1830
rect 140 -1850 160 -1830
rect 180 -1850 200 -1830
rect 220 -1850 240 -1830
rect 260 -1850 280 -1830
rect 300 -1850 320 -1830
rect 340 -1850 360 -1830
rect 380 -1850 400 -1830
rect 420 -1850 440 -1830
rect 460 -1850 480 -1830
rect 500 -1850 520 -1830
rect 540 -1850 560 -1830
rect 580 -1850 600 -1830
rect 620 -1850 640 -1830
rect 660 -1850 680 -1830
rect 700 -1850 720 -1830
rect 740 -1850 760 -1830
rect 780 -1850 800 -1830
rect 820 -1850 840 -1830
rect 860 -1850 880 -1830
rect 900 -1850 920 -1830
rect 940 -1850 960 -1830
rect 980 -1850 1000 -1830
rect 1020 -1850 1040 -1830
rect 1060 -1850 1080 -1830
rect 1100 -1850 1120 -1830
rect 1140 -1850 1160 -1830
rect 1180 -1850 1200 -1830
rect 1220 -1850 1240 -1830
rect 1260 -1850 1280 -1830
rect 1300 -1850 1320 -1830
rect 1340 -1850 1360 -1830
rect 1380 -1850 1400 -1830
rect 1420 -1850 1440 -1830
rect 1460 -1850 1480 -1830
rect 1500 -1850 1520 -1830
rect 1540 -1850 1560 -1830
rect 1580 -1850 1600 -1830
rect 1620 -1850 1640 -1830
rect 1660 -1850 1680 -1830
rect 1700 -1850 1720 -1830
rect 1740 -1850 1760 -1830
rect 1780 -1850 1800 -1830
rect 1820 -1850 1840 -1830
rect 1860 -1850 1880 -1830
rect 1900 -1850 1920 -1830
rect 1940 -1850 1960 -1830
rect 1980 -1850 2000 -1830
rect 2020 -1850 2040 -1830
rect 2060 -1850 2080 -1830
rect 2100 -1850 2120 -1830
rect 2140 -1850 2160 -1830
rect 2180 -1850 2200 -1830
rect 2220 -1850 2240 -1830
rect 2260 -1850 2280 -1830
rect 2300 -1850 2320 -1830
rect 2340 -1850 2360 -1830
rect 2380 -1850 2400 -1830
rect 2420 -1850 2440 -1830
rect 2460 -1850 2480 -1830
rect 2500 -1850 2520 -1830
rect 2540 -1850 2560 -1830
rect 2590 -1850 2605 -1830
rect 105 -1865 2605 -1850
rect 105 -1925 2605 -1910
rect 105 -1945 120 -1925
rect 140 -1945 160 -1925
rect 180 -1945 200 -1925
rect 220 -1945 240 -1925
rect 260 -1945 280 -1925
rect 300 -1945 320 -1925
rect 340 -1945 360 -1925
rect 380 -1945 400 -1925
rect 420 -1945 440 -1925
rect 460 -1945 480 -1925
rect 500 -1945 520 -1925
rect 540 -1945 560 -1925
rect 580 -1945 600 -1925
rect 620 -1945 640 -1925
rect 660 -1945 680 -1925
rect 700 -1945 720 -1925
rect 740 -1945 760 -1925
rect 780 -1945 800 -1925
rect 820 -1945 840 -1925
rect 860 -1945 880 -1925
rect 900 -1945 920 -1925
rect 940 -1945 960 -1925
rect 980 -1945 1000 -1925
rect 1020 -1945 1040 -1925
rect 1060 -1945 1080 -1925
rect 1100 -1945 1120 -1925
rect 1140 -1945 1160 -1925
rect 1180 -1945 1200 -1925
rect 1220 -1945 1240 -1925
rect 1260 -1945 1280 -1925
rect 1300 -1945 1320 -1925
rect 1340 -1945 1360 -1925
rect 1380 -1945 1400 -1925
rect 1420 -1945 1440 -1925
rect 1460 -1945 1480 -1925
rect 1500 -1945 1520 -1925
rect 1540 -1945 1560 -1925
rect 1580 -1945 1600 -1925
rect 1620 -1945 1640 -1925
rect 1660 -1945 1680 -1925
rect 1700 -1945 1720 -1925
rect 1740 -1945 1760 -1925
rect 1780 -1945 1800 -1925
rect 1820 -1945 1840 -1925
rect 1860 -1945 1880 -1925
rect 1900 -1945 1920 -1925
rect 1940 -1945 1960 -1925
rect 1980 -1945 2000 -1925
rect 2020 -1945 2040 -1925
rect 2060 -1945 2080 -1925
rect 2100 -1945 2120 -1925
rect 2140 -1945 2160 -1925
rect 2180 -1945 2200 -1925
rect 2220 -1945 2240 -1925
rect 2260 -1945 2280 -1925
rect 2300 -1945 2320 -1925
rect 2340 -1945 2360 -1925
rect 2380 -1945 2400 -1925
rect 2420 -1945 2440 -1925
rect 2460 -1945 2480 -1925
rect 2500 -1945 2520 -1925
rect 2540 -1945 2560 -1925
rect 2590 -1945 2605 -1925
rect 105 -1960 2605 -1945
rect 105 -2020 2605 -2005
rect 105 -2040 120 -2020
rect 140 -2040 160 -2020
rect 180 -2040 200 -2020
rect 220 -2040 240 -2020
rect 260 -2040 280 -2020
rect 300 -2040 320 -2020
rect 340 -2040 360 -2020
rect 380 -2040 400 -2020
rect 420 -2040 440 -2020
rect 460 -2040 480 -2020
rect 500 -2040 520 -2020
rect 540 -2040 560 -2020
rect 580 -2040 600 -2020
rect 620 -2040 640 -2020
rect 660 -2040 680 -2020
rect 700 -2040 720 -2020
rect 740 -2040 760 -2020
rect 780 -2040 800 -2020
rect 820 -2040 840 -2020
rect 860 -2040 880 -2020
rect 900 -2040 920 -2020
rect 940 -2040 960 -2020
rect 980 -2040 1000 -2020
rect 1020 -2040 1040 -2020
rect 1060 -2040 1080 -2020
rect 1100 -2040 1120 -2020
rect 1140 -2040 1160 -2020
rect 1180 -2040 1200 -2020
rect 1220 -2040 1240 -2020
rect 1260 -2040 1280 -2020
rect 1300 -2040 1320 -2020
rect 1340 -2040 1360 -2020
rect 1380 -2040 1400 -2020
rect 1420 -2040 1440 -2020
rect 1460 -2040 1480 -2020
rect 1500 -2040 1520 -2020
rect 1540 -2040 1560 -2020
rect 1580 -2040 1600 -2020
rect 1620 -2040 1640 -2020
rect 1660 -2040 1680 -2020
rect 1700 -2040 1720 -2020
rect 1740 -2040 1760 -2020
rect 1780 -2040 1800 -2020
rect 1820 -2040 1840 -2020
rect 1860 -2040 1880 -2020
rect 1900 -2040 1920 -2020
rect 1940 -2040 1960 -2020
rect 1980 -2040 2000 -2020
rect 2020 -2040 2040 -2020
rect 2060 -2040 2080 -2020
rect 2100 -2040 2120 -2020
rect 2140 -2040 2160 -2020
rect 2180 -2040 2200 -2020
rect 2220 -2040 2240 -2020
rect 2260 -2040 2280 -2020
rect 2300 -2040 2320 -2020
rect 2340 -2040 2360 -2020
rect 2380 -2040 2400 -2020
rect 2420 -2040 2440 -2020
rect 2460 -2040 2480 -2020
rect 2500 -2040 2520 -2020
rect 2540 -2040 2560 -2020
rect 2590 -2040 2605 -2020
rect 105 -2055 2605 -2040
rect 105 -2115 2605 -2100
rect 105 -2135 120 -2115
rect 140 -2135 160 -2115
rect 180 -2135 200 -2115
rect 220 -2135 240 -2115
rect 260 -2135 280 -2115
rect 300 -2135 320 -2115
rect 340 -2135 360 -2115
rect 380 -2135 400 -2115
rect 420 -2135 440 -2115
rect 460 -2135 480 -2115
rect 500 -2135 520 -2115
rect 540 -2135 560 -2115
rect 580 -2135 600 -2115
rect 620 -2135 640 -2115
rect 660 -2135 680 -2115
rect 700 -2135 720 -2115
rect 740 -2135 760 -2115
rect 780 -2135 800 -2115
rect 820 -2135 840 -2115
rect 860 -2135 880 -2115
rect 900 -2135 920 -2115
rect 940 -2135 960 -2115
rect 980 -2135 1000 -2115
rect 1020 -2135 1040 -2115
rect 1060 -2135 1080 -2115
rect 1100 -2135 1120 -2115
rect 1140 -2135 1160 -2115
rect 1180 -2135 1200 -2115
rect 1220 -2135 1240 -2115
rect 1260 -2135 1280 -2115
rect 1300 -2135 1320 -2115
rect 1340 -2135 1360 -2115
rect 1380 -2135 1400 -2115
rect 1420 -2135 1440 -2115
rect 1460 -2135 1480 -2115
rect 1500 -2135 1520 -2115
rect 1540 -2135 1560 -2115
rect 1580 -2135 1600 -2115
rect 1620 -2135 1640 -2115
rect 1660 -2135 1680 -2115
rect 1700 -2135 1720 -2115
rect 1740 -2135 1760 -2115
rect 1780 -2135 1800 -2115
rect 1820 -2135 1840 -2115
rect 1860 -2135 1880 -2115
rect 1900 -2135 1920 -2115
rect 1940 -2135 1960 -2115
rect 1980 -2135 2000 -2115
rect 2020 -2135 2040 -2115
rect 2060 -2135 2080 -2115
rect 2100 -2135 2120 -2115
rect 2140 -2135 2160 -2115
rect 2180 -2135 2200 -2115
rect 2220 -2135 2240 -2115
rect 2260 -2135 2280 -2115
rect 2300 -2135 2320 -2115
rect 2340 -2135 2360 -2115
rect 2380 -2135 2400 -2115
rect 2420 -2135 2440 -2115
rect 2460 -2135 2480 -2115
rect 2500 -2135 2520 -2115
rect 2540 -2135 2560 -2115
rect 2590 -2135 2605 -2115
rect 105 -2150 2605 -2135
rect 105 -2210 2605 -2195
rect 105 -2230 120 -2210
rect 140 -2230 160 -2210
rect 180 -2230 200 -2210
rect 220 -2230 240 -2210
rect 260 -2230 280 -2210
rect 300 -2230 320 -2210
rect 340 -2230 360 -2210
rect 380 -2230 400 -2210
rect 420 -2230 440 -2210
rect 460 -2230 480 -2210
rect 500 -2230 520 -2210
rect 540 -2230 560 -2210
rect 580 -2230 600 -2210
rect 620 -2230 640 -2210
rect 660 -2230 680 -2210
rect 700 -2230 720 -2210
rect 740 -2230 760 -2210
rect 780 -2230 800 -2210
rect 820 -2230 840 -2210
rect 860 -2230 880 -2210
rect 900 -2230 920 -2210
rect 940 -2230 960 -2210
rect 980 -2230 1000 -2210
rect 1020 -2230 1040 -2210
rect 1060 -2230 1080 -2210
rect 1100 -2230 1120 -2210
rect 1140 -2230 1160 -2210
rect 1180 -2230 1200 -2210
rect 1220 -2230 1240 -2210
rect 1260 -2230 1280 -2210
rect 1300 -2230 1320 -2210
rect 1340 -2230 1360 -2210
rect 1380 -2230 1400 -2210
rect 1420 -2230 1440 -2210
rect 1460 -2230 1480 -2210
rect 1500 -2230 1520 -2210
rect 1540 -2230 1560 -2210
rect 1580 -2230 1600 -2210
rect 1620 -2230 1640 -2210
rect 1660 -2230 1680 -2210
rect 1700 -2230 1720 -2210
rect 1740 -2230 1760 -2210
rect 1780 -2230 1800 -2210
rect 1820 -2230 1840 -2210
rect 1860 -2230 1880 -2210
rect 1900 -2230 1920 -2210
rect 1940 -2230 1960 -2210
rect 1980 -2230 2000 -2210
rect 2020 -2230 2040 -2210
rect 2060 -2230 2080 -2210
rect 2100 -2230 2120 -2210
rect 2140 -2230 2160 -2210
rect 2180 -2230 2200 -2210
rect 2220 -2230 2240 -2210
rect 2260 -2230 2280 -2210
rect 2300 -2230 2320 -2210
rect 2340 -2230 2360 -2210
rect 2380 -2230 2400 -2210
rect 2420 -2230 2440 -2210
rect 2460 -2230 2480 -2210
rect 2500 -2230 2520 -2210
rect 2540 -2230 2560 -2210
rect 2590 -2230 2605 -2210
rect 105 -2245 2605 -2230
rect 105 -2305 2605 -2290
rect 105 -2325 120 -2305
rect 140 -2325 160 -2305
rect 180 -2325 200 -2305
rect 220 -2325 240 -2305
rect 260 -2325 280 -2305
rect 300 -2325 320 -2305
rect 340 -2325 360 -2305
rect 380 -2325 400 -2305
rect 420 -2325 440 -2305
rect 460 -2325 480 -2305
rect 500 -2325 520 -2305
rect 540 -2325 560 -2305
rect 580 -2325 600 -2305
rect 620 -2325 640 -2305
rect 660 -2325 680 -2305
rect 700 -2325 720 -2305
rect 740 -2325 760 -2305
rect 780 -2325 800 -2305
rect 820 -2325 840 -2305
rect 860 -2325 880 -2305
rect 900 -2325 920 -2305
rect 940 -2325 960 -2305
rect 980 -2325 1000 -2305
rect 1020 -2325 1040 -2305
rect 1060 -2325 1080 -2305
rect 1100 -2325 1120 -2305
rect 1140 -2325 1160 -2305
rect 1180 -2325 1200 -2305
rect 1220 -2325 1240 -2305
rect 1260 -2325 1280 -2305
rect 1300 -2325 1320 -2305
rect 1340 -2325 1360 -2305
rect 1380 -2325 1400 -2305
rect 1420 -2325 1440 -2305
rect 1460 -2325 1480 -2305
rect 1500 -2325 1520 -2305
rect 1540 -2325 1560 -2305
rect 1580 -2325 1600 -2305
rect 1620 -2325 1640 -2305
rect 1660 -2325 1680 -2305
rect 1700 -2325 1720 -2305
rect 1740 -2325 1760 -2305
rect 1780 -2325 1800 -2305
rect 1820 -2325 1840 -2305
rect 1860 -2325 1880 -2305
rect 1900 -2325 1920 -2305
rect 1940 -2325 1960 -2305
rect 1980 -2325 2000 -2305
rect 2020 -2325 2040 -2305
rect 2060 -2325 2080 -2305
rect 2100 -2325 2120 -2305
rect 2140 -2325 2160 -2305
rect 2180 -2325 2200 -2305
rect 2220 -2325 2240 -2305
rect 2260 -2325 2280 -2305
rect 2300 -2325 2320 -2305
rect 2340 -2325 2360 -2305
rect 2380 -2325 2400 -2305
rect 2420 -2325 2440 -2305
rect 2460 -2325 2480 -2305
rect 2500 -2325 2520 -2305
rect 2540 -2325 2560 -2305
rect 2590 -2325 2605 -2305
rect 105 -2340 2605 -2325
rect 105 -2400 2605 -2385
rect 105 -2420 120 -2400
rect 140 -2420 160 -2400
rect 180 -2420 200 -2400
rect 220 -2420 240 -2400
rect 260 -2420 280 -2400
rect 300 -2420 320 -2400
rect 340 -2420 360 -2400
rect 380 -2420 400 -2400
rect 420 -2420 440 -2400
rect 460 -2420 480 -2400
rect 500 -2420 520 -2400
rect 540 -2420 560 -2400
rect 580 -2420 600 -2400
rect 620 -2420 640 -2400
rect 660 -2420 680 -2400
rect 700 -2420 720 -2400
rect 740 -2420 760 -2400
rect 780 -2420 800 -2400
rect 820 -2420 840 -2400
rect 860 -2420 880 -2400
rect 900 -2420 920 -2400
rect 940 -2420 960 -2400
rect 980 -2420 1000 -2400
rect 1020 -2420 1040 -2400
rect 1060 -2420 1080 -2400
rect 1100 -2420 1120 -2400
rect 1140 -2420 1160 -2400
rect 1180 -2420 1200 -2400
rect 1220 -2420 1240 -2400
rect 1260 -2420 1280 -2400
rect 1300 -2420 1320 -2400
rect 1340 -2420 1360 -2400
rect 1380 -2420 1400 -2400
rect 1420 -2420 1440 -2400
rect 1460 -2420 1480 -2400
rect 1500 -2420 1520 -2400
rect 1540 -2420 1560 -2400
rect 1580 -2420 1600 -2400
rect 1620 -2420 1640 -2400
rect 1660 -2420 1680 -2400
rect 1700 -2420 1720 -2400
rect 1740 -2420 1760 -2400
rect 1780 -2420 1800 -2400
rect 1820 -2420 1840 -2400
rect 1860 -2420 1880 -2400
rect 1900 -2420 1920 -2400
rect 1940 -2420 1960 -2400
rect 1980 -2420 2000 -2400
rect 2020 -2420 2040 -2400
rect 2060 -2420 2080 -2400
rect 2100 -2420 2120 -2400
rect 2140 -2420 2160 -2400
rect 2180 -2420 2200 -2400
rect 2220 -2420 2240 -2400
rect 2260 -2420 2280 -2400
rect 2300 -2420 2320 -2400
rect 2340 -2420 2360 -2400
rect 2380 -2420 2400 -2400
rect 2420 -2420 2440 -2400
rect 2460 -2420 2480 -2400
rect 2500 -2420 2520 -2400
rect 2540 -2420 2560 -2400
rect 2590 -2420 2605 -2400
rect 105 -2435 2605 -2420
rect 105 -2495 2605 -2480
rect 105 -2515 120 -2495
rect 140 -2515 160 -2495
rect 180 -2515 200 -2495
rect 220 -2515 240 -2495
rect 260 -2515 280 -2495
rect 300 -2515 320 -2495
rect 340 -2515 360 -2495
rect 380 -2515 400 -2495
rect 420 -2515 440 -2495
rect 460 -2515 480 -2495
rect 500 -2515 520 -2495
rect 540 -2515 560 -2495
rect 580 -2515 600 -2495
rect 620 -2515 640 -2495
rect 660 -2515 680 -2495
rect 700 -2515 720 -2495
rect 740 -2515 760 -2495
rect 780 -2515 800 -2495
rect 820 -2515 840 -2495
rect 860 -2515 880 -2495
rect 900 -2515 920 -2495
rect 940 -2515 960 -2495
rect 980 -2515 1000 -2495
rect 1020 -2515 1040 -2495
rect 1060 -2515 1080 -2495
rect 1100 -2515 1120 -2495
rect 1140 -2515 1160 -2495
rect 1180 -2515 1200 -2495
rect 1220 -2515 1240 -2495
rect 1260 -2515 1280 -2495
rect 1300 -2515 1320 -2495
rect 1340 -2515 1360 -2495
rect 1380 -2515 1400 -2495
rect 1420 -2515 1440 -2495
rect 1460 -2515 1480 -2495
rect 1500 -2515 1520 -2495
rect 1540 -2515 1560 -2495
rect 1580 -2515 1600 -2495
rect 1620 -2515 1640 -2495
rect 1660 -2515 1680 -2495
rect 1700 -2515 1720 -2495
rect 1740 -2515 1760 -2495
rect 1780 -2515 1800 -2495
rect 1820 -2515 1840 -2495
rect 1860 -2515 1880 -2495
rect 1900 -2515 1920 -2495
rect 1940 -2515 1960 -2495
rect 1980 -2515 2000 -2495
rect 2020 -2515 2040 -2495
rect 2060 -2515 2080 -2495
rect 2100 -2515 2120 -2495
rect 2140 -2515 2160 -2495
rect 2180 -2515 2200 -2495
rect 2220 -2515 2240 -2495
rect 2260 -2515 2280 -2495
rect 2300 -2515 2320 -2495
rect 2340 -2515 2360 -2495
rect 2380 -2515 2400 -2495
rect 2420 -2515 2440 -2495
rect 2460 -2515 2480 -2495
rect 2500 -2515 2520 -2495
rect 2540 -2515 2560 -2495
rect 2590 -2515 2605 -2495
rect 105 -2530 2605 -2515
rect 105 -2590 2605 -2575
rect 105 -2610 120 -2590
rect 140 -2610 160 -2590
rect 180 -2610 200 -2590
rect 220 -2610 240 -2590
rect 260 -2610 280 -2590
rect 300 -2610 320 -2590
rect 340 -2610 360 -2590
rect 380 -2610 400 -2590
rect 420 -2610 440 -2590
rect 460 -2610 480 -2590
rect 500 -2610 520 -2590
rect 540 -2610 560 -2590
rect 580 -2610 600 -2590
rect 620 -2610 640 -2590
rect 660 -2610 680 -2590
rect 700 -2610 720 -2590
rect 740 -2610 760 -2590
rect 780 -2610 800 -2590
rect 820 -2610 840 -2590
rect 860 -2610 880 -2590
rect 900 -2610 920 -2590
rect 940 -2610 960 -2590
rect 980 -2610 1000 -2590
rect 1020 -2610 1040 -2590
rect 1060 -2610 1080 -2590
rect 1100 -2610 1120 -2590
rect 1140 -2610 1160 -2590
rect 1180 -2610 1200 -2590
rect 1220 -2610 1240 -2590
rect 1260 -2610 1280 -2590
rect 1300 -2610 1320 -2590
rect 1340 -2610 1360 -2590
rect 1380 -2610 1400 -2590
rect 1420 -2610 1440 -2590
rect 1460 -2610 1480 -2590
rect 1500 -2610 1520 -2590
rect 1540 -2610 1560 -2590
rect 1580 -2610 1600 -2590
rect 1620 -2610 1640 -2590
rect 1660 -2610 1680 -2590
rect 1700 -2610 1720 -2590
rect 1740 -2610 1760 -2590
rect 1780 -2610 1800 -2590
rect 1820 -2610 1840 -2590
rect 1860 -2610 1880 -2590
rect 1900 -2610 1920 -2590
rect 1940 -2610 1960 -2590
rect 1980 -2610 2000 -2590
rect 2020 -2610 2040 -2590
rect 2060 -2610 2080 -2590
rect 2100 -2610 2120 -2590
rect 2140 -2610 2160 -2590
rect 2180 -2610 2200 -2590
rect 2220 -2610 2240 -2590
rect 2260 -2610 2280 -2590
rect 2300 -2610 2320 -2590
rect 2340 -2610 2360 -2590
rect 2380 -2610 2400 -2590
rect 2420 -2610 2440 -2590
rect 2460 -2610 2480 -2590
rect 2500 -2610 2520 -2590
rect 2540 -2610 2560 -2590
rect 2590 -2610 2605 -2590
rect 105 -2625 2605 -2610
rect 105 -2685 2605 -2670
rect 105 -2705 120 -2685
rect 140 -2705 160 -2685
rect 180 -2705 200 -2685
rect 220 -2705 240 -2685
rect 260 -2705 280 -2685
rect 300 -2705 320 -2685
rect 340 -2705 360 -2685
rect 380 -2705 400 -2685
rect 420 -2705 440 -2685
rect 460 -2705 480 -2685
rect 500 -2705 520 -2685
rect 540 -2705 560 -2685
rect 580 -2705 600 -2685
rect 620 -2705 640 -2685
rect 660 -2705 680 -2685
rect 700 -2705 720 -2685
rect 740 -2705 760 -2685
rect 780 -2705 800 -2685
rect 820 -2705 840 -2685
rect 860 -2705 880 -2685
rect 900 -2705 920 -2685
rect 940 -2705 960 -2685
rect 980 -2705 1000 -2685
rect 1020 -2705 1040 -2685
rect 1060 -2705 1080 -2685
rect 1100 -2705 1120 -2685
rect 1140 -2705 1160 -2685
rect 1180 -2705 1200 -2685
rect 1220 -2705 1240 -2685
rect 1260 -2705 1280 -2685
rect 1300 -2705 1320 -2685
rect 1340 -2705 1360 -2685
rect 1380 -2705 1400 -2685
rect 1420 -2705 1440 -2685
rect 1460 -2705 1480 -2685
rect 1500 -2705 1520 -2685
rect 1540 -2705 1560 -2685
rect 1580 -2705 1600 -2685
rect 1620 -2705 1640 -2685
rect 1660 -2705 1680 -2685
rect 1700 -2705 1720 -2685
rect 1740 -2705 1760 -2685
rect 1780 -2705 1800 -2685
rect 1820 -2705 1840 -2685
rect 1860 -2705 1880 -2685
rect 1900 -2705 1920 -2685
rect 1940 -2705 1960 -2685
rect 1980 -2705 2000 -2685
rect 2020 -2705 2040 -2685
rect 2060 -2705 2080 -2685
rect 2100 -2705 2120 -2685
rect 2140 -2705 2160 -2685
rect 2180 -2705 2200 -2685
rect 2220 -2705 2240 -2685
rect 2260 -2705 2280 -2685
rect 2300 -2705 2320 -2685
rect 2340 -2705 2360 -2685
rect 2380 -2705 2400 -2685
rect 2420 -2705 2440 -2685
rect 2460 -2705 2480 -2685
rect 2500 -2705 2520 -2685
rect 2540 -2705 2560 -2685
rect 2590 -2705 2605 -2685
rect 105 -2715 2605 -2705
<< ndiffc >>
rect 200 2197 220 2217
rect 240 2197 260 2217
rect 280 2197 300 2217
rect 320 2197 340 2217
rect 360 2197 380 2217
rect 400 2197 420 2217
rect 440 2197 460 2217
rect 480 2197 500 2217
rect 520 2197 540 2217
rect 560 2197 580 2217
rect 600 2197 620 2217
rect 640 2197 660 2217
rect 680 2197 700 2217
rect 720 2197 740 2217
rect 760 2197 780 2217
rect 800 2197 820 2217
rect 840 2197 860 2217
rect 880 2197 900 2217
rect 920 2197 940 2217
rect 960 2197 980 2217
rect 1000 2197 1020 2217
rect 1040 2197 1060 2217
rect 1080 2197 1100 2217
rect 1120 2197 1140 2217
rect 1160 2197 1180 2217
rect 1200 2197 1220 2217
rect 1240 2197 1260 2217
rect 1280 2197 1300 2217
rect 1320 2197 1340 2217
rect 1360 2197 1380 2217
rect 1400 2197 1420 2217
rect 1440 2197 1460 2217
rect 1480 2197 1500 2217
rect 1520 2197 1540 2217
rect 1560 2197 1580 2217
rect 1600 2197 1620 2217
rect 1640 2197 1660 2217
rect 1680 2197 1700 2217
rect 1720 2197 1740 2217
rect 1760 2197 1780 2217
rect 1800 2197 1820 2217
rect 1840 2197 1860 2217
rect 1880 2197 1900 2217
rect 1920 2197 1940 2217
rect 1960 2197 1980 2217
rect 2000 2197 2020 2217
rect 2040 2197 2060 2217
rect 2080 2197 2100 2217
rect 2120 2197 2140 2217
rect 2160 2197 2180 2217
rect 2200 2197 2220 2217
rect 2240 2197 2260 2217
rect 2280 2197 2300 2217
rect 2320 2197 2340 2217
rect 2360 2197 2380 2217
rect 2400 2197 2420 2217
rect 2440 2197 2460 2217
rect 2480 2197 2500 2217
rect 2520 2197 2540 2217
rect 2560 2197 2580 2217
rect 2600 2197 2620 2217
rect 2640 2197 2660 2217
rect 200 2115 220 2135
rect 240 2115 260 2135
rect 280 2115 300 2135
rect 320 2115 340 2135
rect 360 2115 380 2135
rect 400 2115 420 2135
rect 440 2115 460 2135
rect 480 2115 500 2135
rect 520 2115 540 2135
rect 560 2115 580 2135
rect 600 2115 620 2135
rect 640 2115 660 2135
rect 680 2115 700 2135
rect 720 2115 740 2135
rect 760 2115 780 2135
rect 800 2115 820 2135
rect 840 2115 860 2135
rect 880 2115 900 2135
rect 920 2115 940 2135
rect 960 2115 980 2135
rect 1000 2115 1020 2135
rect 1040 2115 1060 2135
rect 1080 2115 1100 2135
rect 1120 2115 1140 2135
rect 1160 2115 1180 2135
rect 1200 2115 1220 2135
rect 1240 2115 1260 2135
rect 1280 2115 1300 2135
rect 1320 2115 1340 2135
rect 1360 2115 1380 2135
rect 1400 2115 1420 2135
rect 1440 2115 1460 2135
rect 1480 2115 1500 2135
rect 1520 2115 1540 2135
rect 1560 2115 1580 2135
rect 1600 2115 1620 2135
rect 1640 2115 1660 2135
rect 1680 2115 1700 2135
rect 1720 2115 1740 2135
rect 1760 2115 1780 2135
rect 1800 2115 1820 2135
rect 1840 2115 1860 2135
rect 1880 2115 1900 2135
rect 1920 2115 1940 2135
rect 1960 2115 1980 2135
rect 2000 2115 2020 2135
rect 2040 2115 2060 2135
rect 2080 2115 2100 2135
rect 2120 2115 2140 2135
rect 2160 2115 2180 2135
rect 2200 2115 2220 2135
rect 2240 2115 2260 2135
rect 2280 2115 2300 2135
rect 2320 2115 2340 2135
rect 2360 2115 2380 2135
rect 2400 2115 2420 2135
rect 2440 2115 2460 2135
rect 2480 2115 2500 2135
rect 2520 2115 2540 2135
rect 2560 2115 2580 2135
rect 2600 2115 2620 2135
rect 2640 2115 2660 2135
rect 200 2033 220 2053
rect 240 2033 260 2053
rect 280 2033 300 2053
rect 320 2033 340 2053
rect 360 2033 380 2053
rect 400 2033 420 2053
rect 440 2033 460 2053
rect 480 2033 500 2053
rect 520 2033 540 2053
rect 560 2033 580 2053
rect 600 2033 620 2053
rect 640 2033 660 2053
rect 680 2033 700 2053
rect 720 2033 740 2053
rect 760 2033 780 2053
rect 800 2033 820 2053
rect 840 2033 860 2053
rect 880 2033 900 2053
rect 920 2033 940 2053
rect 960 2033 980 2053
rect 1000 2033 1020 2053
rect 1040 2033 1060 2053
rect 1080 2033 1100 2053
rect 1120 2033 1140 2053
rect 1160 2033 1180 2053
rect 1200 2033 1220 2053
rect 1240 2033 1260 2053
rect 1280 2033 1300 2053
rect 1320 2033 1340 2053
rect 1360 2033 1380 2053
rect 1400 2033 1420 2053
rect 1440 2033 1460 2053
rect 1480 2033 1500 2053
rect 1520 2033 1540 2053
rect 1560 2033 1580 2053
rect 1600 2033 1620 2053
rect 1640 2033 1660 2053
rect 1680 2033 1700 2053
rect 1720 2033 1740 2053
rect 1760 2033 1780 2053
rect 1800 2033 1820 2053
rect 1840 2033 1860 2053
rect 1880 2033 1900 2053
rect 1920 2033 1940 2053
rect 1960 2033 1980 2053
rect 2000 2033 2020 2053
rect 2040 2033 2060 2053
rect 2080 2033 2100 2053
rect 2120 2033 2140 2053
rect 2160 2033 2180 2053
rect 2200 2033 2220 2053
rect 2240 2033 2260 2053
rect 2280 2033 2300 2053
rect 2320 2033 2340 2053
rect 2360 2033 2380 2053
rect 2400 2033 2420 2053
rect 2440 2033 2460 2053
rect 2480 2033 2500 2053
rect 2520 2033 2540 2053
rect 2560 2033 2580 2053
rect 2600 2033 2620 2053
rect 2640 2033 2660 2053
rect 200 1951 220 1971
rect 240 1951 260 1971
rect 280 1951 300 1971
rect 320 1951 340 1971
rect 360 1951 380 1971
rect 400 1951 420 1971
rect 440 1951 460 1971
rect 480 1951 500 1971
rect 520 1951 540 1971
rect 560 1951 580 1971
rect 600 1951 620 1971
rect 640 1951 660 1971
rect 680 1951 700 1971
rect 720 1951 740 1971
rect 760 1951 780 1971
rect 800 1951 820 1971
rect 840 1951 860 1971
rect 880 1951 900 1971
rect 920 1951 940 1971
rect 960 1951 980 1971
rect 1000 1951 1020 1971
rect 1040 1951 1060 1971
rect 1080 1951 1100 1971
rect 1120 1951 1140 1971
rect 1160 1951 1180 1971
rect 1200 1951 1220 1971
rect 1240 1951 1260 1971
rect 1280 1951 1300 1971
rect 1320 1951 1340 1971
rect 1360 1951 1380 1971
rect 1400 1951 1420 1971
rect 1440 1951 1460 1971
rect 1480 1951 1500 1971
rect 1520 1951 1540 1971
rect 1560 1951 1580 1971
rect 1600 1951 1620 1971
rect 1640 1951 1660 1971
rect 1680 1951 1700 1971
rect 1720 1951 1740 1971
rect 1760 1951 1780 1971
rect 1800 1951 1820 1971
rect 1840 1951 1860 1971
rect 1880 1951 1900 1971
rect 1920 1951 1940 1971
rect 1960 1951 1980 1971
rect 2000 1951 2020 1971
rect 2040 1951 2060 1971
rect 2080 1951 2100 1971
rect 2120 1951 2140 1971
rect 2160 1951 2180 1971
rect 2200 1951 2220 1971
rect 2240 1951 2260 1971
rect 2280 1951 2300 1971
rect 2320 1951 2340 1971
rect 2360 1951 2380 1971
rect 2400 1951 2420 1971
rect 2440 1951 2460 1971
rect 2480 1951 2500 1971
rect 2520 1951 2540 1971
rect 2560 1951 2580 1971
rect 2600 1951 2620 1971
rect 2640 1951 2660 1971
rect 200 1869 220 1889
rect 240 1869 260 1889
rect 280 1869 300 1889
rect 320 1869 340 1889
rect 360 1869 380 1889
rect 400 1869 420 1889
rect 440 1869 460 1889
rect 480 1869 500 1889
rect 520 1869 540 1889
rect 560 1869 580 1889
rect 600 1869 620 1889
rect 640 1869 660 1889
rect 680 1869 700 1889
rect 720 1869 740 1889
rect 760 1869 780 1889
rect 800 1869 820 1889
rect 840 1869 860 1889
rect 880 1869 900 1889
rect 920 1869 940 1889
rect 960 1869 980 1889
rect 1000 1869 1020 1889
rect 1040 1869 1060 1889
rect 1080 1869 1100 1889
rect 1120 1869 1140 1889
rect 1160 1869 1180 1889
rect 1200 1869 1220 1889
rect 1240 1869 1260 1889
rect 1280 1869 1300 1889
rect 1320 1869 1340 1889
rect 1360 1869 1380 1889
rect 1400 1869 1420 1889
rect 1440 1869 1460 1889
rect 1480 1869 1500 1889
rect 1520 1869 1540 1889
rect 1560 1869 1580 1889
rect 1600 1869 1620 1889
rect 1640 1869 1660 1889
rect 1680 1869 1700 1889
rect 1720 1869 1740 1889
rect 1760 1869 1780 1889
rect 1800 1869 1820 1889
rect 1840 1869 1860 1889
rect 1880 1869 1900 1889
rect 1920 1869 1940 1889
rect 1960 1869 1980 1889
rect 2000 1869 2020 1889
rect 2040 1869 2060 1889
rect 2080 1869 2100 1889
rect 2120 1869 2140 1889
rect 2160 1869 2180 1889
rect 2200 1869 2220 1889
rect 2240 1869 2260 1889
rect 2280 1869 2300 1889
rect 2320 1869 2340 1889
rect 2360 1869 2380 1889
rect 2400 1869 2420 1889
rect 2440 1869 2460 1889
rect 2480 1869 2500 1889
rect 2520 1869 2540 1889
rect 2560 1869 2580 1889
rect 2600 1869 2620 1889
rect 2640 1869 2660 1889
rect 200 1787 220 1807
rect 240 1787 260 1807
rect 280 1787 300 1807
rect 320 1787 340 1807
rect 360 1787 380 1807
rect 400 1787 420 1807
rect 440 1787 460 1807
rect 480 1787 500 1807
rect 520 1787 540 1807
rect 560 1787 580 1807
rect 600 1787 620 1807
rect 640 1787 660 1807
rect 680 1787 700 1807
rect 720 1787 740 1807
rect 760 1787 780 1807
rect 800 1787 820 1807
rect 840 1787 860 1807
rect 880 1787 900 1807
rect 920 1787 940 1807
rect 960 1787 980 1807
rect 1000 1787 1020 1807
rect 1040 1787 1060 1807
rect 1080 1787 1100 1807
rect 1120 1787 1140 1807
rect 1160 1787 1180 1807
rect 1200 1787 1220 1807
rect 1240 1787 1260 1807
rect 1280 1787 1300 1807
rect 1320 1787 1340 1807
rect 1360 1787 1380 1807
rect 1400 1787 1420 1807
rect 1440 1787 1460 1807
rect 1480 1787 1500 1807
rect 1520 1787 1540 1807
rect 1560 1787 1580 1807
rect 1600 1787 1620 1807
rect 1640 1787 1660 1807
rect 1680 1787 1700 1807
rect 1720 1787 1740 1807
rect 1760 1787 1780 1807
rect 1800 1787 1820 1807
rect 1840 1787 1860 1807
rect 1880 1787 1900 1807
rect 1920 1787 1940 1807
rect 1960 1787 1980 1807
rect 2000 1787 2020 1807
rect 2040 1787 2060 1807
rect 2080 1787 2100 1807
rect 2120 1787 2140 1807
rect 2160 1787 2180 1807
rect 2200 1787 2220 1807
rect 2240 1787 2260 1807
rect 2280 1787 2300 1807
rect 2320 1787 2340 1807
rect 2360 1787 2380 1807
rect 2400 1787 2420 1807
rect 2440 1787 2460 1807
rect 2480 1787 2500 1807
rect 2520 1787 2540 1807
rect 2560 1787 2580 1807
rect 2600 1787 2620 1807
rect 2640 1787 2660 1807
rect 200 1705 220 1725
rect 240 1705 260 1725
rect 280 1705 300 1725
rect 320 1705 340 1725
rect 360 1705 380 1725
rect 400 1705 420 1725
rect 440 1705 460 1725
rect 480 1705 500 1725
rect 520 1705 540 1725
rect 560 1705 580 1725
rect 600 1705 620 1725
rect 640 1705 660 1725
rect 680 1705 700 1725
rect 720 1705 740 1725
rect 760 1705 780 1725
rect 800 1705 820 1725
rect 840 1705 860 1725
rect 880 1705 900 1725
rect 920 1705 940 1725
rect 960 1705 980 1725
rect 1000 1705 1020 1725
rect 1040 1705 1060 1725
rect 1080 1705 1100 1725
rect 1120 1705 1140 1725
rect 1160 1705 1180 1725
rect 1200 1705 1220 1725
rect 1240 1705 1260 1725
rect 1280 1705 1300 1725
rect 1320 1705 1340 1725
rect 1360 1705 1380 1725
rect 1400 1705 1420 1725
rect 1440 1705 1460 1725
rect 1480 1705 1500 1725
rect 1520 1705 1540 1725
rect 1560 1705 1580 1725
rect 1600 1705 1620 1725
rect 1640 1705 1660 1725
rect 1680 1705 1700 1725
rect 1720 1705 1740 1725
rect 1760 1705 1780 1725
rect 1800 1705 1820 1725
rect 1840 1705 1860 1725
rect 1880 1705 1900 1725
rect 1920 1705 1940 1725
rect 1960 1705 1980 1725
rect 2000 1705 2020 1725
rect 2040 1705 2060 1725
rect 2080 1705 2100 1725
rect 2120 1705 2140 1725
rect 2160 1705 2180 1725
rect 2200 1705 2220 1725
rect 2240 1705 2260 1725
rect 2280 1705 2300 1725
rect 2320 1705 2340 1725
rect 2360 1705 2380 1725
rect 2400 1705 2420 1725
rect 2440 1705 2460 1725
rect 2480 1705 2500 1725
rect 2520 1705 2540 1725
rect 2560 1705 2580 1725
rect 2600 1705 2620 1725
rect 2640 1705 2660 1725
rect 200 1623 220 1643
rect 240 1623 260 1643
rect 280 1623 300 1643
rect 320 1623 340 1643
rect 360 1623 380 1643
rect 400 1623 420 1643
rect 440 1623 460 1643
rect 480 1623 500 1643
rect 520 1623 540 1643
rect 560 1623 580 1643
rect 600 1623 620 1643
rect 640 1623 660 1643
rect 680 1623 700 1643
rect 720 1623 740 1643
rect 760 1623 780 1643
rect 800 1623 820 1643
rect 840 1623 860 1643
rect 880 1623 900 1643
rect 920 1623 940 1643
rect 960 1623 980 1643
rect 1000 1623 1020 1643
rect 1040 1623 1060 1643
rect 1080 1623 1100 1643
rect 1120 1623 1140 1643
rect 1160 1623 1180 1643
rect 1200 1623 1220 1643
rect 1240 1623 1260 1643
rect 1280 1623 1300 1643
rect 1320 1623 1340 1643
rect 1360 1623 1380 1643
rect 1400 1623 1420 1643
rect 1440 1623 1460 1643
rect 1480 1623 1500 1643
rect 1520 1623 1540 1643
rect 1560 1623 1580 1643
rect 1600 1623 1620 1643
rect 1640 1623 1660 1643
rect 1680 1623 1700 1643
rect 1720 1623 1740 1643
rect 1760 1623 1780 1643
rect 1800 1623 1820 1643
rect 1840 1623 1860 1643
rect 1880 1623 1900 1643
rect 1920 1623 1940 1643
rect 1960 1623 1980 1643
rect 2000 1623 2020 1643
rect 2040 1623 2060 1643
rect 2080 1623 2100 1643
rect 2120 1623 2140 1643
rect 2160 1623 2180 1643
rect 2200 1623 2220 1643
rect 2240 1623 2260 1643
rect 2280 1623 2300 1643
rect 2320 1623 2340 1643
rect 2360 1623 2380 1643
rect 2400 1623 2420 1643
rect 2440 1623 2460 1643
rect 2480 1623 2500 1643
rect 2520 1623 2540 1643
rect 2560 1623 2580 1643
rect 2600 1623 2620 1643
rect 2640 1623 2660 1643
rect 200 1541 220 1561
rect 240 1541 260 1561
rect 280 1541 300 1561
rect 320 1541 340 1561
rect 360 1541 380 1561
rect 400 1541 420 1561
rect 440 1541 460 1561
rect 480 1541 500 1561
rect 520 1541 540 1561
rect 560 1541 580 1561
rect 600 1541 620 1561
rect 640 1541 660 1561
rect 680 1541 700 1561
rect 720 1541 740 1561
rect 760 1541 780 1561
rect 800 1541 820 1561
rect 840 1541 860 1561
rect 880 1541 900 1561
rect 920 1541 940 1561
rect 960 1541 980 1561
rect 1000 1541 1020 1561
rect 1040 1541 1060 1561
rect 1080 1541 1100 1561
rect 1120 1541 1140 1561
rect 1160 1541 1180 1561
rect 1200 1541 1220 1561
rect 1240 1541 1260 1561
rect 1280 1541 1300 1561
rect 1320 1541 1340 1561
rect 1360 1541 1380 1561
rect 1400 1541 1420 1561
rect 1440 1541 1460 1561
rect 1480 1541 1500 1561
rect 1520 1541 1540 1561
rect 1560 1541 1580 1561
rect 1600 1541 1620 1561
rect 1640 1541 1660 1561
rect 1680 1541 1700 1561
rect 1720 1541 1740 1561
rect 1760 1541 1780 1561
rect 1800 1541 1820 1561
rect 1840 1541 1860 1561
rect 1880 1541 1900 1561
rect 1920 1541 1940 1561
rect 1960 1541 1980 1561
rect 2000 1541 2020 1561
rect 2040 1541 2060 1561
rect 2080 1541 2100 1561
rect 2120 1541 2140 1561
rect 2160 1541 2180 1561
rect 2200 1541 2220 1561
rect 2240 1541 2260 1561
rect 2280 1541 2300 1561
rect 2320 1541 2340 1561
rect 2360 1541 2380 1561
rect 2400 1541 2420 1561
rect 2440 1541 2460 1561
rect 2480 1541 2500 1561
rect 2520 1541 2540 1561
rect 2560 1541 2580 1561
rect 2600 1541 2620 1561
rect 2640 1541 2660 1561
rect 200 1459 220 1479
rect 240 1459 260 1479
rect 280 1459 300 1479
rect 320 1459 340 1479
rect 360 1459 380 1479
rect 400 1459 420 1479
rect 440 1459 460 1479
rect 480 1459 500 1479
rect 520 1459 540 1479
rect 560 1459 580 1479
rect 600 1459 620 1479
rect 640 1459 660 1479
rect 680 1459 700 1479
rect 720 1459 740 1479
rect 760 1459 780 1479
rect 800 1459 820 1479
rect 840 1459 860 1479
rect 880 1459 900 1479
rect 920 1459 940 1479
rect 960 1459 980 1479
rect 1000 1459 1020 1479
rect 1040 1459 1060 1479
rect 1080 1459 1100 1479
rect 1120 1459 1140 1479
rect 1160 1459 1180 1479
rect 1200 1459 1220 1479
rect 1240 1459 1260 1479
rect 1280 1459 1300 1479
rect 1320 1459 1340 1479
rect 1360 1459 1380 1479
rect 1400 1459 1420 1479
rect 1440 1459 1460 1479
rect 1480 1459 1500 1479
rect 1520 1459 1540 1479
rect 1560 1459 1580 1479
rect 1600 1459 1620 1479
rect 1640 1459 1660 1479
rect 1680 1459 1700 1479
rect 1720 1459 1740 1479
rect 1760 1459 1780 1479
rect 1800 1459 1820 1479
rect 1840 1459 1860 1479
rect 1880 1459 1900 1479
rect 1920 1459 1940 1479
rect 1960 1459 1980 1479
rect 2000 1459 2020 1479
rect 2040 1459 2060 1479
rect 2080 1459 2100 1479
rect 2120 1459 2140 1479
rect 2160 1459 2180 1479
rect 2200 1459 2220 1479
rect 2240 1459 2260 1479
rect 2280 1459 2300 1479
rect 2320 1459 2340 1479
rect 2360 1459 2380 1479
rect 2400 1459 2420 1479
rect 2440 1459 2460 1479
rect 2480 1459 2500 1479
rect 2520 1459 2540 1479
rect 2560 1459 2580 1479
rect 2600 1459 2620 1479
rect 2640 1459 2660 1479
rect 200 1377 220 1397
rect 240 1377 260 1397
rect 280 1377 300 1397
rect 320 1377 340 1397
rect 360 1377 380 1397
rect 400 1377 420 1397
rect 440 1377 460 1397
rect 480 1377 500 1397
rect 520 1377 540 1397
rect 560 1377 580 1397
rect 600 1377 620 1397
rect 640 1377 660 1397
rect 680 1377 700 1397
rect 720 1377 740 1397
rect 760 1377 780 1397
rect 800 1377 820 1397
rect 840 1377 860 1397
rect 880 1377 900 1397
rect 920 1377 940 1397
rect 960 1377 980 1397
rect 1000 1377 1020 1397
rect 1040 1377 1060 1397
rect 1080 1377 1100 1397
rect 1120 1377 1140 1397
rect 1160 1377 1180 1397
rect 1200 1377 1220 1397
rect 1240 1377 1260 1397
rect 1280 1377 1300 1397
rect 1320 1377 1340 1397
rect 1360 1377 1380 1397
rect 1400 1377 1420 1397
rect 1440 1377 1460 1397
rect 1480 1377 1500 1397
rect 1520 1377 1540 1397
rect 1560 1377 1580 1397
rect 1600 1377 1620 1397
rect 1640 1377 1660 1397
rect 1680 1377 1700 1397
rect 1720 1377 1740 1397
rect 1760 1377 1780 1397
rect 1800 1377 1820 1397
rect 1840 1377 1860 1397
rect 1880 1377 1900 1397
rect 1920 1377 1940 1397
rect 1960 1377 1980 1397
rect 2000 1377 2020 1397
rect 2040 1377 2060 1397
rect 2080 1377 2100 1397
rect 2120 1377 2140 1397
rect 2160 1377 2180 1397
rect 2200 1377 2220 1397
rect 2240 1377 2260 1397
rect 2280 1377 2300 1397
rect 2320 1377 2340 1397
rect 2360 1377 2380 1397
rect 2400 1377 2420 1397
rect 2440 1377 2460 1397
rect 2480 1377 2500 1397
rect 2520 1377 2540 1397
rect 2560 1377 2580 1397
rect 2600 1377 2620 1397
rect 2640 1377 2660 1397
rect 200 1295 220 1315
rect 240 1295 260 1315
rect 280 1295 300 1315
rect 320 1295 340 1315
rect 360 1295 380 1315
rect 400 1295 420 1315
rect 440 1295 460 1315
rect 480 1295 500 1315
rect 520 1295 540 1315
rect 560 1295 580 1315
rect 600 1295 620 1315
rect 640 1295 660 1315
rect 680 1295 700 1315
rect 720 1295 740 1315
rect 760 1295 780 1315
rect 800 1295 820 1315
rect 840 1295 860 1315
rect 880 1295 900 1315
rect 920 1295 940 1315
rect 960 1295 980 1315
rect 1000 1295 1020 1315
rect 1040 1295 1060 1315
rect 1080 1295 1100 1315
rect 1120 1295 1140 1315
rect 1160 1295 1180 1315
rect 1200 1295 1220 1315
rect 1240 1295 1260 1315
rect 1280 1295 1300 1315
rect 1320 1295 1340 1315
rect 1360 1295 1380 1315
rect 1400 1295 1420 1315
rect 1440 1295 1460 1315
rect 1480 1295 1500 1315
rect 1520 1295 1540 1315
rect 1560 1295 1580 1315
rect 1600 1295 1620 1315
rect 1640 1295 1660 1315
rect 1680 1295 1700 1315
rect 1720 1295 1740 1315
rect 1760 1295 1780 1315
rect 1800 1295 1820 1315
rect 1840 1295 1860 1315
rect 1880 1295 1900 1315
rect 1920 1295 1940 1315
rect 1960 1295 1980 1315
rect 2000 1295 2020 1315
rect 2040 1295 2060 1315
rect 2080 1295 2100 1315
rect 2120 1295 2140 1315
rect 2160 1295 2180 1315
rect 2200 1295 2220 1315
rect 2240 1295 2260 1315
rect 2280 1295 2300 1315
rect 2320 1295 2340 1315
rect 2360 1295 2380 1315
rect 2400 1295 2420 1315
rect 2440 1295 2460 1315
rect 2480 1295 2500 1315
rect 2520 1295 2540 1315
rect 2560 1295 2580 1315
rect 2600 1295 2620 1315
rect 2640 1295 2660 1315
rect 200 1213 220 1233
rect 240 1213 260 1233
rect 280 1213 300 1233
rect 320 1213 340 1233
rect 360 1213 380 1233
rect 400 1213 420 1233
rect 440 1213 460 1233
rect 480 1213 500 1233
rect 520 1213 540 1233
rect 560 1213 580 1233
rect 600 1213 620 1233
rect 640 1213 660 1233
rect 680 1213 700 1233
rect 720 1213 740 1233
rect 760 1213 780 1233
rect 800 1213 820 1233
rect 840 1213 860 1233
rect 880 1213 900 1233
rect 920 1213 940 1233
rect 960 1213 980 1233
rect 1000 1213 1020 1233
rect 1040 1213 1060 1233
rect 1080 1213 1100 1233
rect 1120 1213 1140 1233
rect 1160 1213 1180 1233
rect 1200 1213 1220 1233
rect 1240 1213 1260 1233
rect 1280 1213 1300 1233
rect 1320 1213 1340 1233
rect 1360 1213 1380 1233
rect 1400 1213 1420 1233
rect 1440 1213 1460 1233
rect 1480 1213 1500 1233
rect 1520 1213 1540 1233
rect 1560 1213 1580 1233
rect 1600 1213 1620 1233
rect 1640 1213 1660 1233
rect 1680 1213 1700 1233
rect 1720 1213 1740 1233
rect 1760 1213 1780 1233
rect 1800 1213 1820 1233
rect 1840 1213 1860 1233
rect 1880 1213 1900 1233
rect 1920 1213 1940 1233
rect 1960 1213 1980 1233
rect 2000 1213 2020 1233
rect 2040 1213 2060 1233
rect 2080 1213 2100 1233
rect 2120 1213 2140 1233
rect 2160 1213 2180 1233
rect 2200 1213 2220 1233
rect 2240 1213 2260 1233
rect 2280 1213 2300 1233
rect 2320 1213 2340 1233
rect 2360 1213 2380 1233
rect 2400 1213 2420 1233
rect 2440 1213 2460 1233
rect 2480 1213 2500 1233
rect 2520 1213 2540 1233
rect 2560 1213 2580 1233
rect 2600 1213 2620 1233
rect 2640 1213 2660 1233
rect 200 1131 220 1151
rect 240 1131 260 1151
rect 280 1131 300 1151
rect 320 1131 340 1151
rect 360 1131 380 1151
rect 400 1131 420 1151
rect 440 1131 460 1151
rect 480 1131 500 1151
rect 520 1131 540 1151
rect 560 1131 580 1151
rect 600 1131 620 1151
rect 640 1131 660 1151
rect 680 1131 700 1151
rect 720 1131 740 1151
rect 760 1131 780 1151
rect 800 1131 820 1151
rect 840 1131 860 1151
rect 880 1131 900 1151
rect 920 1131 940 1151
rect 960 1131 980 1151
rect 1000 1131 1020 1151
rect 1040 1131 1060 1151
rect 1080 1131 1100 1151
rect 1120 1131 1140 1151
rect 1160 1131 1180 1151
rect 1200 1131 1220 1151
rect 1240 1131 1260 1151
rect 1280 1131 1300 1151
rect 1320 1131 1340 1151
rect 1360 1131 1380 1151
rect 1400 1131 1420 1151
rect 1440 1131 1460 1151
rect 1480 1131 1500 1151
rect 1520 1131 1540 1151
rect 1560 1131 1580 1151
rect 1600 1131 1620 1151
rect 1640 1131 1660 1151
rect 1680 1131 1700 1151
rect 1720 1131 1740 1151
rect 1760 1131 1780 1151
rect 1800 1131 1820 1151
rect 1840 1131 1860 1151
rect 1880 1131 1900 1151
rect 1920 1131 1940 1151
rect 1960 1131 1980 1151
rect 2000 1131 2020 1151
rect 2040 1131 2060 1151
rect 2080 1131 2100 1151
rect 2120 1131 2140 1151
rect 2160 1131 2180 1151
rect 2200 1131 2220 1151
rect 2240 1131 2260 1151
rect 2280 1131 2300 1151
rect 2320 1131 2340 1151
rect 2360 1131 2380 1151
rect 2400 1131 2420 1151
rect 2440 1131 2460 1151
rect 2480 1131 2500 1151
rect 2520 1131 2540 1151
rect 2560 1131 2580 1151
rect 2600 1131 2620 1151
rect 2640 1131 2660 1151
rect 200 1049 220 1069
rect 240 1049 260 1069
rect 280 1049 300 1069
rect 320 1049 340 1069
rect 360 1049 380 1069
rect 400 1049 420 1069
rect 440 1049 460 1069
rect 480 1049 500 1069
rect 520 1049 540 1069
rect 560 1049 580 1069
rect 600 1049 620 1069
rect 640 1049 660 1069
rect 680 1049 700 1069
rect 720 1049 740 1069
rect 760 1049 780 1069
rect 800 1049 820 1069
rect 840 1049 860 1069
rect 880 1049 900 1069
rect 920 1049 940 1069
rect 960 1049 980 1069
rect 1000 1049 1020 1069
rect 1040 1049 1060 1069
rect 1080 1049 1100 1069
rect 1120 1049 1140 1069
rect 1160 1049 1180 1069
rect 1200 1049 1220 1069
rect 1240 1049 1260 1069
rect 1280 1049 1300 1069
rect 1320 1049 1340 1069
rect 1360 1049 1380 1069
rect 1400 1049 1420 1069
rect 1440 1049 1460 1069
rect 1480 1049 1500 1069
rect 1520 1049 1540 1069
rect 1560 1049 1580 1069
rect 1600 1049 1620 1069
rect 1640 1049 1660 1069
rect 1680 1049 1700 1069
rect 1720 1049 1740 1069
rect 1760 1049 1780 1069
rect 1800 1049 1820 1069
rect 1840 1049 1860 1069
rect 1880 1049 1900 1069
rect 1920 1049 1940 1069
rect 1960 1049 1980 1069
rect 2000 1049 2020 1069
rect 2040 1049 2060 1069
rect 2080 1049 2100 1069
rect 2120 1049 2140 1069
rect 2160 1049 2180 1069
rect 2200 1049 2220 1069
rect 2240 1049 2260 1069
rect 2280 1049 2300 1069
rect 2320 1049 2340 1069
rect 2360 1049 2380 1069
rect 2400 1049 2420 1069
rect 2440 1049 2460 1069
rect 2480 1049 2500 1069
rect 2520 1049 2540 1069
rect 2560 1049 2580 1069
rect 2600 1049 2620 1069
rect 2640 1049 2660 1069
rect 200 967 220 987
rect 240 967 260 987
rect 280 967 300 987
rect 320 967 340 987
rect 360 967 380 987
rect 400 967 420 987
rect 440 967 460 987
rect 480 967 500 987
rect 520 967 540 987
rect 560 967 580 987
rect 600 967 620 987
rect 640 967 660 987
rect 680 967 700 987
rect 720 967 740 987
rect 760 967 780 987
rect 800 967 820 987
rect 840 967 860 987
rect 880 967 900 987
rect 920 967 940 987
rect 960 967 980 987
rect 1000 967 1020 987
rect 1040 967 1060 987
rect 1080 967 1100 987
rect 1120 967 1140 987
rect 1160 967 1180 987
rect 1200 967 1220 987
rect 1240 967 1260 987
rect 1280 967 1300 987
rect 1320 967 1340 987
rect 1360 967 1380 987
rect 1400 967 1420 987
rect 1440 967 1460 987
rect 1480 967 1500 987
rect 1520 967 1540 987
rect 1560 967 1580 987
rect 1600 967 1620 987
rect 1640 967 1660 987
rect 1680 967 1700 987
rect 1720 967 1740 987
rect 1760 967 1780 987
rect 1800 967 1820 987
rect 1840 967 1860 987
rect 1880 967 1900 987
rect 1920 967 1940 987
rect 1960 967 1980 987
rect 2000 967 2020 987
rect 2040 967 2060 987
rect 2080 967 2100 987
rect 2120 967 2140 987
rect 2160 967 2180 987
rect 2200 967 2220 987
rect 2240 967 2260 987
rect 2280 967 2300 987
rect 2320 967 2340 987
rect 2360 967 2380 987
rect 2400 967 2420 987
rect 2440 967 2460 987
rect 2480 967 2500 987
rect 2520 967 2540 987
rect 2560 967 2580 987
rect 2600 967 2620 987
rect 2640 967 2660 987
rect 200 885 220 905
rect 240 885 260 905
rect 280 885 300 905
rect 320 885 340 905
rect 360 885 380 905
rect 400 885 420 905
rect 440 885 460 905
rect 480 885 500 905
rect 520 885 540 905
rect 560 885 580 905
rect 600 885 620 905
rect 640 885 660 905
rect 680 885 700 905
rect 720 885 740 905
rect 760 885 780 905
rect 800 885 820 905
rect 840 885 860 905
rect 880 885 900 905
rect 920 885 940 905
rect 960 885 980 905
rect 1000 885 1020 905
rect 1040 885 1060 905
rect 1080 885 1100 905
rect 1120 885 1140 905
rect 1160 885 1180 905
rect 1200 885 1220 905
rect 1240 885 1260 905
rect 1280 885 1300 905
rect 1320 885 1340 905
rect 1360 885 1380 905
rect 1400 885 1420 905
rect 1440 885 1460 905
rect 1480 885 1500 905
rect 1520 885 1540 905
rect 1560 885 1580 905
rect 1600 885 1620 905
rect 1640 885 1660 905
rect 1680 885 1700 905
rect 1720 885 1740 905
rect 1760 885 1780 905
rect 1800 885 1820 905
rect 1840 885 1860 905
rect 1880 885 1900 905
rect 1920 885 1940 905
rect 1960 885 1980 905
rect 2000 885 2020 905
rect 2040 885 2060 905
rect 2080 885 2100 905
rect 2120 885 2140 905
rect 2160 885 2180 905
rect 2200 885 2220 905
rect 2240 885 2260 905
rect 2280 885 2300 905
rect 2320 885 2340 905
rect 2360 885 2380 905
rect 2400 885 2420 905
rect 2440 885 2460 905
rect 2480 885 2500 905
rect 2520 885 2540 905
rect 2560 885 2580 905
rect 2600 885 2620 905
rect 2640 885 2660 905
rect 200 803 220 823
rect 240 803 260 823
rect 280 803 300 823
rect 320 803 340 823
rect 360 803 380 823
rect 400 803 420 823
rect 440 803 460 823
rect 480 803 500 823
rect 520 803 540 823
rect 560 803 580 823
rect 600 803 620 823
rect 640 803 660 823
rect 680 803 700 823
rect 720 803 740 823
rect 760 803 780 823
rect 800 803 820 823
rect 840 803 860 823
rect 880 803 900 823
rect 920 803 940 823
rect 960 803 980 823
rect 1000 803 1020 823
rect 1040 803 1060 823
rect 1080 803 1100 823
rect 1120 803 1140 823
rect 1160 803 1180 823
rect 1200 803 1220 823
rect 1240 803 1260 823
rect 1280 803 1300 823
rect 1320 803 1340 823
rect 1360 803 1380 823
rect 1400 803 1420 823
rect 1440 803 1460 823
rect 1480 803 1500 823
rect 1520 803 1540 823
rect 1560 803 1580 823
rect 1600 803 1620 823
rect 1640 803 1660 823
rect 1680 803 1700 823
rect 1720 803 1740 823
rect 1760 803 1780 823
rect 1800 803 1820 823
rect 1840 803 1860 823
rect 1880 803 1900 823
rect 1920 803 1940 823
rect 1960 803 1980 823
rect 2000 803 2020 823
rect 2040 803 2060 823
rect 2080 803 2100 823
rect 2120 803 2140 823
rect 2160 803 2180 823
rect 2200 803 2220 823
rect 2240 803 2260 823
rect 2280 803 2300 823
rect 2320 803 2340 823
rect 2360 803 2380 823
rect 2400 803 2420 823
rect 2440 803 2460 823
rect 2480 803 2500 823
rect 2520 803 2540 823
rect 2560 803 2580 823
rect 2600 803 2620 823
rect 2640 803 2660 823
rect 200 721 220 741
rect 240 721 260 741
rect 280 721 300 741
rect 320 721 340 741
rect 360 721 380 741
rect 400 721 420 741
rect 440 721 460 741
rect 480 721 500 741
rect 520 721 540 741
rect 560 721 580 741
rect 600 721 620 741
rect 640 721 660 741
rect 680 721 700 741
rect 720 721 740 741
rect 760 721 780 741
rect 800 721 820 741
rect 840 721 860 741
rect 880 721 900 741
rect 920 721 940 741
rect 960 721 980 741
rect 1000 721 1020 741
rect 1040 721 1060 741
rect 1080 721 1100 741
rect 1120 721 1140 741
rect 1160 721 1180 741
rect 1200 721 1220 741
rect 1240 721 1260 741
rect 1280 721 1300 741
rect 1320 721 1340 741
rect 1360 721 1380 741
rect 1400 721 1420 741
rect 1440 721 1460 741
rect 1480 721 1500 741
rect 1520 721 1540 741
rect 1560 721 1580 741
rect 1600 721 1620 741
rect 1640 721 1660 741
rect 1680 721 1700 741
rect 1720 721 1740 741
rect 1760 721 1780 741
rect 1800 721 1820 741
rect 1840 721 1860 741
rect 1880 721 1900 741
rect 1920 721 1940 741
rect 1960 721 1980 741
rect 2000 721 2020 741
rect 2040 721 2060 741
rect 2080 721 2100 741
rect 2120 721 2140 741
rect 2160 721 2180 741
rect 2200 721 2220 741
rect 2240 721 2260 741
rect 2280 721 2300 741
rect 2320 721 2340 741
rect 2360 721 2380 741
rect 2400 721 2420 741
rect 2440 721 2460 741
rect 2480 721 2500 741
rect 2520 721 2540 741
rect 2560 721 2580 741
rect 2600 721 2620 741
rect 2640 721 2660 741
rect 200 639 220 659
rect 240 639 260 659
rect 280 639 300 659
rect 320 639 340 659
rect 360 639 380 659
rect 400 639 420 659
rect 440 639 460 659
rect 480 639 500 659
rect 520 639 540 659
rect 560 639 580 659
rect 600 639 620 659
rect 640 639 660 659
rect 680 639 700 659
rect 720 639 740 659
rect 760 639 780 659
rect 800 639 820 659
rect 840 639 860 659
rect 880 639 900 659
rect 920 639 940 659
rect 960 639 980 659
rect 1000 639 1020 659
rect 1040 639 1060 659
rect 1080 639 1100 659
rect 1120 639 1140 659
rect 1160 639 1180 659
rect 1200 639 1220 659
rect 1240 639 1260 659
rect 1280 639 1300 659
rect 1320 639 1340 659
rect 1360 639 1380 659
rect 1400 639 1420 659
rect 1440 639 1460 659
rect 1480 639 1500 659
rect 1520 639 1540 659
rect 1560 639 1580 659
rect 1600 639 1620 659
rect 1640 639 1660 659
rect 1680 639 1700 659
rect 1720 639 1740 659
rect 1760 639 1780 659
rect 1800 639 1820 659
rect 1840 639 1860 659
rect 1880 639 1900 659
rect 1920 639 1940 659
rect 1960 639 1980 659
rect 2000 639 2020 659
rect 2040 639 2060 659
rect 2080 639 2100 659
rect 2120 639 2140 659
rect 2160 639 2180 659
rect 2200 639 2220 659
rect 2240 639 2260 659
rect 2280 639 2300 659
rect 2320 639 2340 659
rect 2360 639 2380 659
rect 2400 639 2420 659
rect 2440 639 2460 659
rect 2480 639 2500 659
rect 2520 639 2540 659
rect 2560 639 2580 659
rect 2600 639 2620 659
rect 2640 639 2660 659
rect 200 557 220 577
rect 240 557 260 577
rect 280 557 300 577
rect 320 557 340 577
rect 360 557 380 577
rect 400 557 420 577
rect 440 557 460 577
rect 480 557 500 577
rect 520 557 540 577
rect 560 557 580 577
rect 600 557 620 577
rect 640 557 660 577
rect 680 557 700 577
rect 720 557 740 577
rect 760 557 780 577
rect 800 557 820 577
rect 840 557 860 577
rect 880 557 900 577
rect 920 557 940 577
rect 960 557 980 577
rect 1000 557 1020 577
rect 1040 557 1060 577
rect 1080 557 1100 577
rect 1120 557 1140 577
rect 1160 557 1180 577
rect 1200 557 1220 577
rect 1240 557 1260 577
rect 1280 557 1300 577
rect 1320 557 1340 577
rect 1360 557 1380 577
rect 1400 557 1420 577
rect 1440 557 1460 577
rect 1480 557 1500 577
rect 1520 557 1540 577
rect 1560 557 1580 577
rect 1600 557 1620 577
rect 1640 557 1660 577
rect 1680 557 1700 577
rect 1720 557 1740 577
rect 1760 557 1780 577
rect 1800 557 1820 577
rect 1840 557 1860 577
rect 1880 557 1900 577
rect 1920 557 1940 577
rect 1960 557 1980 577
rect 2000 557 2020 577
rect 2040 557 2060 577
rect 2080 557 2100 577
rect 2120 557 2140 577
rect 2160 557 2180 577
rect 2200 557 2220 577
rect 2240 557 2260 577
rect 2280 557 2300 577
rect 2320 557 2340 577
rect 2360 557 2380 577
rect 2400 557 2420 577
rect 2440 557 2460 577
rect 2480 557 2500 577
rect 2520 557 2540 577
rect 2560 557 2580 577
rect 2600 557 2620 577
rect 2640 557 2660 577
rect 200 475 220 495
rect 240 475 260 495
rect 280 475 300 495
rect 320 475 340 495
rect 360 475 380 495
rect 400 475 420 495
rect 440 475 460 495
rect 480 475 500 495
rect 520 475 540 495
rect 560 475 580 495
rect 600 475 620 495
rect 640 475 660 495
rect 680 475 700 495
rect 720 475 740 495
rect 760 475 780 495
rect 800 475 820 495
rect 840 475 860 495
rect 880 475 900 495
rect 920 475 940 495
rect 960 475 980 495
rect 1000 475 1020 495
rect 1040 475 1060 495
rect 1080 475 1100 495
rect 1120 475 1140 495
rect 1160 475 1180 495
rect 1200 475 1220 495
rect 1240 475 1260 495
rect 1280 475 1300 495
rect 1320 475 1340 495
rect 1360 475 1380 495
rect 1400 475 1420 495
rect 1440 475 1460 495
rect 1480 475 1500 495
rect 1520 475 1540 495
rect 1560 475 1580 495
rect 1600 475 1620 495
rect 1640 475 1660 495
rect 1680 475 1700 495
rect 1720 475 1740 495
rect 1760 475 1780 495
rect 1800 475 1820 495
rect 1840 475 1860 495
rect 1880 475 1900 495
rect 1920 475 1940 495
rect 1960 475 1980 495
rect 2000 475 2020 495
rect 2040 475 2060 495
rect 2080 475 2100 495
rect 2120 475 2140 495
rect 2160 475 2180 495
rect 2200 475 2220 495
rect 2240 475 2260 495
rect 2280 475 2300 495
rect 2320 475 2340 495
rect 2360 475 2380 495
rect 2400 475 2420 495
rect 2440 475 2460 495
rect 2480 475 2500 495
rect 2520 475 2540 495
rect 2560 475 2580 495
rect 2600 475 2620 495
rect 2640 475 2660 495
rect 200 393 220 413
rect 240 393 260 413
rect 280 393 300 413
rect 320 393 340 413
rect 360 393 380 413
rect 400 393 420 413
rect 440 393 460 413
rect 480 393 500 413
rect 520 393 540 413
rect 560 393 580 413
rect 600 393 620 413
rect 640 393 660 413
rect 680 393 700 413
rect 720 393 740 413
rect 760 393 780 413
rect 800 393 820 413
rect 840 393 860 413
rect 880 393 900 413
rect 920 393 940 413
rect 960 393 980 413
rect 1000 393 1020 413
rect 1040 393 1060 413
rect 1080 393 1100 413
rect 1120 393 1140 413
rect 1160 393 1180 413
rect 1200 393 1220 413
rect 1240 393 1260 413
rect 1280 393 1300 413
rect 1320 393 1340 413
rect 1360 393 1380 413
rect 1400 393 1420 413
rect 1440 393 1460 413
rect 1480 393 1500 413
rect 1520 393 1540 413
rect 1560 393 1580 413
rect 1600 393 1620 413
rect 1640 393 1660 413
rect 1680 393 1700 413
rect 1720 393 1740 413
rect 1760 393 1780 413
rect 1800 393 1820 413
rect 1840 393 1860 413
rect 1880 393 1900 413
rect 1920 393 1940 413
rect 1960 393 1980 413
rect 2000 393 2020 413
rect 2040 393 2060 413
rect 2080 393 2100 413
rect 2120 393 2140 413
rect 2160 393 2180 413
rect 2200 393 2220 413
rect 2240 393 2260 413
rect 2280 393 2300 413
rect 2320 393 2340 413
rect 2360 393 2380 413
rect 2400 393 2420 413
rect 2440 393 2460 413
rect 2480 393 2500 413
rect 2520 393 2540 413
rect 2560 393 2580 413
rect 2600 393 2620 413
rect 2640 393 2660 413
rect 200 311 220 331
rect 240 311 260 331
rect 280 311 300 331
rect 320 311 340 331
rect 360 311 380 331
rect 400 311 420 331
rect 440 311 460 331
rect 480 311 500 331
rect 520 311 540 331
rect 560 311 580 331
rect 600 311 620 331
rect 640 311 660 331
rect 680 311 700 331
rect 720 311 740 331
rect 760 311 780 331
rect 800 311 820 331
rect 840 311 860 331
rect 880 311 900 331
rect 920 311 940 331
rect 960 311 980 331
rect 1000 311 1020 331
rect 1040 311 1060 331
rect 1080 311 1100 331
rect 1120 311 1140 331
rect 1160 311 1180 331
rect 1200 311 1220 331
rect 1240 311 1260 331
rect 1280 311 1300 331
rect 1320 311 1340 331
rect 1360 311 1380 331
rect 1400 311 1420 331
rect 1440 311 1460 331
rect 1480 311 1500 331
rect 1520 311 1540 331
rect 1560 311 1580 331
rect 1600 311 1620 331
rect 1640 311 1660 331
rect 1680 311 1700 331
rect 1720 311 1740 331
rect 1760 311 1780 331
rect 1800 311 1820 331
rect 1840 311 1860 331
rect 1880 311 1900 331
rect 1920 311 1940 331
rect 1960 311 1980 331
rect 2000 311 2020 331
rect 2040 311 2060 331
rect 2080 311 2100 331
rect 2120 311 2140 331
rect 2160 311 2180 331
rect 2200 311 2220 331
rect 2240 311 2260 331
rect 2280 311 2300 331
rect 2320 311 2340 331
rect 2360 311 2380 331
rect 2400 311 2420 331
rect 2440 311 2460 331
rect 2480 311 2500 331
rect 2520 311 2540 331
rect 2560 311 2580 331
rect 2600 311 2620 331
rect 2640 311 2660 331
rect 200 229 220 249
rect 240 229 260 249
rect 280 229 300 249
rect 320 229 340 249
rect 360 229 380 249
rect 400 229 420 249
rect 440 229 460 249
rect 480 229 500 249
rect 520 229 540 249
rect 560 229 580 249
rect 600 229 620 249
rect 640 229 660 249
rect 680 229 700 249
rect 720 229 740 249
rect 760 229 780 249
rect 800 229 820 249
rect 840 229 860 249
rect 880 229 900 249
rect 920 229 940 249
rect 960 229 980 249
rect 1000 229 1020 249
rect 1040 229 1060 249
rect 1080 229 1100 249
rect 1120 229 1140 249
rect 1160 229 1180 249
rect 1200 229 1220 249
rect 1240 229 1260 249
rect 1280 229 1300 249
rect 1320 229 1340 249
rect 1360 229 1380 249
rect 1400 229 1420 249
rect 1440 229 1460 249
rect 1480 229 1500 249
rect 1520 229 1540 249
rect 1560 229 1580 249
rect 1600 229 1620 249
rect 1640 229 1660 249
rect 1680 229 1700 249
rect 1720 229 1740 249
rect 1760 229 1780 249
rect 1800 229 1820 249
rect 1840 229 1860 249
rect 1880 229 1900 249
rect 1920 229 1940 249
rect 1960 229 1980 249
rect 2000 229 2020 249
rect 2040 229 2060 249
rect 2080 229 2100 249
rect 2120 229 2140 249
rect 2160 229 2180 249
rect 2200 229 2220 249
rect 2240 229 2260 249
rect 2280 229 2300 249
rect 2320 229 2340 249
rect 2360 229 2380 249
rect 2400 229 2420 249
rect 2440 229 2460 249
rect 2480 229 2500 249
rect 2520 229 2540 249
rect 2560 229 2580 249
rect 2600 229 2620 249
rect 2640 229 2660 249
rect 200 147 220 167
rect 240 147 260 167
rect 280 147 300 167
rect 320 147 340 167
rect 360 147 380 167
rect 400 147 420 167
rect 440 147 460 167
rect 480 147 500 167
rect 520 147 540 167
rect 560 147 580 167
rect 600 147 620 167
rect 640 147 660 167
rect 680 147 700 167
rect 720 147 740 167
rect 760 147 780 167
rect 800 147 820 167
rect 840 147 860 167
rect 880 147 900 167
rect 920 147 940 167
rect 960 147 980 167
rect 1000 147 1020 167
rect 1040 147 1060 167
rect 1080 147 1100 167
rect 1120 147 1140 167
rect 1160 147 1180 167
rect 1200 147 1220 167
rect 1240 147 1260 167
rect 1280 147 1300 167
rect 1320 147 1340 167
rect 1360 147 1380 167
rect 1400 147 1420 167
rect 1440 147 1460 167
rect 1480 147 1500 167
rect 1520 147 1540 167
rect 1560 147 1580 167
rect 1600 147 1620 167
rect 1640 147 1660 167
rect 1680 147 1700 167
rect 1720 147 1740 167
rect 1760 147 1780 167
rect 1800 147 1820 167
rect 1840 147 1860 167
rect 1880 147 1900 167
rect 1920 147 1940 167
rect 1960 147 1980 167
rect 2000 147 2020 167
rect 2040 147 2060 167
rect 2080 147 2100 167
rect 2120 147 2140 167
rect 2160 147 2180 167
rect 2200 147 2220 167
rect 2240 147 2260 167
rect 2280 147 2300 167
rect 2320 147 2340 167
rect 2360 147 2380 167
rect 2400 147 2420 167
rect 2440 147 2460 167
rect 2480 147 2500 167
rect 2520 147 2540 167
rect 2560 147 2580 167
rect 2600 147 2620 167
rect 2640 147 2660 167
rect 200 65 220 85
rect 240 65 260 85
rect 280 65 300 85
rect 320 65 340 85
rect 360 65 380 85
rect 400 65 420 85
rect 440 65 460 85
rect 480 65 500 85
rect 520 65 540 85
rect 560 65 580 85
rect 600 65 620 85
rect 640 65 660 85
rect 680 65 700 85
rect 720 65 740 85
rect 760 65 780 85
rect 800 65 820 85
rect 840 65 860 85
rect 880 65 900 85
rect 920 65 940 85
rect 960 65 980 85
rect 1000 65 1020 85
rect 1040 65 1060 85
rect 1080 65 1100 85
rect 1120 65 1140 85
rect 1160 65 1180 85
rect 1200 65 1220 85
rect 1240 65 1260 85
rect 1280 65 1300 85
rect 1320 65 1340 85
rect 1360 65 1380 85
rect 1400 65 1420 85
rect 1440 65 1460 85
rect 1480 65 1500 85
rect 1520 65 1540 85
rect 1560 65 1580 85
rect 1600 65 1620 85
rect 1640 65 1660 85
rect 1680 65 1700 85
rect 1720 65 1740 85
rect 1760 65 1780 85
rect 1800 65 1820 85
rect 1840 65 1860 85
rect 1880 65 1900 85
rect 1920 65 1940 85
rect 1960 65 1980 85
rect 2000 65 2020 85
rect 2040 65 2060 85
rect 2080 65 2100 85
rect 2120 65 2140 85
rect 2160 65 2180 85
rect 2200 65 2220 85
rect 2240 65 2260 85
rect 2280 65 2300 85
rect 2320 65 2340 85
rect 2360 65 2380 85
rect 2400 65 2420 85
rect 2440 65 2460 85
rect 2480 65 2500 85
rect 2520 65 2540 85
rect 2560 65 2580 85
rect 2600 65 2620 85
rect 2640 65 2660 85
rect 120 -235 140 -215
rect 160 -235 180 -215
rect 200 -235 220 -215
rect 240 -235 260 -215
rect 280 -235 300 -215
rect 320 -235 340 -215
rect 360 -235 380 -215
rect 400 -235 420 -215
rect 440 -235 460 -215
rect 480 -235 500 -215
rect 520 -235 540 -215
rect 560 -235 580 -215
rect 600 -235 620 -215
rect 640 -235 660 -215
rect 680 -235 700 -215
rect 720 -235 740 -215
rect 760 -235 780 -215
rect 800 -235 820 -215
rect 840 -235 860 -215
rect 880 -235 900 -215
rect 920 -235 940 -215
rect 960 -235 980 -215
rect 1000 -235 1020 -215
rect 1040 -235 1060 -215
rect 1080 -235 1100 -215
rect 1120 -235 1140 -215
rect 1160 -235 1180 -215
rect 1200 -235 1220 -215
rect 1240 -235 1260 -215
rect 1280 -235 1300 -215
rect 1320 -235 1340 -215
rect 1360 -235 1380 -215
rect 1400 -235 1420 -215
rect 1440 -235 1460 -215
rect 1480 -235 1500 -215
rect 1520 -235 1540 -215
rect 1560 -235 1580 -215
rect 1600 -235 1620 -215
rect 1640 -235 1660 -215
rect 1680 -235 1700 -215
rect 1720 -235 1740 -215
rect 1760 -235 1780 -215
rect 1800 -235 1820 -215
rect 1840 -235 1860 -215
rect 1880 -235 1900 -215
rect 1920 -235 1940 -215
rect 1960 -235 1980 -215
rect 2000 -235 2020 -215
rect 2040 -235 2060 -215
rect 2080 -235 2100 -215
rect 2120 -235 2140 -215
rect 2160 -235 2180 -215
rect 2200 -235 2220 -215
rect 2240 -235 2260 -215
rect 2280 -235 2300 -215
rect 2320 -235 2340 -215
rect 2360 -235 2380 -215
rect 2400 -235 2420 -215
rect 2440 -235 2460 -215
rect 2480 -235 2500 -215
rect 2520 -235 2540 -215
rect 2560 -235 2590 -215
rect 120 -330 140 -310
rect 160 -330 180 -310
rect 200 -330 220 -310
rect 240 -330 260 -310
rect 280 -330 300 -310
rect 320 -330 340 -310
rect 360 -330 380 -310
rect 400 -330 420 -310
rect 440 -330 460 -310
rect 480 -330 500 -310
rect 520 -330 540 -310
rect 560 -330 580 -310
rect 600 -330 620 -310
rect 640 -330 660 -310
rect 680 -330 700 -310
rect 720 -330 740 -310
rect 760 -330 780 -310
rect 800 -330 820 -310
rect 840 -330 860 -310
rect 880 -330 900 -310
rect 920 -330 940 -310
rect 960 -330 980 -310
rect 1000 -330 1020 -310
rect 1040 -330 1060 -310
rect 1080 -330 1100 -310
rect 1120 -330 1140 -310
rect 1160 -330 1180 -310
rect 1200 -330 1220 -310
rect 1240 -330 1260 -310
rect 1280 -330 1300 -310
rect 1320 -330 1340 -310
rect 1360 -330 1380 -310
rect 1400 -330 1420 -310
rect 1440 -330 1460 -310
rect 1480 -330 1500 -310
rect 1520 -330 1540 -310
rect 1560 -330 1580 -310
rect 1600 -330 1620 -310
rect 1640 -330 1660 -310
rect 1680 -330 1700 -310
rect 1720 -330 1740 -310
rect 1760 -330 1780 -310
rect 1800 -330 1820 -310
rect 1840 -330 1860 -310
rect 1880 -330 1900 -310
rect 1920 -330 1940 -310
rect 1960 -330 1980 -310
rect 2000 -330 2020 -310
rect 2040 -330 2060 -310
rect 2080 -330 2100 -310
rect 2120 -330 2140 -310
rect 2160 -330 2180 -310
rect 2200 -330 2220 -310
rect 2240 -330 2260 -310
rect 2280 -330 2300 -310
rect 2320 -330 2340 -310
rect 2360 -330 2380 -310
rect 2400 -330 2420 -310
rect 2440 -330 2460 -310
rect 2480 -330 2500 -310
rect 2520 -330 2540 -310
rect 2560 -330 2590 -310
rect 120 -425 140 -405
rect 160 -425 180 -405
rect 200 -425 220 -405
rect 240 -425 260 -405
rect 280 -425 300 -405
rect 320 -425 340 -405
rect 360 -425 380 -405
rect 400 -425 420 -405
rect 440 -425 460 -405
rect 480 -425 500 -405
rect 520 -425 540 -405
rect 560 -425 580 -405
rect 600 -425 620 -405
rect 640 -425 660 -405
rect 680 -425 700 -405
rect 720 -425 740 -405
rect 760 -425 780 -405
rect 800 -425 820 -405
rect 840 -425 860 -405
rect 880 -425 900 -405
rect 920 -425 940 -405
rect 960 -425 980 -405
rect 1000 -425 1020 -405
rect 1040 -425 1060 -405
rect 1080 -425 1100 -405
rect 1120 -425 1140 -405
rect 1160 -425 1180 -405
rect 1200 -425 1220 -405
rect 1240 -425 1260 -405
rect 1280 -425 1300 -405
rect 1320 -425 1340 -405
rect 1360 -425 1380 -405
rect 1400 -425 1420 -405
rect 1440 -425 1460 -405
rect 1480 -425 1500 -405
rect 1520 -425 1540 -405
rect 1560 -425 1580 -405
rect 1600 -425 1620 -405
rect 1640 -425 1660 -405
rect 1680 -425 1700 -405
rect 1720 -425 1740 -405
rect 1760 -425 1780 -405
rect 1800 -425 1820 -405
rect 1840 -425 1860 -405
rect 1880 -425 1900 -405
rect 1920 -425 1940 -405
rect 1960 -425 1980 -405
rect 2000 -425 2020 -405
rect 2040 -425 2060 -405
rect 2080 -425 2100 -405
rect 2120 -425 2140 -405
rect 2160 -425 2180 -405
rect 2200 -425 2220 -405
rect 2240 -425 2260 -405
rect 2280 -425 2300 -405
rect 2320 -425 2340 -405
rect 2360 -425 2380 -405
rect 2400 -425 2420 -405
rect 2440 -425 2460 -405
rect 2480 -425 2500 -405
rect 2520 -425 2540 -405
rect 2560 -425 2590 -405
rect 120 -520 140 -500
rect 160 -520 180 -500
rect 200 -520 220 -500
rect 240 -520 260 -500
rect 280 -520 300 -500
rect 320 -520 340 -500
rect 360 -520 380 -500
rect 400 -520 420 -500
rect 440 -520 460 -500
rect 480 -520 500 -500
rect 520 -520 540 -500
rect 560 -520 580 -500
rect 600 -520 620 -500
rect 640 -520 660 -500
rect 680 -520 700 -500
rect 720 -520 740 -500
rect 760 -520 780 -500
rect 800 -520 820 -500
rect 840 -520 860 -500
rect 880 -520 900 -500
rect 920 -520 940 -500
rect 960 -520 980 -500
rect 1000 -520 1020 -500
rect 1040 -520 1060 -500
rect 1080 -520 1100 -500
rect 1120 -520 1140 -500
rect 1160 -520 1180 -500
rect 1200 -520 1220 -500
rect 1240 -520 1260 -500
rect 1280 -520 1300 -500
rect 1320 -520 1340 -500
rect 1360 -520 1380 -500
rect 1400 -520 1420 -500
rect 1440 -520 1460 -500
rect 1480 -520 1500 -500
rect 1520 -520 1540 -500
rect 1560 -520 1580 -500
rect 1600 -520 1620 -500
rect 1640 -520 1660 -500
rect 1680 -520 1700 -500
rect 1720 -520 1740 -500
rect 1760 -520 1780 -500
rect 1800 -520 1820 -500
rect 1840 -520 1860 -500
rect 1880 -520 1900 -500
rect 1920 -520 1940 -500
rect 1960 -520 1980 -500
rect 2000 -520 2020 -500
rect 2040 -520 2060 -500
rect 2080 -520 2100 -500
rect 2120 -520 2140 -500
rect 2160 -520 2180 -500
rect 2200 -520 2220 -500
rect 2240 -520 2260 -500
rect 2280 -520 2300 -500
rect 2320 -520 2340 -500
rect 2360 -520 2380 -500
rect 2400 -520 2420 -500
rect 2440 -520 2460 -500
rect 2480 -520 2500 -500
rect 2520 -520 2540 -500
rect 2560 -520 2590 -500
rect 120 -615 140 -595
rect 160 -615 180 -595
rect 200 -615 220 -595
rect 240 -615 260 -595
rect 280 -615 300 -595
rect 320 -615 340 -595
rect 360 -615 380 -595
rect 400 -615 420 -595
rect 440 -615 460 -595
rect 480 -615 500 -595
rect 520 -615 540 -595
rect 560 -615 580 -595
rect 600 -615 620 -595
rect 640 -615 660 -595
rect 680 -615 700 -595
rect 720 -615 740 -595
rect 760 -615 780 -595
rect 800 -615 820 -595
rect 840 -615 860 -595
rect 880 -615 900 -595
rect 920 -615 940 -595
rect 960 -615 980 -595
rect 1000 -615 1020 -595
rect 1040 -615 1060 -595
rect 1080 -615 1100 -595
rect 1120 -615 1140 -595
rect 1160 -615 1180 -595
rect 1200 -615 1220 -595
rect 1240 -615 1260 -595
rect 1280 -615 1300 -595
rect 1320 -615 1340 -595
rect 1360 -615 1380 -595
rect 1400 -615 1420 -595
rect 1440 -615 1460 -595
rect 1480 -615 1500 -595
rect 1520 -615 1540 -595
rect 1560 -615 1580 -595
rect 1600 -615 1620 -595
rect 1640 -615 1660 -595
rect 1680 -615 1700 -595
rect 1720 -615 1740 -595
rect 1760 -615 1780 -595
rect 1800 -615 1820 -595
rect 1840 -615 1860 -595
rect 1880 -615 1900 -595
rect 1920 -615 1940 -595
rect 1960 -615 1980 -595
rect 2000 -615 2020 -595
rect 2040 -615 2060 -595
rect 2080 -615 2100 -595
rect 2120 -615 2140 -595
rect 2160 -615 2180 -595
rect 2200 -615 2220 -595
rect 2240 -615 2260 -595
rect 2280 -615 2300 -595
rect 2320 -615 2340 -595
rect 2360 -615 2380 -595
rect 2400 -615 2420 -595
rect 2440 -615 2460 -595
rect 2480 -615 2500 -595
rect 2520 -615 2540 -595
rect 2560 -615 2590 -595
rect 120 -710 140 -690
rect 160 -710 180 -690
rect 200 -710 220 -690
rect 240 -710 260 -690
rect 280 -710 300 -690
rect 320 -710 340 -690
rect 360 -710 380 -690
rect 400 -710 420 -690
rect 440 -710 460 -690
rect 480 -710 500 -690
rect 520 -710 540 -690
rect 560 -710 580 -690
rect 600 -710 620 -690
rect 640 -710 660 -690
rect 680 -710 700 -690
rect 720 -710 740 -690
rect 760 -710 780 -690
rect 800 -710 820 -690
rect 840 -710 860 -690
rect 880 -710 900 -690
rect 920 -710 940 -690
rect 960 -710 980 -690
rect 1000 -710 1020 -690
rect 1040 -710 1060 -690
rect 1080 -710 1100 -690
rect 1120 -710 1140 -690
rect 1160 -710 1180 -690
rect 1200 -710 1220 -690
rect 1240 -710 1260 -690
rect 1280 -710 1300 -690
rect 1320 -710 1340 -690
rect 1360 -710 1380 -690
rect 1400 -710 1420 -690
rect 1440 -710 1460 -690
rect 1480 -710 1500 -690
rect 1520 -710 1540 -690
rect 1560 -710 1580 -690
rect 1600 -710 1620 -690
rect 1640 -710 1660 -690
rect 1680 -710 1700 -690
rect 1720 -710 1740 -690
rect 1760 -710 1780 -690
rect 1800 -710 1820 -690
rect 1840 -710 1860 -690
rect 1880 -710 1900 -690
rect 1920 -710 1940 -690
rect 1960 -710 1980 -690
rect 2000 -710 2020 -690
rect 2040 -710 2060 -690
rect 2080 -710 2100 -690
rect 2120 -710 2140 -690
rect 2160 -710 2180 -690
rect 2200 -710 2220 -690
rect 2240 -710 2260 -690
rect 2280 -710 2300 -690
rect 2320 -710 2340 -690
rect 2360 -710 2380 -690
rect 2400 -710 2420 -690
rect 2440 -710 2460 -690
rect 2480 -710 2500 -690
rect 2520 -710 2540 -690
rect 2560 -710 2590 -690
rect 120 -805 140 -785
rect 160 -805 180 -785
rect 200 -805 220 -785
rect 240 -805 260 -785
rect 280 -805 300 -785
rect 320 -805 340 -785
rect 360 -805 380 -785
rect 400 -805 420 -785
rect 440 -805 460 -785
rect 480 -805 500 -785
rect 520 -805 540 -785
rect 560 -805 580 -785
rect 600 -805 620 -785
rect 640 -805 660 -785
rect 680 -805 700 -785
rect 720 -805 740 -785
rect 760 -805 780 -785
rect 800 -805 820 -785
rect 840 -805 860 -785
rect 880 -805 900 -785
rect 920 -805 940 -785
rect 960 -805 980 -785
rect 1000 -805 1020 -785
rect 1040 -805 1060 -785
rect 1080 -805 1100 -785
rect 1120 -805 1140 -785
rect 1160 -805 1180 -785
rect 1200 -805 1220 -785
rect 1240 -805 1260 -785
rect 1280 -805 1300 -785
rect 1320 -805 1340 -785
rect 1360 -805 1380 -785
rect 1400 -805 1420 -785
rect 1440 -805 1460 -785
rect 1480 -805 1500 -785
rect 1520 -805 1540 -785
rect 1560 -805 1580 -785
rect 1600 -805 1620 -785
rect 1640 -805 1660 -785
rect 1680 -805 1700 -785
rect 1720 -805 1740 -785
rect 1760 -805 1780 -785
rect 1800 -805 1820 -785
rect 1840 -805 1860 -785
rect 1880 -805 1900 -785
rect 1920 -805 1940 -785
rect 1960 -805 1980 -785
rect 2000 -805 2020 -785
rect 2040 -805 2060 -785
rect 2080 -805 2100 -785
rect 2120 -805 2140 -785
rect 2160 -805 2180 -785
rect 2200 -805 2220 -785
rect 2240 -805 2260 -785
rect 2280 -805 2300 -785
rect 2320 -805 2340 -785
rect 2360 -805 2380 -785
rect 2400 -805 2420 -785
rect 2440 -805 2460 -785
rect 2480 -805 2500 -785
rect 2520 -805 2540 -785
rect 2560 -805 2590 -785
rect 120 -900 140 -880
rect 160 -900 180 -880
rect 200 -900 220 -880
rect 240 -900 260 -880
rect 280 -900 300 -880
rect 320 -900 340 -880
rect 360 -900 380 -880
rect 400 -900 420 -880
rect 440 -900 460 -880
rect 480 -900 500 -880
rect 520 -900 540 -880
rect 560 -900 580 -880
rect 600 -900 620 -880
rect 640 -900 660 -880
rect 680 -900 700 -880
rect 720 -900 740 -880
rect 760 -900 780 -880
rect 800 -900 820 -880
rect 840 -900 860 -880
rect 880 -900 900 -880
rect 920 -900 940 -880
rect 960 -900 980 -880
rect 1000 -900 1020 -880
rect 1040 -900 1060 -880
rect 1080 -900 1100 -880
rect 1120 -900 1140 -880
rect 1160 -900 1180 -880
rect 1200 -900 1220 -880
rect 1240 -900 1260 -880
rect 1280 -900 1300 -880
rect 1320 -900 1340 -880
rect 1360 -900 1380 -880
rect 1400 -900 1420 -880
rect 1440 -900 1460 -880
rect 1480 -900 1500 -880
rect 1520 -900 1540 -880
rect 1560 -900 1580 -880
rect 1600 -900 1620 -880
rect 1640 -900 1660 -880
rect 1680 -900 1700 -880
rect 1720 -900 1740 -880
rect 1760 -900 1780 -880
rect 1800 -900 1820 -880
rect 1840 -900 1860 -880
rect 1880 -900 1900 -880
rect 1920 -900 1940 -880
rect 1960 -900 1980 -880
rect 2000 -900 2020 -880
rect 2040 -900 2060 -880
rect 2080 -900 2100 -880
rect 2120 -900 2140 -880
rect 2160 -900 2180 -880
rect 2200 -900 2220 -880
rect 2240 -900 2260 -880
rect 2280 -900 2300 -880
rect 2320 -900 2340 -880
rect 2360 -900 2380 -880
rect 2400 -900 2420 -880
rect 2440 -900 2460 -880
rect 2480 -900 2500 -880
rect 2520 -900 2540 -880
rect 2560 -900 2590 -880
rect 120 -995 140 -975
rect 160 -995 180 -975
rect 200 -995 220 -975
rect 240 -995 260 -975
rect 280 -995 300 -975
rect 320 -995 340 -975
rect 360 -995 380 -975
rect 400 -995 420 -975
rect 440 -995 460 -975
rect 480 -995 500 -975
rect 520 -995 540 -975
rect 560 -995 580 -975
rect 600 -995 620 -975
rect 640 -995 660 -975
rect 680 -995 700 -975
rect 720 -995 740 -975
rect 760 -995 780 -975
rect 800 -995 820 -975
rect 840 -995 860 -975
rect 880 -995 900 -975
rect 920 -995 940 -975
rect 960 -995 980 -975
rect 1000 -995 1020 -975
rect 1040 -995 1060 -975
rect 1080 -995 1100 -975
rect 1120 -995 1140 -975
rect 1160 -995 1180 -975
rect 1200 -995 1220 -975
rect 1240 -995 1260 -975
rect 1280 -995 1300 -975
rect 1320 -995 1340 -975
rect 1360 -995 1380 -975
rect 1400 -995 1420 -975
rect 1440 -995 1460 -975
rect 1480 -995 1500 -975
rect 1520 -995 1540 -975
rect 1560 -995 1580 -975
rect 1600 -995 1620 -975
rect 1640 -995 1660 -975
rect 1680 -995 1700 -975
rect 1720 -995 1740 -975
rect 1760 -995 1780 -975
rect 1800 -995 1820 -975
rect 1840 -995 1860 -975
rect 1880 -995 1900 -975
rect 1920 -995 1940 -975
rect 1960 -995 1980 -975
rect 2000 -995 2020 -975
rect 2040 -995 2060 -975
rect 2080 -995 2100 -975
rect 2120 -995 2140 -975
rect 2160 -995 2180 -975
rect 2200 -995 2220 -975
rect 2240 -995 2260 -975
rect 2280 -995 2300 -975
rect 2320 -995 2340 -975
rect 2360 -995 2380 -975
rect 2400 -995 2420 -975
rect 2440 -995 2460 -975
rect 2480 -995 2500 -975
rect 2520 -995 2540 -975
rect 2560 -995 2590 -975
rect 120 -1090 140 -1070
rect 160 -1090 180 -1070
rect 200 -1090 220 -1070
rect 240 -1090 260 -1070
rect 280 -1090 300 -1070
rect 320 -1090 340 -1070
rect 360 -1090 380 -1070
rect 400 -1090 420 -1070
rect 440 -1090 460 -1070
rect 480 -1090 500 -1070
rect 520 -1090 540 -1070
rect 560 -1090 580 -1070
rect 600 -1090 620 -1070
rect 640 -1090 660 -1070
rect 680 -1090 700 -1070
rect 720 -1090 740 -1070
rect 760 -1090 780 -1070
rect 800 -1090 820 -1070
rect 840 -1090 860 -1070
rect 880 -1090 900 -1070
rect 920 -1090 940 -1070
rect 960 -1090 980 -1070
rect 1000 -1090 1020 -1070
rect 1040 -1090 1060 -1070
rect 1080 -1090 1100 -1070
rect 1120 -1090 1140 -1070
rect 1160 -1090 1180 -1070
rect 1200 -1090 1220 -1070
rect 1240 -1090 1260 -1070
rect 1280 -1090 1300 -1070
rect 1320 -1090 1340 -1070
rect 1360 -1090 1380 -1070
rect 1400 -1090 1420 -1070
rect 1440 -1090 1460 -1070
rect 1480 -1090 1500 -1070
rect 1520 -1090 1540 -1070
rect 1560 -1090 1580 -1070
rect 1600 -1090 1620 -1070
rect 1640 -1090 1660 -1070
rect 1680 -1090 1700 -1070
rect 1720 -1090 1740 -1070
rect 1760 -1090 1780 -1070
rect 1800 -1090 1820 -1070
rect 1840 -1090 1860 -1070
rect 1880 -1090 1900 -1070
rect 1920 -1090 1940 -1070
rect 1960 -1090 1980 -1070
rect 2000 -1090 2020 -1070
rect 2040 -1090 2060 -1070
rect 2080 -1090 2100 -1070
rect 2120 -1090 2140 -1070
rect 2160 -1090 2180 -1070
rect 2200 -1090 2220 -1070
rect 2240 -1090 2260 -1070
rect 2280 -1090 2300 -1070
rect 2320 -1090 2340 -1070
rect 2360 -1090 2380 -1070
rect 2400 -1090 2420 -1070
rect 2440 -1090 2460 -1070
rect 2480 -1090 2500 -1070
rect 2520 -1090 2540 -1070
rect 2560 -1090 2590 -1070
rect 120 -1185 140 -1165
rect 160 -1185 180 -1165
rect 200 -1185 220 -1165
rect 240 -1185 260 -1165
rect 280 -1185 300 -1165
rect 320 -1185 340 -1165
rect 360 -1185 380 -1165
rect 400 -1185 420 -1165
rect 440 -1185 460 -1165
rect 480 -1185 500 -1165
rect 520 -1185 540 -1165
rect 560 -1185 580 -1165
rect 600 -1185 620 -1165
rect 640 -1185 660 -1165
rect 680 -1185 700 -1165
rect 720 -1185 740 -1165
rect 760 -1185 780 -1165
rect 800 -1185 820 -1165
rect 840 -1185 860 -1165
rect 880 -1185 900 -1165
rect 920 -1185 940 -1165
rect 960 -1185 980 -1165
rect 1000 -1185 1020 -1165
rect 1040 -1185 1060 -1165
rect 1080 -1185 1100 -1165
rect 1120 -1185 1140 -1165
rect 1160 -1185 1180 -1165
rect 1200 -1185 1220 -1165
rect 1240 -1185 1260 -1165
rect 1280 -1185 1300 -1165
rect 1320 -1185 1340 -1165
rect 1360 -1185 1380 -1165
rect 1400 -1185 1420 -1165
rect 1440 -1185 1460 -1165
rect 1480 -1185 1500 -1165
rect 1520 -1185 1540 -1165
rect 1560 -1185 1580 -1165
rect 1600 -1185 1620 -1165
rect 1640 -1185 1660 -1165
rect 1680 -1185 1700 -1165
rect 1720 -1185 1740 -1165
rect 1760 -1185 1780 -1165
rect 1800 -1185 1820 -1165
rect 1840 -1185 1860 -1165
rect 1880 -1185 1900 -1165
rect 1920 -1185 1940 -1165
rect 1960 -1185 1980 -1165
rect 2000 -1185 2020 -1165
rect 2040 -1185 2060 -1165
rect 2080 -1185 2100 -1165
rect 2120 -1185 2140 -1165
rect 2160 -1185 2180 -1165
rect 2200 -1185 2220 -1165
rect 2240 -1185 2260 -1165
rect 2280 -1185 2300 -1165
rect 2320 -1185 2340 -1165
rect 2360 -1185 2380 -1165
rect 2400 -1185 2420 -1165
rect 2440 -1185 2460 -1165
rect 2480 -1185 2500 -1165
rect 2520 -1185 2540 -1165
rect 2560 -1185 2590 -1165
rect 120 -1280 140 -1260
rect 160 -1280 180 -1260
rect 200 -1280 220 -1260
rect 240 -1280 260 -1260
rect 280 -1280 300 -1260
rect 320 -1280 340 -1260
rect 360 -1280 380 -1260
rect 400 -1280 420 -1260
rect 440 -1280 460 -1260
rect 480 -1280 500 -1260
rect 520 -1280 540 -1260
rect 560 -1280 580 -1260
rect 600 -1280 620 -1260
rect 640 -1280 660 -1260
rect 680 -1280 700 -1260
rect 720 -1280 740 -1260
rect 760 -1280 780 -1260
rect 800 -1280 820 -1260
rect 840 -1280 860 -1260
rect 880 -1280 900 -1260
rect 920 -1280 940 -1260
rect 960 -1280 980 -1260
rect 1000 -1280 1020 -1260
rect 1040 -1280 1060 -1260
rect 1080 -1280 1100 -1260
rect 1120 -1280 1140 -1260
rect 1160 -1280 1180 -1260
rect 1200 -1280 1220 -1260
rect 1240 -1280 1260 -1260
rect 1280 -1280 1300 -1260
rect 1320 -1280 1340 -1260
rect 1360 -1280 1380 -1260
rect 1400 -1280 1420 -1260
rect 1440 -1280 1460 -1260
rect 1480 -1280 1500 -1260
rect 1520 -1280 1540 -1260
rect 1560 -1280 1580 -1260
rect 1600 -1280 1620 -1260
rect 1640 -1280 1660 -1260
rect 1680 -1280 1700 -1260
rect 1720 -1280 1740 -1260
rect 1760 -1280 1780 -1260
rect 1800 -1280 1820 -1260
rect 1840 -1280 1860 -1260
rect 1880 -1280 1900 -1260
rect 1920 -1280 1940 -1260
rect 1960 -1280 1980 -1260
rect 2000 -1280 2020 -1260
rect 2040 -1280 2060 -1260
rect 2080 -1280 2100 -1260
rect 2120 -1280 2140 -1260
rect 2160 -1280 2180 -1260
rect 2200 -1280 2220 -1260
rect 2240 -1280 2260 -1260
rect 2280 -1280 2300 -1260
rect 2320 -1280 2340 -1260
rect 2360 -1280 2380 -1260
rect 2400 -1280 2420 -1260
rect 2440 -1280 2460 -1260
rect 2480 -1280 2500 -1260
rect 2520 -1280 2540 -1260
rect 2560 -1280 2590 -1260
rect 120 -1375 140 -1355
rect 160 -1375 180 -1355
rect 200 -1375 220 -1355
rect 240 -1375 260 -1355
rect 280 -1375 300 -1355
rect 320 -1375 340 -1355
rect 360 -1375 380 -1355
rect 400 -1375 420 -1355
rect 440 -1375 460 -1355
rect 480 -1375 500 -1355
rect 520 -1375 540 -1355
rect 560 -1375 580 -1355
rect 600 -1375 620 -1355
rect 640 -1375 660 -1355
rect 680 -1375 700 -1355
rect 720 -1375 740 -1355
rect 760 -1375 780 -1355
rect 800 -1375 820 -1355
rect 840 -1375 860 -1355
rect 880 -1375 900 -1355
rect 920 -1375 940 -1355
rect 960 -1375 980 -1355
rect 1000 -1375 1020 -1355
rect 1040 -1375 1060 -1355
rect 1080 -1375 1100 -1355
rect 1120 -1375 1140 -1355
rect 1160 -1375 1180 -1355
rect 1200 -1375 1220 -1355
rect 1240 -1375 1260 -1355
rect 1280 -1375 1300 -1355
rect 1320 -1375 1340 -1355
rect 1360 -1375 1380 -1355
rect 1400 -1375 1420 -1355
rect 1440 -1375 1460 -1355
rect 1480 -1375 1500 -1355
rect 1520 -1375 1540 -1355
rect 1560 -1375 1580 -1355
rect 1600 -1375 1620 -1355
rect 1640 -1375 1660 -1355
rect 1680 -1375 1700 -1355
rect 1720 -1375 1740 -1355
rect 1760 -1375 1780 -1355
rect 1800 -1375 1820 -1355
rect 1840 -1375 1860 -1355
rect 1880 -1375 1900 -1355
rect 1920 -1375 1940 -1355
rect 1960 -1375 1980 -1355
rect 2000 -1375 2020 -1355
rect 2040 -1375 2060 -1355
rect 2080 -1375 2100 -1355
rect 2120 -1375 2140 -1355
rect 2160 -1375 2180 -1355
rect 2200 -1375 2220 -1355
rect 2240 -1375 2260 -1355
rect 2280 -1375 2300 -1355
rect 2320 -1375 2340 -1355
rect 2360 -1375 2380 -1355
rect 2400 -1375 2420 -1355
rect 2440 -1375 2460 -1355
rect 2480 -1375 2500 -1355
rect 2520 -1375 2540 -1355
rect 2560 -1375 2590 -1355
rect 120 -1470 140 -1450
rect 160 -1470 180 -1450
rect 200 -1470 220 -1450
rect 240 -1470 260 -1450
rect 280 -1470 300 -1450
rect 320 -1470 340 -1450
rect 360 -1470 380 -1450
rect 400 -1470 420 -1450
rect 440 -1470 460 -1450
rect 480 -1470 500 -1450
rect 520 -1470 540 -1450
rect 560 -1470 580 -1450
rect 600 -1470 620 -1450
rect 640 -1470 660 -1450
rect 680 -1470 700 -1450
rect 720 -1470 740 -1450
rect 760 -1470 780 -1450
rect 800 -1470 820 -1450
rect 840 -1470 860 -1450
rect 880 -1470 900 -1450
rect 920 -1470 940 -1450
rect 960 -1470 980 -1450
rect 1000 -1470 1020 -1450
rect 1040 -1470 1060 -1450
rect 1080 -1470 1100 -1450
rect 1120 -1470 1140 -1450
rect 1160 -1470 1180 -1450
rect 1200 -1470 1220 -1450
rect 1240 -1470 1260 -1450
rect 1280 -1470 1300 -1450
rect 1320 -1470 1340 -1450
rect 1360 -1470 1380 -1450
rect 1400 -1470 1420 -1450
rect 1440 -1470 1460 -1450
rect 1480 -1470 1500 -1450
rect 1520 -1470 1540 -1450
rect 1560 -1470 1580 -1450
rect 1600 -1470 1620 -1450
rect 1640 -1470 1660 -1450
rect 1680 -1470 1700 -1450
rect 1720 -1470 1740 -1450
rect 1760 -1470 1780 -1450
rect 1800 -1470 1820 -1450
rect 1840 -1470 1860 -1450
rect 1880 -1470 1900 -1450
rect 1920 -1470 1940 -1450
rect 1960 -1470 1980 -1450
rect 2000 -1470 2020 -1450
rect 2040 -1470 2060 -1450
rect 2080 -1470 2100 -1450
rect 2120 -1470 2140 -1450
rect 2160 -1470 2180 -1450
rect 2200 -1470 2220 -1450
rect 2240 -1470 2260 -1450
rect 2280 -1470 2300 -1450
rect 2320 -1470 2340 -1450
rect 2360 -1470 2380 -1450
rect 2400 -1470 2420 -1450
rect 2440 -1470 2460 -1450
rect 2480 -1470 2500 -1450
rect 2520 -1470 2540 -1450
rect 2560 -1470 2590 -1450
rect 120 -1565 140 -1545
rect 160 -1565 180 -1545
rect 200 -1565 220 -1545
rect 240 -1565 260 -1545
rect 280 -1565 300 -1545
rect 320 -1565 340 -1545
rect 360 -1565 380 -1545
rect 400 -1565 420 -1545
rect 440 -1565 460 -1545
rect 480 -1565 500 -1545
rect 520 -1565 540 -1545
rect 560 -1565 580 -1545
rect 600 -1565 620 -1545
rect 640 -1565 660 -1545
rect 680 -1565 700 -1545
rect 720 -1565 740 -1545
rect 760 -1565 780 -1545
rect 800 -1565 820 -1545
rect 840 -1565 860 -1545
rect 880 -1565 900 -1545
rect 920 -1565 940 -1545
rect 960 -1565 980 -1545
rect 1000 -1565 1020 -1545
rect 1040 -1565 1060 -1545
rect 1080 -1565 1100 -1545
rect 1120 -1565 1140 -1545
rect 1160 -1565 1180 -1545
rect 1200 -1565 1220 -1545
rect 1240 -1565 1260 -1545
rect 1280 -1565 1300 -1545
rect 1320 -1565 1340 -1545
rect 1360 -1565 1380 -1545
rect 1400 -1565 1420 -1545
rect 1440 -1565 1460 -1545
rect 1480 -1565 1500 -1545
rect 1520 -1565 1540 -1545
rect 1560 -1565 1580 -1545
rect 1600 -1565 1620 -1545
rect 1640 -1565 1660 -1545
rect 1680 -1565 1700 -1545
rect 1720 -1565 1740 -1545
rect 1760 -1565 1780 -1545
rect 1800 -1565 1820 -1545
rect 1840 -1565 1860 -1545
rect 1880 -1565 1900 -1545
rect 1920 -1565 1940 -1545
rect 1960 -1565 1980 -1545
rect 2000 -1565 2020 -1545
rect 2040 -1565 2060 -1545
rect 2080 -1565 2100 -1545
rect 2120 -1565 2140 -1545
rect 2160 -1565 2180 -1545
rect 2200 -1565 2220 -1545
rect 2240 -1565 2260 -1545
rect 2280 -1565 2300 -1545
rect 2320 -1565 2340 -1545
rect 2360 -1565 2380 -1545
rect 2400 -1565 2420 -1545
rect 2440 -1565 2460 -1545
rect 2480 -1565 2500 -1545
rect 2520 -1565 2540 -1545
rect 2560 -1565 2590 -1545
rect 120 -1660 140 -1640
rect 160 -1660 180 -1640
rect 200 -1660 220 -1640
rect 240 -1660 260 -1640
rect 280 -1660 300 -1640
rect 320 -1660 340 -1640
rect 360 -1660 380 -1640
rect 400 -1660 420 -1640
rect 440 -1660 460 -1640
rect 480 -1660 500 -1640
rect 520 -1660 540 -1640
rect 560 -1660 580 -1640
rect 600 -1660 620 -1640
rect 640 -1660 660 -1640
rect 680 -1660 700 -1640
rect 720 -1660 740 -1640
rect 760 -1660 780 -1640
rect 800 -1660 820 -1640
rect 840 -1660 860 -1640
rect 880 -1660 900 -1640
rect 920 -1660 940 -1640
rect 960 -1660 980 -1640
rect 1000 -1660 1020 -1640
rect 1040 -1660 1060 -1640
rect 1080 -1660 1100 -1640
rect 1120 -1660 1140 -1640
rect 1160 -1660 1180 -1640
rect 1200 -1660 1220 -1640
rect 1240 -1660 1260 -1640
rect 1280 -1660 1300 -1640
rect 1320 -1660 1340 -1640
rect 1360 -1660 1380 -1640
rect 1400 -1660 1420 -1640
rect 1440 -1660 1460 -1640
rect 1480 -1660 1500 -1640
rect 1520 -1660 1540 -1640
rect 1560 -1660 1580 -1640
rect 1600 -1660 1620 -1640
rect 1640 -1660 1660 -1640
rect 1680 -1660 1700 -1640
rect 1720 -1660 1740 -1640
rect 1760 -1660 1780 -1640
rect 1800 -1660 1820 -1640
rect 1840 -1660 1860 -1640
rect 1880 -1660 1900 -1640
rect 1920 -1660 1940 -1640
rect 1960 -1660 1980 -1640
rect 2000 -1660 2020 -1640
rect 2040 -1660 2060 -1640
rect 2080 -1660 2100 -1640
rect 2120 -1660 2140 -1640
rect 2160 -1660 2180 -1640
rect 2200 -1660 2220 -1640
rect 2240 -1660 2260 -1640
rect 2280 -1660 2300 -1640
rect 2320 -1660 2340 -1640
rect 2360 -1660 2380 -1640
rect 2400 -1660 2420 -1640
rect 2440 -1660 2460 -1640
rect 2480 -1660 2500 -1640
rect 2520 -1660 2540 -1640
rect 2560 -1660 2590 -1640
rect 120 -1755 140 -1735
rect 160 -1755 180 -1735
rect 200 -1755 220 -1735
rect 240 -1755 260 -1735
rect 280 -1755 300 -1735
rect 320 -1755 340 -1735
rect 360 -1755 380 -1735
rect 400 -1755 420 -1735
rect 440 -1755 460 -1735
rect 480 -1755 500 -1735
rect 520 -1755 540 -1735
rect 560 -1755 580 -1735
rect 600 -1755 620 -1735
rect 640 -1755 660 -1735
rect 680 -1755 700 -1735
rect 720 -1755 740 -1735
rect 760 -1755 780 -1735
rect 800 -1755 820 -1735
rect 840 -1755 860 -1735
rect 880 -1755 900 -1735
rect 920 -1755 940 -1735
rect 960 -1755 980 -1735
rect 1000 -1755 1020 -1735
rect 1040 -1755 1060 -1735
rect 1080 -1755 1100 -1735
rect 1120 -1755 1140 -1735
rect 1160 -1755 1180 -1735
rect 1200 -1755 1220 -1735
rect 1240 -1755 1260 -1735
rect 1280 -1755 1300 -1735
rect 1320 -1755 1340 -1735
rect 1360 -1755 1380 -1735
rect 1400 -1755 1420 -1735
rect 1440 -1755 1460 -1735
rect 1480 -1755 1500 -1735
rect 1520 -1755 1540 -1735
rect 1560 -1755 1580 -1735
rect 1600 -1755 1620 -1735
rect 1640 -1755 1660 -1735
rect 1680 -1755 1700 -1735
rect 1720 -1755 1740 -1735
rect 1760 -1755 1780 -1735
rect 1800 -1755 1820 -1735
rect 1840 -1755 1860 -1735
rect 1880 -1755 1900 -1735
rect 1920 -1755 1940 -1735
rect 1960 -1755 1980 -1735
rect 2000 -1755 2020 -1735
rect 2040 -1755 2060 -1735
rect 2080 -1755 2100 -1735
rect 2120 -1755 2140 -1735
rect 2160 -1755 2180 -1735
rect 2200 -1755 2220 -1735
rect 2240 -1755 2260 -1735
rect 2280 -1755 2300 -1735
rect 2320 -1755 2340 -1735
rect 2360 -1755 2380 -1735
rect 2400 -1755 2420 -1735
rect 2440 -1755 2460 -1735
rect 2480 -1755 2500 -1735
rect 2520 -1755 2540 -1735
rect 2560 -1755 2590 -1735
rect 120 -1850 140 -1830
rect 160 -1850 180 -1830
rect 200 -1850 220 -1830
rect 240 -1850 260 -1830
rect 280 -1850 300 -1830
rect 320 -1850 340 -1830
rect 360 -1850 380 -1830
rect 400 -1850 420 -1830
rect 440 -1850 460 -1830
rect 480 -1850 500 -1830
rect 520 -1850 540 -1830
rect 560 -1850 580 -1830
rect 600 -1850 620 -1830
rect 640 -1850 660 -1830
rect 680 -1850 700 -1830
rect 720 -1850 740 -1830
rect 760 -1850 780 -1830
rect 800 -1850 820 -1830
rect 840 -1850 860 -1830
rect 880 -1850 900 -1830
rect 920 -1850 940 -1830
rect 960 -1850 980 -1830
rect 1000 -1850 1020 -1830
rect 1040 -1850 1060 -1830
rect 1080 -1850 1100 -1830
rect 1120 -1850 1140 -1830
rect 1160 -1850 1180 -1830
rect 1200 -1850 1220 -1830
rect 1240 -1850 1260 -1830
rect 1280 -1850 1300 -1830
rect 1320 -1850 1340 -1830
rect 1360 -1850 1380 -1830
rect 1400 -1850 1420 -1830
rect 1440 -1850 1460 -1830
rect 1480 -1850 1500 -1830
rect 1520 -1850 1540 -1830
rect 1560 -1850 1580 -1830
rect 1600 -1850 1620 -1830
rect 1640 -1850 1660 -1830
rect 1680 -1850 1700 -1830
rect 1720 -1850 1740 -1830
rect 1760 -1850 1780 -1830
rect 1800 -1850 1820 -1830
rect 1840 -1850 1860 -1830
rect 1880 -1850 1900 -1830
rect 1920 -1850 1940 -1830
rect 1960 -1850 1980 -1830
rect 2000 -1850 2020 -1830
rect 2040 -1850 2060 -1830
rect 2080 -1850 2100 -1830
rect 2120 -1850 2140 -1830
rect 2160 -1850 2180 -1830
rect 2200 -1850 2220 -1830
rect 2240 -1850 2260 -1830
rect 2280 -1850 2300 -1830
rect 2320 -1850 2340 -1830
rect 2360 -1850 2380 -1830
rect 2400 -1850 2420 -1830
rect 2440 -1850 2460 -1830
rect 2480 -1850 2500 -1830
rect 2520 -1850 2540 -1830
rect 2560 -1850 2590 -1830
rect 120 -1945 140 -1925
rect 160 -1945 180 -1925
rect 200 -1945 220 -1925
rect 240 -1945 260 -1925
rect 280 -1945 300 -1925
rect 320 -1945 340 -1925
rect 360 -1945 380 -1925
rect 400 -1945 420 -1925
rect 440 -1945 460 -1925
rect 480 -1945 500 -1925
rect 520 -1945 540 -1925
rect 560 -1945 580 -1925
rect 600 -1945 620 -1925
rect 640 -1945 660 -1925
rect 680 -1945 700 -1925
rect 720 -1945 740 -1925
rect 760 -1945 780 -1925
rect 800 -1945 820 -1925
rect 840 -1945 860 -1925
rect 880 -1945 900 -1925
rect 920 -1945 940 -1925
rect 960 -1945 980 -1925
rect 1000 -1945 1020 -1925
rect 1040 -1945 1060 -1925
rect 1080 -1945 1100 -1925
rect 1120 -1945 1140 -1925
rect 1160 -1945 1180 -1925
rect 1200 -1945 1220 -1925
rect 1240 -1945 1260 -1925
rect 1280 -1945 1300 -1925
rect 1320 -1945 1340 -1925
rect 1360 -1945 1380 -1925
rect 1400 -1945 1420 -1925
rect 1440 -1945 1460 -1925
rect 1480 -1945 1500 -1925
rect 1520 -1945 1540 -1925
rect 1560 -1945 1580 -1925
rect 1600 -1945 1620 -1925
rect 1640 -1945 1660 -1925
rect 1680 -1945 1700 -1925
rect 1720 -1945 1740 -1925
rect 1760 -1945 1780 -1925
rect 1800 -1945 1820 -1925
rect 1840 -1945 1860 -1925
rect 1880 -1945 1900 -1925
rect 1920 -1945 1940 -1925
rect 1960 -1945 1980 -1925
rect 2000 -1945 2020 -1925
rect 2040 -1945 2060 -1925
rect 2080 -1945 2100 -1925
rect 2120 -1945 2140 -1925
rect 2160 -1945 2180 -1925
rect 2200 -1945 2220 -1925
rect 2240 -1945 2260 -1925
rect 2280 -1945 2300 -1925
rect 2320 -1945 2340 -1925
rect 2360 -1945 2380 -1925
rect 2400 -1945 2420 -1925
rect 2440 -1945 2460 -1925
rect 2480 -1945 2500 -1925
rect 2520 -1945 2540 -1925
rect 2560 -1945 2590 -1925
rect 120 -2040 140 -2020
rect 160 -2040 180 -2020
rect 200 -2040 220 -2020
rect 240 -2040 260 -2020
rect 280 -2040 300 -2020
rect 320 -2040 340 -2020
rect 360 -2040 380 -2020
rect 400 -2040 420 -2020
rect 440 -2040 460 -2020
rect 480 -2040 500 -2020
rect 520 -2040 540 -2020
rect 560 -2040 580 -2020
rect 600 -2040 620 -2020
rect 640 -2040 660 -2020
rect 680 -2040 700 -2020
rect 720 -2040 740 -2020
rect 760 -2040 780 -2020
rect 800 -2040 820 -2020
rect 840 -2040 860 -2020
rect 880 -2040 900 -2020
rect 920 -2040 940 -2020
rect 960 -2040 980 -2020
rect 1000 -2040 1020 -2020
rect 1040 -2040 1060 -2020
rect 1080 -2040 1100 -2020
rect 1120 -2040 1140 -2020
rect 1160 -2040 1180 -2020
rect 1200 -2040 1220 -2020
rect 1240 -2040 1260 -2020
rect 1280 -2040 1300 -2020
rect 1320 -2040 1340 -2020
rect 1360 -2040 1380 -2020
rect 1400 -2040 1420 -2020
rect 1440 -2040 1460 -2020
rect 1480 -2040 1500 -2020
rect 1520 -2040 1540 -2020
rect 1560 -2040 1580 -2020
rect 1600 -2040 1620 -2020
rect 1640 -2040 1660 -2020
rect 1680 -2040 1700 -2020
rect 1720 -2040 1740 -2020
rect 1760 -2040 1780 -2020
rect 1800 -2040 1820 -2020
rect 1840 -2040 1860 -2020
rect 1880 -2040 1900 -2020
rect 1920 -2040 1940 -2020
rect 1960 -2040 1980 -2020
rect 2000 -2040 2020 -2020
rect 2040 -2040 2060 -2020
rect 2080 -2040 2100 -2020
rect 2120 -2040 2140 -2020
rect 2160 -2040 2180 -2020
rect 2200 -2040 2220 -2020
rect 2240 -2040 2260 -2020
rect 2280 -2040 2300 -2020
rect 2320 -2040 2340 -2020
rect 2360 -2040 2380 -2020
rect 2400 -2040 2420 -2020
rect 2440 -2040 2460 -2020
rect 2480 -2040 2500 -2020
rect 2520 -2040 2540 -2020
rect 2560 -2040 2590 -2020
rect 120 -2135 140 -2115
rect 160 -2135 180 -2115
rect 200 -2135 220 -2115
rect 240 -2135 260 -2115
rect 280 -2135 300 -2115
rect 320 -2135 340 -2115
rect 360 -2135 380 -2115
rect 400 -2135 420 -2115
rect 440 -2135 460 -2115
rect 480 -2135 500 -2115
rect 520 -2135 540 -2115
rect 560 -2135 580 -2115
rect 600 -2135 620 -2115
rect 640 -2135 660 -2115
rect 680 -2135 700 -2115
rect 720 -2135 740 -2115
rect 760 -2135 780 -2115
rect 800 -2135 820 -2115
rect 840 -2135 860 -2115
rect 880 -2135 900 -2115
rect 920 -2135 940 -2115
rect 960 -2135 980 -2115
rect 1000 -2135 1020 -2115
rect 1040 -2135 1060 -2115
rect 1080 -2135 1100 -2115
rect 1120 -2135 1140 -2115
rect 1160 -2135 1180 -2115
rect 1200 -2135 1220 -2115
rect 1240 -2135 1260 -2115
rect 1280 -2135 1300 -2115
rect 1320 -2135 1340 -2115
rect 1360 -2135 1380 -2115
rect 1400 -2135 1420 -2115
rect 1440 -2135 1460 -2115
rect 1480 -2135 1500 -2115
rect 1520 -2135 1540 -2115
rect 1560 -2135 1580 -2115
rect 1600 -2135 1620 -2115
rect 1640 -2135 1660 -2115
rect 1680 -2135 1700 -2115
rect 1720 -2135 1740 -2115
rect 1760 -2135 1780 -2115
rect 1800 -2135 1820 -2115
rect 1840 -2135 1860 -2115
rect 1880 -2135 1900 -2115
rect 1920 -2135 1940 -2115
rect 1960 -2135 1980 -2115
rect 2000 -2135 2020 -2115
rect 2040 -2135 2060 -2115
rect 2080 -2135 2100 -2115
rect 2120 -2135 2140 -2115
rect 2160 -2135 2180 -2115
rect 2200 -2135 2220 -2115
rect 2240 -2135 2260 -2115
rect 2280 -2135 2300 -2115
rect 2320 -2135 2340 -2115
rect 2360 -2135 2380 -2115
rect 2400 -2135 2420 -2115
rect 2440 -2135 2460 -2115
rect 2480 -2135 2500 -2115
rect 2520 -2135 2540 -2115
rect 2560 -2135 2590 -2115
rect 120 -2230 140 -2210
rect 160 -2230 180 -2210
rect 200 -2230 220 -2210
rect 240 -2230 260 -2210
rect 280 -2230 300 -2210
rect 320 -2230 340 -2210
rect 360 -2230 380 -2210
rect 400 -2230 420 -2210
rect 440 -2230 460 -2210
rect 480 -2230 500 -2210
rect 520 -2230 540 -2210
rect 560 -2230 580 -2210
rect 600 -2230 620 -2210
rect 640 -2230 660 -2210
rect 680 -2230 700 -2210
rect 720 -2230 740 -2210
rect 760 -2230 780 -2210
rect 800 -2230 820 -2210
rect 840 -2230 860 -2210
rect 880 -2230 900 -2210
rect 920 -2230 940 -2210
rect 960 -2230 980 -2210
rect 1000 -2230 1020 -2210
rect 1040 -2230 1060 -2210
rect 1080 -2230 1100 -2210
rect 1120 -2230 1140 -2210
rect 1160 -2230 1180 -2210
rect 1200 -2230 1220 -2210
rect 1240 -2230 1260 -2210
rect 1280 -2230 1300 -2210
rect 1320 -2230 1340 -2210
rect 1360 -2230 1380 -2210
rect 1400 -2230 1420 -2210
rect 1440 -2230 1460 -2210
rect 1480 -2230 1500 -2210
rect 1520 -2230 1540 -2210
rect 1560 -2230 1580 -2210
rect 1600 -2230 1620 -2210
rect 1640 -2230 1660 -2210
rect 1680 -2230 1700 -2210
rect 1720 -2230 1740 -2210
rect 1760 -2230 1780 -2210
rect 1800 -2230 1820 -2210
rect 1840 -2230 1860 -2210
rect 1880 -2230 1900 -2210
rect 1920 -2230 1940 -2210
rect 1960 -2230 1980 -2210
rect 2000 -2230 2020 -2210
rect 2040 -2230 2060 -2210
rect 2080 -2230 2100 -2210
rect 2120 -2230 2140 -2210
rect 2160 -2230 2180 -2210
rect 2200 -2230 2220 -2210
rect 2240 -2230 2260 -2210
rect 2280 -2230 2300 -2210
rect 2320 -2230 2340 -2210
rect 2360 -2230 2380 -2210
rect 2400 -2230 2420 -2210
rect 2440 -2230 2460 -2210
rect 2480 -2230 2500 -2210
rect 2520 -2230 2540 -2210
rect 2560 -2230 2590 -2210
rect 120 -2325 140 -2305
rect 160 -2325 180 -2305
rect 200 -2325 220 -2305
rect 240 -2325 260 -2305
rect 280 -2325 300 -2305
rect 320 -2325 340 -2305
rect 360 -2325 380 -2305
rect 400 -2325 420 -2305
rect 440 -2325 460 -2305
rect 480 -2325 500 -2305
rect 520 -2325 540 -2305
rect 560 -2325 580 -2305
rect 600 -2325 620 -2305
rect 640 -2325 660 -2305
rect 680 -2325 700 -2305
rect 720 -2325 740 -2305
rect 760 -2325 780 -2305
rect 800 -2325 820 -2305
rect 840 -2325 860 -2305
rect 880 -2325 900 -2305
rect 920 -2325 940 -2305
rect 960 -2325 980 -2305
rect 1000 -2325 1020 -2305
rect 1040 -2325 1060 -2305
rect 1080 -2325 1100 -2305
rect 1120 -2325 1140 -2305
rect 1160 -2325 1180 -2305
rect 1200 -2325 1220 -2305
rect 1240 -2325 1260 -2305
rect 1280 -2325 1300 -2305
rect 1320 -2325 1340 -2305
rect 1360 -2325 1380 -2305
rect 1400 -2325 1420 -2305
rect 1440 -2325 1460 -2305
rect 1480 -2325 1500 -2305
rect 1520 -2325 1540 -2305
rect 1560 -2325 1580 -2305
rect 1600 -2325 1620 -2305
rect 1640 -2325 1660 -2305
rect 1680 -2325 1700 -2305
rect 1720 -2325 1740 -2305
rect 1760 -2325 1780 -2305
rect 1800 -2325 1820 -2305
rect 1840 -2325 1860 -2305
rect 1880 -2325 1900 -2305
rect 1920 -2325 1940 -2305
rect 1960 -2325 1980 -2305
rect 2000 -2325 2020 -2305
rect 2040 -2325 2060 -2305
rect 2080 -2325 2100 -2305
rect 2120 -2325 2140 -2305
rect 2160 -2325 2180 -2305
rect 2200 -2325 2220 -2305
rect 2240 -2325 2260 -2305
rect 2280 -2325 2300 -2305
rect 2320 -2325 2340 -2305
rect 2360 -2325 2380 -2305
rect 2400 -2325 2420 -2305
rect 2440 -2325 2460 -2305
rect 2480 -2325 2500 -2305
rect 2520 -2325 2540 -2305
rect 2560 -2325 2590 -2305
rect 120 -2420 140 -2400
rect 160 -2420 180 -2400
rect 200 -2420 220 -2400
rect 240 -2420 260 -2400
rect 280 -2420 300 -2400
rect 320 -2420 340 -2400
rect 360 -2420 380 -2400
rect 400 -2420 420 -2400
rect 440 -2420 460 -2400
rect 480 -2420 500 -2400
rect 520 -2420 540 -2400
rect 560 -2420 580 -2400
rect 600 -2420 620 -2400
rect 640 -2420 660 -2400
rect 680 -2420 700 -2400
rect 720 -2420 740 -2400
rect 760 -2420 780 -2400
rect 800 -2420 820 -2400
rect 840 -2420 860 -2400
rect 880 -2420 900 -2400
rect 920 -2420 940 -2400
rect 960 -2420 980 -2400
rect 1000 -2420 1020 -2400
rect 1040 -2420 1060 -2400
rect 1080 -2420 1100 -2400
rect 1120 -2420 1140 -2400
rect 1160 -2420 1180 -2400
rect 1200 -2420 1220 -2400
rect 1240 -2420 1260 -2400
rect 1280 -2420 1300 -2400
rect 1320 -2420 1340 -2400
rect 1360 -2420 1380 -2400
rect 1400 -2420 1420 -2400
rect 1440 -2420 1460 -2400
rect 1480 -2420 1500 -2400
rect 1520 -2420 1540 -2400
rect 1560 -2420 1580 -2400
rect 1600 -2420 1620 -2400
rect 1640 -2420 1660 -2400
rect 1680 -2420 1700 -2400
rect 1720 -2420 1740 -2400
rect 1760 -2420 1780 -2400
rect 1800 -2420 1820 -2400
rect 1840 -2420 1860 -2400
rect 1880 -2420 1900 -2400
rect 1920 -2420 1940 -2400
rect 1960 -2420 1980 -2400
rect 2000 -2420 2020 -2400
rect 2040 -2420 2060 -2400
rect 2080 -2420 2100 -2400
rect 2120 -2420 2140 -2400
rect 2160 -2420 2180 -2400
rect 2200 -2420 2220 -2400
rect 2240 -2420 2260 -2400
rect 2280 -2420 2300 -2400
rect 2320 -2420 2340 -2400
rect 2360 -2420 2380 -2400
rect 2400 -2420 2420 -2400
rect 2440 -2420 2460 -2400
rect 2480 -2420 2500 -2400
rect 2520 -2420 2540 -2400
rect 2560 -2420 2590 -2400
rect 120 -2515 140 -2495
rect 160 -2515 180 -2495
rect 200 -2515 220 -2495
rect 240 -2515 260 -2495
rect 280 -2515 300 -2495
rect 320 -2515 340 -2495
rect 360 -2515 380 -2495
rect 400 -2515 420 -2495
rect 440 -2515 460 -2495
rect 480 -2515 500 -2495
rect 520 -2515 540 -2495
rect 560 -2515 580 -2495
rect 600 -2515 620 -2495
rect 640 -2515 660 -2495
rect 680 -2515 700 -2495
rect 720 -2515 740 -2495
rect 760 -2515 780 -2495
rect 800 -2515 820 -2495
rect 840 -2515 860 -2495
rect 880 -2515 900 -2495
rect 920 -2515 940 -2495
rect 960 -2515 980 -2495
rect 1000 -2515 1020 -2495
rect 1040 -2515 1060 -2495
rect 1080 -2515 1100 -2495
rect 1120 -2515 1140 -2495
rect 1160 -2515 1180 -2495
rect 1200 -2515 1220 -2495
rect 1240 -2515 1260 -2495
rect 1280 -2515 1300 -2495
rect 1320 -2515 1340 -2495
rect 1360 -2515 1380 -2495
rect 1400 -2515 1420 -2495
rect 1440 -2515 1460 -2495
rect 1480 -2515 1500 -2495
rect 1520 -2515 1540 -2495
rect 1560 -2515 1580 -2495
rect 1600 -2515 1620 -2495
rect 1640 -2515 1660 -2495
rect 1680 -2515 1700 -2495
rect 1720 -2515 1740 -2495
rect 1760 -2515 1780 -2495
rect 1800 -2515 1820 -2495
rect 1840 -2515 1860 -2495
rect 1880 -2515 1900 -2495
rect 1920 -2515 1940 -2495
rect 1960 -2515 1980 -2495
rect 2000 -2515 2020 -2495
rect 2040 -2515 2060 -2495
rect 2080 -2515 2100 -2495
rect 2120 -2515 2140 -2495
rect 2160 -2515 2180 -2495
rect 2200 -2515 2220 -2495
rect 2240 -2515 2260 -2495
rect 2280 -2515 2300 -2495
rect 2320 -2515 2340 -2495
rect 2360 -2515 2380 -2495
rect 2400 -2515 2420 -2495
rect 2440 -2515 2460 -2495
rect 2480 -2515 2500 -2495
rect 2520 -2515 2540 -2495
rect 2560 -2515 2590 -2495
rect 120 -2610 140 -2590
rect 160 -2610 180 -2590
rect 200 -2610 220 -2590
rect 240 -2610 260 -2590
rect 280 -2610 300 -2590
rect 320 -2610 340 -2590
rect 360 -2610 380 -2590
rect 400 -2610 420 -2590
rect 440 -2610 460 -2590
rect 480 -2610 500 -2590
rect 520 -2610 540 -2590
rect 560 -2610 580 -2590
rect 600 -2610 620 -2590
rect 640 -2610 660 -2590
rect 680 -2610 700 -2590
rect 720 -2610 740 -2590
rect 760 -2610 780 -2590
rect 800 -2610 820 -2590
rect 840 -2610 860 -2590
rect 880 -2610 900 -2590
rect 920 -2610 940 -2590
rect 960 -2610 980 -2590
rect 1000 -2610 1020 -2590
rect 1040 -2610 1060 -2590
rect 1080 -2610 1100 -2590
rect 1120 -2610 1140 -2590
rect 1160 -2610 1180 -2590
rect 1200 -2610 1220 -2590
rect 1240 -2610 1260 -2590
rect 1280 -2610 1300 -2590
rect 1320 -2610 1340 -2590
rect 1360 -2610 1380 -2590
rect 1400 -2610 1420 -2590
rect 1440 -2610 1460 -2590
rect 1480 -2610 1500 -2590
rect 1520 -2610 1540 -2590
rect 1560 -2610 1580 -2590
rect 1600 -2610 1620 -2590
rect 1640 -2610 1660 -2590
rect 1680 -2610 1700 -2590
rect 1720 -2610 1740 -2590
rect 1760 -2610 1780 -2590
rect 1800 -2610 1820 -2590
rect 1840 -2610 1860 -2590
rect 1880 -2610 1900 -2590
rect 1920 -2610 1940 -2590
rect 1960 -2610 1980 -2590
rect 2000 -2610 2020 -2590
rect 2040 -2610 2060 -2590
rect 2080 -2610 2100 -2590
rect 2120 -2610 2140 -2590
rect 2160 -2610 2180 -2590
rect 2200 -2610 2220 -2590
rect 2240 -2610 2260 -2590
rect 2280 -2610 2300 -2590
rect 2320 -2610 2340 -2590
rect 2360 -2610 2380 -2590
rect 2400 -2610 2420 -2590
rect 2440 -2610 2460 -2590
rect 2480 -2610 2500 -2590
rect 2520 -2610 2540 -2590
rect 2560 -2610 2590 -2590
rect 120 -2705 140 -2685
rect 160 -2705 180 -2685
rect 200 -2705 220 -2685
rect 240 -2705 260 -2685
rect 280 -2705 300 -2685
rect 320 -2705 340 -2685
rect 360 -2705 380 -2685
rect 400 -2705 420 -2685
rect 440 -2705 460 -2685
rect 480 -2705 500 -2685
rect 520 -2705 540 -2685
rect 560 -2705 580 -2685
rect 600 -2705 620 -2685
rect 640 -2705 660 -2685
rect 680 -2705 700 -2685
rect 720 -2705 740 -2685
rect 760 -2705 780 -2685
rect 800 -2705 820 -2685
rect 840 -2705 860 -2685
rect 880 -2705 900 -2685
rect 920 -2705 940 -2685
rect 960 -2705 980 -2685
rect 1000 -2705 1020 -2685
rect 1040 -2705 1060 -2685
rect 1080 -2705 1100 -2685
rect 1120 -2705 1140 -2685
rect 1160 -2705 1180 -2685
rect 1200 -2705 1220 -2685
rect 1240 -2705 1260 -2685
rect 1280 -2705 1300 -2685
rect 1320 -2705 1340 -2685
rect 1360 -2705 1380 -2685
rect 1400 -2705 1420 -2685
rect 1440 -2705 1460 -2685
rect 1480 -2705 1500 -2685
rect 1520 -2705 1540 -2685
rect 1560 -2705 1580 -2685
rect 1600 -2705 1620 -2685
rect 1640 -2705 1660 -2685
rect 1680 -2705 1700 -2685
rect 1720 -2705 1740 -2685
rect 1760 -2705 1780 -2685
rect 1800 -2705 1820 -2685
rect 1840 -2705 1860 -2685
rect 1880 -2705 1900 -2685
rect 1920 -2705 1940 -2685
rect 1960 -2705 1980 -2685
rect 2000 -2705 2020 -2685
rect 2040 -2705 2060 -2685
rect 2080 -2705 2100 -2685
rect 2120 -2705 2140 -2685
rect 2160 -2705 2180 -2685
rect 2200 -2705 2220 -2685
rect 2240 -2705 2260 -2685
rect 2280 -2705 2300 -2685
rect 2320 -2705 2340 -2685
rect 2360 -2705 2380 -2685
rect 2400 -2705 2420 -2685
rect 2440 -2705 2460 -2685
rect 2480 -2705 2500 -2685
rect 2520 -2705 2540 -2685
rect 2560 -2705 2590 -2685
<< psubdiff >>
rect 175 2260 2675 2270
rect 175 2240 200 2260
rect 220 2240 240 2260
rect 260 2240 280 2260
rect 300 2240 320 2260
rect 340 2240 360 2260
rect 380 2240 400 2260
rect 420 2240 440 2260
rect 460 2240 480 2260
rect 500 2240 520 2260
rect 540 2240 560 2260
rect 580 2240 600 2260
rect 620 2240 640 2260
rect 660 2240 680 2260
rect 700 2240 720 2260
rect 740 2240 760 2260
rect 780 2240 800 2260
rect 820 2240 840 2260
rect 860 2240 880 2260
rect 900 2240 920 2260
rect 940 2240 960 2260
rect 980 2240 1000 2260
rect 1020 2240 1040 2260
rect 1060 2240 1080 2260
rect 1100 2240 1120 2260
rect 1140 2240 1160 2260
rect 1180 2240 1200 2260
rect 1220 2240 1240 2260
rect 1260 2240 1280 2260
rect 1300 2240 1320 2260
rect 1340 2240 1360 2260
rect 1380 2240 1400 2260
rect 1420 2240 1440 2260
rect 1460 2240 1480 2260
rect 1500 2240 1520 2260
rect 1540 2240 1560 2260
rect 1580 2240 1600 2260
rect 1620 2240 1640 2260
rect 1660 2240 1680 2260
rect 1700 2240 1720 2260
rect 1740 2240 1760 2260
rect 1780 2240 1800 2260
rect 1820 2240 1840 2260
rect 1860 2240 1880 2260
rect 1900 2240 1920 2260
rect 1940 2240 1960 2260
rect 1980 2240 2000 2260
rect 2020 2240 2040 2260
rect 2060 2240 2080 2260
rect 2100 2240 2120 2260
rect 2140 2240 2160 2260
rect 2180 2240 2200 2260
rect 2220 2240 2240 2260
rect 2260 2240 2280 2260
rect 2300 2240 2320 2260
rect 2340 2240 2360 2260
rect 2380 2240 2400 2260
rect 2420 2240 2440 2260
rect 2460 2240 2480 2260
rect 2500 2240 2520 2260
rect 2540 2240 2560 2260
rect 2580 2240 2600 2260
rect 2620 2240 2640 2260
rect 2660 2240 2675 2260
rect 175 2230 2675 2240
rect 175 45 2675 55
rect 175 25 200 45
rect 220 25 240 45
rect 260 25 280 45
rect 300 25 320 45
rect 340 25 360 45
rect 380 25 400 45
rect 420 25 440 45
rect 460 25 480 45
rect 500 25 520 45
rect 540 25 560 45
rect 580 25 600 45
rect 620 25 640 45
rect 660 25 680 45
rect 700 25 720 45
rect 740 25 760 45
rect 780 25 800 45
rect 820 25 840 45
rect 860 25 880 45
rect 900 25 920 45
rect 940 25 960 45
rect 980 25 1000 45
rect 1020 25 1040 45
rect 1060 25 1080 45
rect 1100 25 1120 45
rect 1140 25 1160 45
rect 1180 25 1200 45
rect 1220 25 1240 45
rect 1260 25 1280 45
rect 1300 25 1320 45
rect 1340 25 1360 45
rect 1380 25 1400 45
rect 1420 25 1440 45
rect 1460 25 1480 45
rect 1500 25 1520 45
rect 1540 25 1560 45
rect 1580 25 1600 45
rect 1620 25 1640 45
rect 1660 25 1680 45
rect 1700 25 1720 45
rect 1740 25 1760 45
rect 1780 25 1800 45
rect 1820 25 1840 45
rect 1860 25 1880 45
rect 1900 25 1920 45
rect 1940 25 1960 45
rect 1980 25 2000 45
rect 2020 25 2040 45
rect 2060 25 2080 45
rect 2100 25 2120 45
rect 2140 25 2160 45
rect 2180 25 2200 45
rect 2220 25 2240 45
rect 2260 25 2280 45
rect 2300 25 2320 45
rect 2340 25 2360 45
rect 2380 25 2400 45
rect 2420 25 2440 45
rect 2460 25 2480 45
rect 2500 25 2520 45
rect 2540 25 2560 45
rect 2580 25 2600 45
rect 2620 25 2640 45
rect 2660 25 2675 45
rect 175 15 2675 25
rect 105 -175 2605 -165
rect 105 -195 120 -175
rect 140 -195 160 -175
rect 180 -195 200 -175
rect 220 -195 240 -175
rect 260 -195 280 -175
rect 300 -195 320 -175
rect 340 -195 360 -175
rect 380 -195 400 -175
rect 420 -195 440 -175
rect 460 -195 480 -175
rect 500 -195 520 -175
rect 540 -195 560 -175
rect 580 -195 600 -175
rect 620 -195 640 -175
rect 660 -195 680 -175
rect 700 -195 720 -175
rect 740 -195 760 -175
rect 780 -195 800 -175
rect 820 -195 840 -175
rect 860 -195 880 -175
rect 900 -195 920 -175
rect 940 -195 960 -175
rect 980 -195 1000 -175
rect 1020 -195 1040 -175
rect 1060 -195 1080 -175
rect 1100 -195 1120 -175
rect 1140 -195 1160 -175
rect 1180 -195 1200 -175
rect 1220 -195 1240 -175
rect 1260 -195 1280 -175
rect 1300 -195 1320 -175
rect 1340 -195 1360 -175
rect 1380 -195 1400 -175
rect 1420 -195 1440 -175
rect 1460 -195 1480 -175
rect 1500 -195 1520 -175
rect 1540 -195 1560 -175
rect 1580 -195 1600 -175
rect 1620 -195 1640 -175
rect 1660 -195 1680 -175
rect 1700 -195 1720 -175
rect 1740 -195 1760 -175
rect 1780 -195 1800 -175
rect 1820 -195 1840 -175
rect 1860 -195 1880 -175
rect 1900 -195 1920 -175
rect 1940 -195 1960 -175
rect 1980 -195 2000 -175
rect 2020 -195 2040 -175
rect 2060 -195 2080 -175
rect 2100 -195 2120 -175
rect 2140 -195 2160 -175
rect 2180 -195 2200 -175
rect 2220 -195 2240 -175
rect 2260 -195 2280 -175
rect 2300 -195 2320 -175
rect 2340 -195 2360 -175
rect 2380 -195 2400 -175
rect 2420 -195 2440 -175
rect 2460 -195 2480 -175
rect 2500 -195 2520 -175
rect 2540 -195 2560 -175
rect 2590 -195 2605 -175
rect 105 -205 2605 -195
rect 105 -2725 2605 -2715
rect 105 -2745 120 -2725
rect 140 -2745 160 -2725
rect 180 -2745 200 -2725
rect 220 -2745 240 -2725
rect 260 -2745 280 -2725
rect 300 -2745 320 -2725
rect 340 -2745 360 -2725
rect 380 -2745 400 -2725
rect 420 -2745 440 -2725
rect 460 -2745 480 -2725
rect 500 -2745 520 -2725
rect 540 -2745 560 -2725
rect 580 -2745 600 -2725
rect 620 -2745 640 -2725
rect 660 -2745 680 -2725
rect 700 -2745 720 -2725
rect 740 -2745 760 -2725
rect 780 -2745 800 -2725
rect 820 -2745 840 -2725
rect 860 -2745 880 -2725
rect 900 -2745 920 -2725
rect 940 -2745 960 -2725
rect 980 -2745 1000 -2725
rect 1020 -2745 1040 -2725
rect 1060 -2745 1080 -2725
rect 1100 -2745 1120 -2725
rect 1140 -2745 1160 -2725
rect 1180 -2745 1200 -2725
rect 1220 -2745 1240 -2725
rect 1260 -2745 1280 -2725
rect 1300 -2745 1320 -2725
rect 1340 -2745 1360 -2725
rect 1380 -2745 1400 -2725
rect 1420 -2745 1440 -2725
rect 1460 -2745 1480 -2725
rect 1500 -2745 1520 -2725
rect 1540 -2745 1560 -2725
rect 1580 -2745 1600 -2725
rect 1620 -2745 1640 -2725
rect 1660 -2745 1680 -2725
rect 1700 -2745 1720 -2725
rect 1740 -2745 1760 -2725
rect 1780 -2745 1800 -2725
rect 1820 -2745 1840 -2725
rect 1860 -2745 1880 -2725
rect 1900 -2745 1920 -2725
rect 1940 -2745 1960 -2725
rect 1980 -2745 2000 -2725
rect 2020 -2745 2040 -2725
rect 2060 -2745 2080 -2725
rect 2100 -2745 2120 -2725
rect 2140 -2745 2160 -2725
rect 2180 -2745 2200 -2725
rect 2220 -2745 2240 -2725
rect 2260 -2745 2280 -2725
rect 2300 -2745 2320 -2725
rect 2340 -2745 2360 -2725
rect 2380 -2745 2400 -2725
rect 2420 -2745 2440 -2725
rect 2460 -2745 2480 -2725
rect 2500 -2745 2520 -2725
rect 2540 -2745 2560 -2725
rect 2590 -2745 2605 -2725
rect 105 -2755 2605 -2745
<< nsubdiff >>
rect -75 2345 2785 2360
rect -75 2325 -20 2345
rect 0 2325 20 2345
rect 40 2325 60 2345
rect 80 2325 100 2345
rect 120 2325 140 2345
rect 160 2325 180 2345
rect 200 2325 220 2345
rect 240 2325 260 2345
rect 280 2325 300 2345
rect 320 2325 340 2345
rect 360 2325 380 2345
rect 400 2325 420 2345
rect 440 2325 460 2345
rect 480 2325 500 2345
rect 520 2325 540 2345
rect 560 2325 580 2345
rect 600 2325 620 2345
rect 640 2325 660 2345
rect 680 2325 700 2345
rect 720 2325 740 2345
rect 760 2325 780 2345
rect 800 2325 820 2345
rect 840 2325 860 2345
rect 880 2325 900 2345
rect 920 2325 940 2345
rect 960 2325 980 2345
rect 1000 2325 1020 2345
rect 1040 2325 1060 2345
rect 1080 2325 1100 2345
rect 1120 2325 1140 2345
rect 1160 2325 1180 2345
rect 1200 2325 1220 2345
rect 1240 2325 1260 2345
rect 1280 2325 1300 2345
rect 1320 2325 1340 2345
rect 1360 2325 1380 2345
rect 1400 2325 1420 2345
rect 1440 2325 1460 2345
rect 1480 2325 1500 2345
rect 1520 2325 1540 2345
rect 1560 2325 1580 2345
rect 1600 2325 1620 2345
rect 1640 2325 1660 2345
rect 1680 2325 1700 2345
rect 1720 2325 1740 2345
rect 1760 2325 1780 2345
rect 1800 2325 1820 2345
rect 1840 2325 1860 2345
rect 1880 2325 1900 2345
rect 1920 2325 1940 2345
rect 1960 2325 1980 2345
rect 2000 2325 2020 2345
rect 2040 2325 2060 2345
rect 2080 2325 2100 2345
rect 2120 2325 2140 2345
rect 2160 2325 2180 2345
rect 2200 2325 2220 2345
rect 2240 2325 2260 2345
rect 2280 2325 2300 2345
rect 2320 2325 2340 2345
rect 2360 2325 2380 2345
rect 2400 2325 2420 2345
rect 2440 2325 2460 2345
rect 2480 2325 2500 2345
rect 2520 2325 2540 2345
rect 2560 2325 2580 2345
rect 2600 2325 2620 2345
rect 2640 2325 2660 2345
rect 2680 2325 2700 2345
rect 2720 2325 2785 2345
rect -75 2310 2785 2325
rect -75 2290 -60 2310
rect -40 2290 -25 2310
rect -75 2270 -25 2290
rect 2735 2290 2750 2310
rect 2770 2290 2785 2310
rect 2735 2270 2785 2290
rect -75 2250 -60 2270
rect -40 2250 -25 2270
rect -75 2230 -25 2250
rect -75 2210 -60 2230
rect -40 2210 -25 2230
rect -75 2190 -25 2210
rect -75 2170 -60 2190
rect -40 2170 -25 2190
rect -75 2150 -25 2170
rect -75 2130 -60 2150
rect -40 2130 -25 2150
rect 2735 2250 2750 2270
rect 2770 2250 2785 2270
rect 2735 2230 2785 2250
rect 2735 2210 2750 2230
rect 2770 2210 2785 2230
rect 2735 2190 2785 2210
rect 2735 2170 2750 2190
rect 2770 2170 2785 2190
rect 2735 2150 2785 2170
rect -75 2110 -25 2130
rect -75 2090 -60 2110
rect -40 2090 -25 2110
rect -75 2070 -25 2090
rect -75 2050 -60 2070
rect -40 2050 -25 2070
rect 2735 2130 2750 2150
rect 2770 2130 2785 2150
rect 2735 2110 2785 2130
rect 2735 2090 2750 2110
rect 2770 2090 2785 2110
rect 2735 2070 2785 2090
rect -75 2030 -25 2050
rect -75 2010 -60 2030
rect -40 2010 -25 2030
rect -75 1990 -25 2010
rect -75 1970 -60 1990
rect -40 1970 -25 1990
rect 2735 2050 2750 2070
rect 2770 2050 2785 2070
rect 2735 2030 2785 2050
rect 2735 2010 2750 2030
rect 2770 2010 2785 2030
rect 2735 1990 2785 2010
rect -75 1950 -25 1970
rect -75 1930 -60 1950
rect -40 1930 -25 1950
rect -75 1910 -25 1930
rect -75 1890 -60 1910
rect -40 1890 -25 1910
rect 2735 1970 2750 1990
rect 2770 1970 2785 1990
rect 2735 1950 2785 1970
rect 2735 1930 2750 1950
rect 2770 1930 2785 1950
rect 2735 1910 2785 1930
rect -75 1870 -25 1890
rect -75 1850 -60 1870
rect -40 1850 -25 1870
rect -75 1830 -25 1850
rect -75 1810 -60 1830
rect -40 1810 -25 1830
rect 2735 1890 2750 1910
rect 2770 1890 2785 1910
rect 2735 1870 2785 1890
rect 2735 1850 2750 1870
rect 2770 1850 2785 1870
rect 2735 1830 2785 1850
rect -75 1790 -25 1810
rect -75 1770 -60 1790
rect -40 1770 -25 1790
rect -75 1750 -25 1770
rect -75 1730 -60 1750
rect -40 1730 -25 1750
rect 2735 1810 2750 1830
rect 2770 1810 2785 1830
rect 2735 1790 2785 1810
rect 2735 1770 2750 1790
rect 2770 1770 2785 1790
rect 2735 1750 2785 1770
rect -75 1710 -25 1730
rect -75 1690 -60 1710
rect -40 1690 -25 1710
rect -75 1670 -25 1690
rect -75 1650 -60 1670
rect -40 1650 -25 1670
rect 2735 1730 2750 1750
rect 2770 1730 2785 1750
rect 2735 1710 2785 1730
rect 2735 1690 2750 1710
rect 2770 1690 2785 1710
rect 2735 1670 2785 1690
rect -75 1630 -25 1650
rect -75 1610 -60 1630
rect -40 1610 -25 1630
rect -75 1590 -25 1610
rect -75 1570 -60 1590
rect -40 1570 -25 1590
rect 2735 1650 2750 1670
rect 2770 1650 2785 1670
rect 2735 1630 2785 1650
rect 2735 1610 2750 1630
rect 2770 1610 2785 1630
rect 2735 1590 2785 1610
rect -75 1550 -25 1570
rect -75 1530 -60 1550
rect -40 1530 -25 1550
rect -75 1510 -25 1530
rect -75 1490 -60 1510
rect -40 1490 -25 1510
rect 2735 1570 2750 1590
rect 2770 1570 2785 1590
rect 2735 1550 2785 1570
rect 2735 1530 2750 1550
rect 2770 1530 2785 1550
rect 2735 1510 2785 1530
rect -75 1470 -25 1490
rect -75 1450 -60 1470
rect -40 1450 -25 1470
rect -75 1430 -25 1450
rect -75 1410 -60 1430
rect -40 1410 -25 1430
rect 2735 1490 2750 1510
rect 2770 1490 2785 1510
rect 2735 1470 2785 1490
rect 2735 1450 2750 1470
rect 2770 1450 2785 1470
rect 2735 1430 2785 1450
rect -75 1390 -25 1410
rect -75 1370 -60 1390
rect -40 1370 -25 1390
rect -75 1350 -25 1370
rect -75 1330 -60 1350
rect -40 1330 -25 1350
rect -75 1310 -25 1330
rect 2735 1410 2750 1430
rect 2770 1410 2785 1430
rect 2735 1390 2785 1410
rect 2735 1370 2750 1390
rect 2770 1370 2785 1390
rect 2735 1350 2785 1370
rect 2735 1330 2750 1350
rect 2770 1330 2785 1350
rect -75 1290 -60 1310
rect -40 1290 -25 1310
rect -75 1270 -25 1290
rect -75 1250 -60 1270
rect -40 1250 -25 1270
rect -75 1230 -25 1250
rect 2735 1310 2785 1330
rect 2735 1290 2750 1310
rect 2770 1290 2785 1310
rect 2735 1270 2785 1290
rect 2735 1250 2750 1270
rect 2770 1250 2785 1270
rect -75 1210 -60 1230
rect -40 1210 -25 1230
rect -75 1190 -25 1210
rect -75 1170 -60 1190
rect -40 1170 -25 1190
rect -75 1150 -25 1170
rect 2735 1230 2785 1250
rect 2735 1210 2750 1230
rect 2770 1210 2785 1230
rect 2735 1190 2785 1210
rect 2735 1170 2750 1190
rect 2770 1170 2785 1190
rect -75 1130 -60 1150
rect -40 1130 -25 1150
rect -75 1110 -25 1130
rect -75 1090 -60 1110
rect -40 1090 -25 1110
rect -75 1070 -25 1090
rect 2735 1150 2785 1170
rect 2735 1130 2750 1150
rect 2770 1130 2785 1150
rect 2735 1110 2785 1130
rect 2735 1090 2750 1110
rect 2770 1090 2785 1110
rect -75 1050 -60 1070
rect -40 1050 -25 1070
rect -75 1030 -25 1050
rect -75 1010 -60 1030
rect -40 1010 -25 1030
rect -75 990 -25 1010
rect 2735 1070 2785 1090
rect 2735 1050 2750 1070
rect 2770 1050 2785 1070
rect 2735 1030 2785 1050
rect 2735 1010 2750 1030
rect 2770 1010 2785 1030
rect -75 970 -60 990
rect -40 970 -25 990
rect -75 950 -25 970
rect -75 930 -60 950
rect -40 930 -25 950
rect -75 910 -25 930
rect 2735 990 2785 1010
rect 2735 970 2750 990
rect 2770 970 2785 990
rect 2735 950 2785 970
rect 2735 930 2750 950
rect 2770 930 2785 950
rect -75 890 -60 910
rect -40 890 -25 910
rect -75 870 -25 890
rect -75 850 -60 870
rect -40 850 -25 870
rect -75 830 -25 850
rect 2735 910 2785 930
rect 2735 890 2750 910
rect 2770 890 2785 910
rect 2735 870 2785 890
rect 2735 850 2750 870
rect 2770 850 2785 870
rect -75 810 -60 830
rect -40 810 -25 830
rect -75 790 -25 810
rect -75 770 -60 790
rect -40 770 -25 790
rect -75 750 -25 770
rect 2735 830 2785 850
rect 2735 810 2750 830
rect 2770 810 2785 830
rect 2735 790 2785 810
rect 2735 770 2750 790
rect 2770 770 2785 790
rect -75 730 -60 750
rect -40 730 -25 750
rect -75 710 -25 730
rect -75 690 -60 710
rect -40 690 -25 710
rect -75 670 -25 690
rect 2735 750 2785 770
rect 2735 730 2750 750
rect 2770 730 2785 750
rect 2735 710 2785 730
rect 2735 690 2750 710
rect 2770 690 2785 710
rect -75 650 -60 670
rect -40 650 -25 670
rect -75 630 -25 650
rect -75 610 -60 630
rect -40 610 -25 630
rect -75 590 -25 610
rect 2735 670 2785 690
rect 2735 650 2750 670
rect 2770 650 2785 670
rect 2735 630 2785 650
rect 2735 610 2750 630
rect 2770 610 2785 630
rect -75 570 -60 590
rect -40 570 -25 590
rect -75 550 -25 570
rect -75 530 -60 550
rect -40 530 -25 550
rect -75 510 -25 530
rect -75 490 -60 510
rect -40 490 -25 510
rect 2735 590 2785 610
rect 2735 570 2750 590
rect 2770 570 2785 590
rect 2735 550 2785 570
rect 2735 530 2750 550
rect 2770 530 2785 550
rect 2735 510 2785 530
rect -75 470 -25 490
rect -75 450 -60 470
rect -40 450 -25 470
rect -75 430 -25 450
rect -75 410 -60 430
rect -40 410 -25 430
rect 2735 490 2750 510
rect 2770 490 2785 510
rect 2735 470 2785 490
rect 2735 450 2750 470
rect 2770 450 2785 470
rect 2735 430 2785 450
rect -75 390 -25 410
rect -75 370 -60 390
rect -40 370 -25 390
rect -75 350 -25 370
rect -75 330 -60 350
rect -40 330 -25 350
rect 2735 410 2750 430
rect 2770 410 2785 430
rect 2735 390 2785 410
rect 2735 370 2750 390
rect 2770 370 2785 390
rect 2735 350 2785 370
rect -75 310 -25 330
rect -75 290 -60 310
rect -40 290 -25 310
rect -75 270 -25 290
rect -75 250 -60 270
rect -40 250 -25 270
rect 2735 330 2750 350
rect 2770 330 2785 350
rect 2735 310 2785 330
rect 2735 290 2750 310
rect 2770 290 2785 310
rect 2735 270 2785 290
rect -75 230 -25 250
rect -75 210 -60 230
rect -40 210 -25 230
rect -75 190 -25 210
rect -75 170 -60 190
rect -40 170 -25 190
rect 2735 250 2750 270
rect 2770 250 2785 270
rect 2735 230 2785 250
rect 2735 210 2750 230
rect 2770 210 2785 230
rect 2735 190 2785 210
rect -75 150 -25 170
rect -75 130 -60 150
rect -40 130 -25 150
rect -75 110 -25 130
rect -75 90 -60 110
rect -40 90 -25 110
rect 2735 170 2750 190
rect 2770 170 2785 190
rect 2735 150 2785 170
rect 2735 130 2750 150
rect 2770 130 2785 150
rect 2735 110 2785 130
rect -75 70 -25 90
rect -75 50 -60 70
rect -40 50 -25 70
rect -75 30 -25 50
rect -75 10 -60 30
rect -40 10 -25 30
rect 2735 90 2750 110
rect 2770 90 2785 110
rect 2735 70 2785 90
rect 2735 50 2750 70
rect 2770 50 2785 70
rect 2735 30 2785 50
rect -75 -10 -25 10
rect -75 -30 -60 -10
rect -40 -25 -25 -10
rect 2735 10 2750 30
rect 2770 10 2785 30
rect 2735 -10 2785 10
rect 2735 -25 2750 -10
rect -40 -30 2750 -25
rect 2770 -30 2785 -10
rect -75 -40 2785 -30
rect -75 -60 -20 -40
rect 0 -60 20 -40
rect 40 -60 60 -40
rect 80 -60 100 -40
rect 120 -60 140 -40
rect 160 -60 180 -40
rect 200 -60 220 -40
rect 240 -60 260 -40
rect 280 -60 300 -40
rect 320 -60 340 -40
rect 360 -60 380 -40
rect 400 -60 420 -40
rect 440 -60 460 -40
rect 480 -60 500 -40
rect 520 -60 540 -40
rect 560 -60 580 -40
rect 600 -60 620 -40
rect 640 -60 660 -40
rect 680 -60 700 -40
rect 720 -60 740 -40
rect 760 -60 780 -40
rect 800 -60 820 -40
rect 840 -60 860 -40
rect 880 -60 900 -40
rect 920 -60 940 -40
rect 960 -60 980 -40
rect 1000 -60 1020 -40
rect 1040 -60 1060 -40
rect 1080 -60 1100 -40
rect 1120 -60 1140 -40
rect 1160 -60 1180 -40
rect 1200 -60 1220 -40
rect 1240 -60 1260 -40
rect 1280 -60 1300 -40
rect 1320 -60 1340 -40
rect 1360 -60 1380 -40
rect 1400 -60 1420 -40
rect 1440 -60 1460 -40
rect 1480 -60 1500 -40
rect 1520 -60 1540 -40
rect 1560 -60 1580 -40
rect 1600 -60 1620 -40
rect 1640 -60 1660 -40
rect 1680 -60 1700 -40
rect 1720 -60 1740 -40
rect 1760 -60 1780 -40
rect 1800 -60 1820 -40
rect 1840 -60 1860 -40
rect 1880 -60 1900 -40
rect 1920 -60 1940 -40
rect 1960 -60 1980 -40
rect 2000 -60 2020 -40
rect 2040 -60 2060 -40
rect 2080 -60 2100 -40
rect 2120 -60 2140 -40
rect 2160 -60 2180 -40
rect 2200 -60 2220 -40
rect 2240 -60 2260 -40
rect 2280 -60 2300 -40
rect 2320 -60 2340 -40
rect 2360 -60 2380 -40
rect 2400 -60 2420 -40
rect 2440 -60 2460 -40
rect 2480 -60 2500 -40
rect 2520 -60 2540 -40
rect 2560 -60 2580 -40
rect 2600 -60 2620 -40
rect 2640 -60 2660 -40
rect 2680 -60 2700 -40
rect 2720 -60 2785 -40
rect -75 -75 2785 -60
<< psubdiffcont >>
rect 200 2240 220 2260
rect 240 2240 260 2260
rect 280 2240 300 2260
rect 320 2240 340 2260
rect 360 2240 380 2260
rect 400 2240 420 2260
rect 440 2240 460 2260
rect 480 2240 500 2260
rect 520 2240 540 2260
rect 560 2240 580 2260
rect 600 2240 620 2260
rect 640 2240 660 2260
rect 680 2240 700 2260
rect 720 2240 740 2260
rect 760 2240 780 2260
rect 800 2240 820 2260
rect 840 2240 860 2260
rect 880 2240 900 2260
rect 920 2240 940 2260
rect 960 2240 980 2260
rect 1000 2240 1020 2260
rect 1040 2240 1060 2260
rect 1080 2240 1100 2260
rect 1120 2240 1140 2260
rect 1160 2240 1180 2260
rect 1200 2240 1220 2260
rect 1240 2240 1260 2260
rect 1280 2240 1300 2260
rect 1320 2240 1340 2260
rect 1360 2240 1380 2260
rect 1400 2240 1420 2260
rect 1440 2240 1460 2260
rect 1480 2240 1500 2260
rect 1520 2240 1540 2260
rect 1560 2240 1580 2260
rect 1600 2240 1620 2260
rect 1640 2240 1660 2260
rect 1680 2240 1700 2260
rect 1720 2240 1740 2260
rect 1760 2240 1780 2260
rect 1800 2240 1820 2260
rect 1840 2240 1860 2260
rect 1880 2240 1900 2260
rect 1920 2240 1940 2260
rect 1960 2240 1980 2260
rect 2000 2240 2020 2260
rect 2040 2240 2060 2260
rect 2080 2240 2100 2260
rect 2120 2240 2140 2260
rect 2160 2240 2180 2260
rect 2200 2240 2220 2260
rect 2240 2240 2260 2260
rect 2280 2240 2300 2260
rect 2320 2240 2340 2260
rect 2360 2240 2380 2260
rect 2400 2240 2420 2260
rect 2440 2240 2460 2260
rect 2480 2240 2500 2260
rect 2520 2240 2540 2260
rect 2560 2240 2580 2260
rect 2600 2240 2620 2260
rect 2640 2240 2660 2260
rect 200 25 220 45
rect 240 25 260 45
rect 280 25 300 45
rect 320 25 340 45
rect 360 25 380 45
rect 400 25 420 45
rect 440 25 460 45
rect 480 25 500 45
rect 520 25 540 45
rect 560 25 580 45
rect 600 25 620 45
rect 640 25 660 45
rect 680 25 700 45
rect 720 25 740 45
rect 760 25 780 45
rect 800 25 820 45
rect 840 25 860 45
rect 880 25 900 45
rect 920 25 940 45
rect 960 25 980 45
rect 1000 25 1020 45
rect 1040 25 1060 45
rect 1080 25 1100 45
rect 1120 25 1140 45
rect 1160 25 1180 45
rect 1200 25 1220 45
rect 1240 25 1260 45
rect 1280 25 1300 45
rect 1320 25 1340 45
rect 1360 25 1380 45
rect 1400 25 1420 45
rect 1440 25 1460 45
rect 1480 25 1500 45
rect 1520 25 1540 45
rect 1560 25 1580 45
rect 1600 25 1620 45
rect 1640 25 1660 45
rect 1680 25 1700 45
rect 1720 25 1740 45
rect 1760 25 1780 45
rect 1800 25 1820 45
rect 1840 25 1860 45
rect 1880 25 1900 45
rect 1920 25 1940 45
rect 1960 25 1980 45
rect 2000 25 2020 45
rect 2040 25 2060 45
rect 2080 25 2100 45
rect 2120 25 2140 45
rect 2160 25 2180 45
rect 2200 25 2220 45
rect 2240 25 2260 45
rect 2280 25 2300 45
rect 2320 25 2340 45
rect 2360 25 2380 45
rect 2400 25 2420 45
rect 2440 25 2460 45
rect 2480 25 2500 45
rect 2520 25 2540 45
rect 2560 25 2580 45
rect 2600 25 2620 45
rect 2640 25 2660 45
rect 120 -195 140 -175
rect 160 -195 180 -175
rect 200 -195 220 -175
rect 240 -195 260 -175
rect 280 -195 300 -175
rect 320 -195 340 -175
rect 360 -195 380 -175
rect 400 -195 420 -175
rect 440 -195 460 -175
rect 480 -195 500 -175
rect 520 -195 540 -175
rect 560 -195 580 -175
rect 600 -195 620 -175
rect 640 -195 660 -175
rect 680 -195 700 -175
rect 720 -195 740 -175
rect 760 -195 780 -175
rect 800 -195 820 -175
rect 840 -195 860 -175
rect 880 -195 900 -175
rect 920 -195 940 -175
rect 960 -195 980 -175
rect 1000 -195 1020 -175
rect 1040 -195 1060 -175
rect 1080 -195 1100 -175
rect 1120 -195 1140 -175
rect 1160 -195 1180 -175
rect 1200 -195 1220 -175
rect 1240 -195 1260 -175
rect 1280 -195 1300 -175
rect 1320 -195 1340 -175
rect 1360 -195 1380 -175
rect 1400 -195 1420 -175
rect 1440 -195 1460 -175
rect 1480 -195 1500 -175
rect 1520 -195 1540 -175
rect 1560 -195 1580 -175
rect 1600 -195 1620 -175
rect 1640 -195 1660 -175
rect 1680 -195 1700 -175
rect 1720 -195 1740 -175
rect 1760 -195 1780 -175
rect 1800 -195 1820 -175
rect 1840 -195 1860 -175
rect 1880 -195 1900 -175
rect 1920 -195 1940 -175
rect 1960 -195 1980 -175
rect 2000 -195 2020 -175
rect 2040 -195 2060 -175
rect 2080 -195 2100 -175
rect 2120 -195 2140 -175
rect 2160 -195 2180 -175
rect 2200 -195 2220 -175
rect 2240 -195 2260 -175
rect 2280 -195 2300 -175
rect 2320 -195 2340 -175
rect 2360 -195 2380 -175
rect 2400 -195 2420 -175
rect 2440 -195 2460 -175
rect 2480 -195 2500 -175
rect 2520 -195 2540 -175
rect 2560 -195 2590 -175
rect 120 -2745 140 -2725
rect 160 -2745 180 -2725
rect 200 -2745 220 -2725
rect 240 -2745 260 -2725
rect 280 -2745 300 -2725
rect 320 -2745 340 -2725
rect 360 -2745 380 -2725
rect 400 -2745 420 -2725
rect 440 -2745 460 -2725
rect 480 -2745 500 -2725
rect 520 -2745 540 -2725
rect 560 -2745 580 -2725
rect 600 -2745 620 -2725
rect 640 -2745 660 -2725
rect 680 -2745 700 -2725
rect 720 -2745 740 -2725
rect 760 -2745 780 -2725
rect 800 -2745 820 -2725
rect 840 -2745 860 -2725
rect 880 -2745 900 -2725
rect 920 -2745 940 -2725
rect 960 -2745 980 -2725
rect 1000 -2745 1020 -2725
rect 1040 -2745 1060 -2725
rect 1080 -2745 1100 -2725
rect 1120 -2745 1140 -2725
rect 1160 -2745 1180 -2725
rect 1200 -2745 1220 -2725
rect 1240 -2745 1260 -2725
rect 1280 -2745 1300 -2725
rect 1320 -2745 1340 -2725
rect 1360 -2745 1380 -2725
rect 1400 -2745 1420 -2725
rect 1440 -2745 1460 -2725
rect 1480 -2745 1500 -2725
rect 1520 -2745 1540 -2725
rect 1560 -2745 1580 -2725
rect 1600 -2745 1620 -2725
rect 1640 -2745 1660 -2725
rect 1680 -2745 1700 -2725
rect 1720 -2745 1740 -2725
rect 1760 -2745 1780 -2725
rect 1800 -2745 1820 -2725
rect 1840 -2745 1860 -2725
rect 1880 -2745 1900 -2725
rect 1920 -2745 1940 -2725
rect 1960 -2745 1980 -2725
rect 2000 -2745 2020 -2725
rect 2040 -2745 2060 -2725
rect 2080 -2745 2100 -2725
rect 2120 -2745 2140 -2725
rect 2160 -2745 2180 -2725
rect 2200 -2745 2220 -2725
rect 2240 -2745 2260 -2725
rect 2280 -2745 2300 -2725
rect 2320 -2745 2340 -2725
rect 2360 -2745 2380 -2725
rect 2400 -2745 2420 -2725
rect 2440 -2745 2460 -2725
rect 2480 -2745 2500 -2725
rect 2520 -2745 2540 -2725
rect 2560 -2745 2590 -2725
<< nsubdiffcont >>
rect -20 2325 0 2345
rect 20 2325 40 2345
rect 60 2325 80 2345
rect 100 2325 120 2345
rect 140 2325 160 2345
rect 180 2325 200 2345
rect 220 2325 240 2345
rect 260 2325 280 2345
rect 300 2325 320 2345
rect 340 2325 360 2345
rect 380 2325 400 2345
rect 420 2325 440 2345
rect 460 2325 480 2345
rect 500 2325 520 2345
rect 540 2325 560 2345
rect 580 2325 600 2345
rect 620 2325 640 2345
rect 660 2325 680 2345
rect 700 2325 720 2345
rect 740 2325 760 2345
rect 780 2325 800 2345
rect 820 2325 840 2345
rect 860 2325 880 2345
rect 900 2325 920 2345
rect 940 2325 960 2345
rect 980 2325 1000 2345
rect 1020 2325 1040 2345
rect 1060 2325 1080 2345
rect 1100 2325 1120 2345
rect 1140 2325 1160 2345
rect 1180 2325 1200 2345
rect 1220 2325 1240 2345
rect 1260 2325 1280 2345
rect 1300 2325 1320 2345
rect 1340 2325 1360 2345
rect 1380 2325 1400 2345
rect 1420 2325 1440 2345
rect 1460 2325 1480 2345
rect 1500 2325 1520 2345
rect 1540 2325 1560 2345
rect 1580 2325 1600 2345
rect 1620 2325 1640 2345
rect 1660 2325 1680 2345
rect 1700 2325 1720 2345
rect 1740 2325 1760 2345
rect 1780 2325 1800 2345
rect 1820 2325 1840 2345
rect 1860 2325 1880 2345
rect 1900 2325 1920 2345
rect 1940 2325 1960 2345
rect 1980 2325 2000 2345
rect 2020 2325 2040 2345
rect 2060 2325 2080 2345
rect 2100 2325 2120 2345
rect 2140 2325 2160 2345
rect 2180 2325 2200 2345
rect 2220 2325 2240 2345
rect 2260 2325 2280 2345
rect 2300 2325 2320 2345
rect 2340 2325 2360 2345
rect 2380 2325 2400 2345
rect 2420 2325 2440 2345
rect 2460 2325 2480 2345
rect 2500 2325 2520 2345
rect 2540 2325 2560 2345
rect 2580 2325 2600 2345
rect 2620 2325 2640 2345
rect 2660 2325 2680 2345
rect 2700 2325 2720 2345
rect -60 2290 -40 2310
rect 2750 2290 2770 2310
rect -60 2250 -40 2270
rect -60 2210 -40 2230
rect -60 2170 -40 2190
rect -60 2130 -40 2150
rect 2750 2250 2770 2270
rect 2750 2210 2770 2230
rect 2750 2170 2770 2190
rect -60 2090 -40 2110
rect -60 2050 -40 2070
rect 2750 2130 2770 2150
rect 2750 2090 2770 2110
rect -60 2010 -40 2030
rect -60 1970 -40 1990
rect 2750 2050 2770 2070
rect 2750 2010 2770 2030
rect -60 1930 -40 1950
rect -60 1890 -40 1910
rect 2750 1970 2770 1990
rect 2750 1930 2770 1950
rect -60 1850 -40 1870
rect -60 1810 -40 1830
rect 2750 1890 2770 1910
rect 2750 1850 2770 1870
rect -60 1770 -40 1790
rect -60 1730 -40 1750
rect 2750 1810 2770 1830
rect 2750 1770 2770 1790
rect -60 1690 -40 1710
rect -60 1650 -40 1670
rect 2750 1730 2770 1750
rect 2750 1690 2770 1710
rect -60 1610 -40 1630
rect -60 1570 -40 1590
rect 2750 1650 2770 1670
rect 2750 1610 2770 1630
rect -60 1530 -40 1550
rect -60 1490 -40 1510
rect 2750 1570 2770 1590
rect 2750 1530 2770 1550
rect -60 1450 -40 1470
rect -60 1410 -40 1430
rect 2750 1490 2770 1510
rect 2750 1450 2770 1470
rect -60 1370 -40 1390
rect -60 1330 -40 1350
rect 2750 1410 2770 1430
rect 2750 1370 2770 1390
rect 2750 1330 2770 1350
rect -60 1290 -40 1310
rect -60 1250 -40 1270
rect 2750 1290 2770 1310
rect 2750 1250 2770 1270
rect -60 1210 -40 1230
rect -60 1170 -40 1190
rect 2750 1210 2770 1230
rect 2750 1170 2770 1190
rect -60 1130 -40 1150
rect -60 1090 -40 1110
rect 2750 1130 2770 1150
rect 2750 1090 2770 1110
rect -60 1050 -40 1070
rect -60 1010 -40 1030
rect 2750 1050 2770 1070
rect 2750 1010 2770 1030
rect -60 970 -40 990
rect -60 930 -40 950
rect 2750 970 2770 990
rect 2750 930 2770 950
rect -60 890 -40 910
rect -60 850 -40 870
rect 2750 890 2770 910
rect 2750 850 2770 870
rect -60 810 -40 830
rect -60 770 -40 790
rect 2750 810 2770 830
rect 2750 770 2770 790
rect -60 730 -40 750
rect -60 690 -40 710
rect 2750 730 2770 750
rect 2750 690 2770 710
rect -60 650 -40 670
rect -60 610 -40 630
rect 2750 650 2770 670
rect 2750 610 2770 630
rect -60 570 -40 590
rect -60 530 -40 550
rect -60 490 -40 510
rect 2750 570 2770 590
rect 2750 530 2770 550
rect -60 450 -40 470
rect -60 410 -40 430
rect 2750 490 2770 510
rect 2750 450 2770 470
rect -60 370 -40 390
rect -60 330 -40 350
rect 2750 410 2770 430
rect 2750 370 2770 390
rect -60 290 -40 310
rect -60 250 -40 270
rect 2750 330 2770 350
rect 2750 290 2770 310
rect -60 210 -40 230
rect -60 170 -40 190
rect 2750 250 2770 270
rect 2750 210 2770 230
rect -60 130 -40 150
rect -60 90 -40 110
rect 2750 170 2770 190
rect 2750 130 2770 150
rect -60 50 -40 70
rect -60 10 -40 30
rect 2750 90 2770 110
rect 2750 50 2770 70
rect -60 -30 -40 -10
rect 2750 10 2770 30
rect 2750 -30 2770 -10
rect -20 -60 0 -40
rect 20 -60 40 -40
rect 60 -60 80 -40
rect 100 -60 120 -40
rect 140 -60 160 -40
rect 180 -60 200 -40
rect 220 -60 240 -40
rect 260 -60 280 -40
rect 300 -60 320 -40
rect 340 -60 360 -40
rect 380 -60 400 -40
rect 420 -60 440 -40
rect 460 -60 480 -40
rect 500 -60 520 -40
rect 540 -60 560 -40
rect 580 -60 600 -40
rect 620 -60 640 -40
rect 660 -60 680 -40
rect 700 -60 720 -40
rect 740 -60 760 -40
rect 780 -60 800 -40
rect 820 -60 840 -40
rect 860 -60 880 -40
rect 900 -60 920 -40
rect 940 -60 960 -40
rect 980 -60 1000 -40
rect 1020 -60 1040 -40
rect 1060 -60 1080 -40
rect 1100 -60 1120 -40
rect 1140 -60 1160 -40
rect 1180 -60 1200 -40
rect 1220 -60 1240 -40
rect 1260 -60 1280 -40
rect 1300 -60 1320 -40
rect 1340 -60 1360 -40
rect 1380 -60 1400 -40
rect 1420 -60 1440 -40
rect 1460 -60 1480 -40
rect 1500 -60 1520 -40
rect 1540 -60 1560 -40
rect 1580 -60 1600 -40
rect 1620 -60 1640 -40
rect 1660 -60 1680 -40
rect 1700 -60 1720 -40
rect 1740 -60 1760 -40
rect 1780 -60 1800 -40
rect 1820 -60 1840 -40
rect 1860 -60 1880 -40
rect 1900 -60 1920 -40
rect 1940 -60 1960 -40
rect 1980 -60 2000 -40
rect 2020 -60 2040 -40
rect 2060 -60 2080 -40
rect 2100 -60 2120 -40
rect 2140 -60 2160 -40
rect 2180 -60 2200 -40
rect 2220 -60 2240 -40
rect 2260 -60 2280 -40
rect 2300 -60 2320 -40
rect 2340 -60 2360 -40
rect 2380 -60 2400 -40
rect 2420 -60 2440 -40
rect 2460 -60 2480 -40
rect 2500 -60 2520 -40
rect 2540 -60 2560 -40
rect 2580 -60 2600 -40
rect 2620 -60 2640 -40
rect 2660 -60 2680 -40
rect 2700 -60 2720 -40
<< poly >>
rect 0 2182 165 2185
rect 0 2175 175 2182
rect 0 2155 10 2175
rect 30 2155 50 2175
rect 70 2155 90 2175
rect 110 2155 130 2175
rect 155 2155 175 2175
rect 0 2150 175 2155
rect 2675 2150 2690 2182
rect 0 2145 165 2150
rect 0 2100 165 2105
rect 0 2095 175 2100
rect 0 2075 10 2095
rect 30 2075 50 2095
rect 70 2075 90 2095
rect 110 2075 130 2095
rect 155 2075 175 2095
rect 0 2068 175 2075
rect 2675 2068 2690 2100
rect 0 2065 165 2068
rect 0 2018 165 2020
rect 0 2010 175 2018
rect 0 1990 10 2010
rect 30 1990 50 2010
rect 70 1990 90 2010
rect 110 1990 130 2010
rect 155 1990 175 2010
rect 0 1986 175 1990
rect 2675 1986 2690 2018
rect 0 1980 165 1986
rect 0 1936 165 1940
rect 0 1930 175 1936
rect 0 1910 10 1930
rect 30 1910 50 1930
rect 70 1910 90 1930
rect 110 1910 130 1930
rect 155 1910 175 1930
rect 0 1904 175 1910
rect 2675 1904 2690 1936
rect 0 1900 165 1904
rect 0 1854 165 1860
rect 0 1850 175 1854
rect 0 1830 10 1850
rect 30 1830 50 1850
rect 70 1830 90 1850
rect 110 1830 130 1850
rect 155 1830 175 1850
rect 0 1822 175 1830
rect 2675 1822 2690 1854
rect 0 1820 165 1822
rect 0 1772 165 1775
rect 0 1765 175 1772
rect 0 1745 10 1765
rect 30 1745 50 1765
rect 70 1745 90 1765
rect 110 1745 130 1765
rect 155 1745 175 1765
rect 0 1740 175 1745
rect 2675 1740 2690 1772
rect 0 1735 165 1740
rect 0 1690 165 1695
rect 0 1685 175 1690
rect 0 1665 10 1685
rect 30 1665 50 1685
rect 70 1665 90 1685
rect 110 1665 130 1685
rect 155 1665 175 1685
rect 0 1658 175 1665
rect 2675 1658 2690 1690
rect 0 1655 165 1658
rect 0 1608 165 1610
rect 0 1600 175 1608
rect 0 1580 10 1600
rect 30 1580 50 1600
rect 70 1580 90 1600
rect 110 1580 130 1600
rect 155 1580 175 1600
rect 0 1576 175 1580
rect 2675 1576 2690 1608
rect 0 1570 165 1576
rect 0 1526 165 1530
rect 0 1520 175 1526
rect 0 1500 10 1520
rect 30 1500 50 1520
rect 70 1500 90 1520
rect 110 1500 130 1520
rect 155 1500 175 1520
rect 0 1494 175 1500
rect 2675 1494 2690 1526
rect 0 1490 165 1494
rect 0 1444 165 1450
rect 0 1440 175 1444
rect 0 1420 10 1440
rect 30 1420 50 1440
rect 70 1420 90 1440
rect 110 1420 130 1440
rect 155 1420 175 1440
rect 0 1412 175 1420
rect 2675 1412 2690 1444
rect 0 1410 165 1412
rect 0 1362 165 1365
rect 0 1355 175 1362
rect 0 1335 10 1355
rect 30 1335 50 1355
rect 70 1335 90 1355
rect 110 1335 130 1355
rect 155 1335 175 1355
rect 0 1330 175 1335
rect 2675 1330 2690 1362
rect 0 1325 165 1330
rect 0 1280 165 1285
rect 0 1275 175 1280
rect 0 1255 10 1275
rect 30 1255 50 1275
rect 70 1255 90 1275
rect 110 1255 130 1275
rect 155 1255 175 1275
rect 0 1248 175 1255
rect 2675 1248 2690 1280
rect 0 1245 165 1248
rect 0 1198 165 1200
rect 0 1190 175 1198
rect 0 1170 10 1190
rect 30 1170 50 1190
rect 70 1170 90 1190
rect 110 1170 130 1190
rect 155 1170 175 1190
rect 0 1166 175 1170
rect 2675 1166 2690 1198
rect 0 1160 165 1166
rect 0 1116 165 1120
rect 0 1110 175 1116
rect 0 1090 10 1110
rect 30 1090 50 1110
rect 70 1090 90 1110
rect 110 1090 130 1110
rect 155 1090 175 1110
rect 0 1084 175 1090
rect 2675 1084 2690 1116
rect 0 1080 165 1084
rect 0 1034 165 1040
rect 0 1030 175 1034
rect 0 1010 10 1030
rect 30 1010 50 1030
rect 70 1010 90 1030
rect 110 1010 130 1030
rect 155 1010 175 1030
rect 0 1002 175 1010
rect 2675 1002 2690 1034
rect 0 1000 165 1002
rect 0 952 165 955
rect 0 945 175 952
rect 0 925 10 945
rect 30 925 50 945
rect 70 925 90 945
rect 110 925 130 945
rect 155 925 175 945
rect 0 920 175 925
rect 2675 920 2690 952
rect 0 915 165 920
rect 0 870 165 875
rect 0 865 175 870
rect 0 845 10 865
rect 30 845 50 865
rect 70 845 90 865
rect 110 845 130 865
rect 155 845 175 865
rect 0 838 175 845
rect 2675 838 2690 870
rect 0 835 165 838
rect 0 788 165 790
rect 0 780 175 788
rect 0 760 10 780
rect 30 760 50 780
rect 70 760 90 780
rect 110 760 130 780
rect 155 760 175 780
rect 0 756 175 760
rect 2675 756 2690 788
rect 0 750 165 756
rect 0 706 165 710
rect 0 700 175 706
rect 0 680 10 700
rect 30 680 50 700
rect 70 680 90 700
rect 110 680 130 700
rect 155 680 175 700
rect 0 674 175 680
rect 2675 674 2690 706
rect 0 670 165 674
rect 0 624 165 630
rect 0 620 175 624
rect 0 600 10 620
rect 30 600 50 620
rect 70 600 90 620
rect 110 600 130 620
rect 155 600 175 620
rect 0 592 175 600
rect 2675 592 2690 624
rect 0 590 165 592
rect 0 542 165 545
rect 0 535 175 542
rect 0 515 10 535
rect 30 515 50 535
rect 70 515 90 535
rect 110 515 130 535
rect 155 515 175 535
rect 0 510 175 515
rect 2675 510 2690 542
rect 0 505 165 510
rect 0 460 165 465
rect 0 455 175 460
rect 0 435 10 455
rect 30 435 50 455
rect 70 435 90 455
rect 110 435 130 455
rect 155 435 175 455
rect 0 428 175 435
rect 2675 428 2690 460
rect 0 425 165 428
rect 0 378 165 385
rect 0 375 175 378
rect 0 355 10 375
rect 30 355 50 375
rect 70 355 90 375
rect 110 355 130 375
rect 155 355 175 375
rect 0 346 175 355
rect 2675 346 2690 378
rect 0 345 165 346
rect 0 296 165 300
rect 0 290 175 296
rect 0 270 10 290
rect 30 270 50 290
rect 70 270 90 290
rect 110 270 130 290
rect 155 270 175 290
rect 0 264 175 270
rect 2675 264 2690 296
rect 0 260 165 264
rect 0 214 165 220
rect 0 210 175 214
rect 0 190 10 210
rect 30 190 50 210
rect 70 190 90 210
rect 110 190 130 210
rect 155 190 175 210
rect 0 182 175 190
rect 2675 182 2690 214
rect 0 180 165 182
rect 0 132 165 140
rect 0 130 175 132
rect 0 110 10 130
rect 30 110 50 130
rect 70 110 90 130
rect 110 110 130 130
rect 155 110 175 130
rect 0 100 175 110
rect 2675 100 2690 132
rect -70 -260 105 -250
rect -70 -285 -60 -260
rect -40 -285 -20 -260
rect 0 -285 20 -260
rect 40 -285 60 -260
rect 85 -285 105 -260
rect -70 -295 105 -285
rect 2605 -295 2620 -250
rect -70 -355 105 -345
rect -70 -380 -60 -355
rect -40 -380 -20 -355
rect 0 -380 20 -355
rect 40 -380 60 -355
rect 85 -380 105 -355
rect -70 -390 105 -380
rect 2605 -390 2620 -345
rect -70 -450 105 -440
rect -70 -475 -60 -450
rect -40 -475 -20 -450
rect 0 -475 20 -450
rect 40 -475 60 -450
rect 85 -475 105 -450
rect -70 -485 105 -475
rect 2605 -485 2620 -440
rect -70 -545 105 -535
rect -70 -570 -60 -545
rect -40 -570 -20 -545
rect 0 -570 20 -545
rect 40 -570 60 -545
rect 85 -570 105 -545
rect -70 -580 105 -570
rect 2605 -580 2620 -535
rect -70 -640 105 -630
rect -70 -665 -60 -640
rect -40 -665 -20 -640
rect 0 -665 20 -640
rect 40 -665 60 -640
rect 85 -665 105 -640
rect -70 -675 105 -665
rect 2605 -675 2620 -630
rect -70 -735 105 -725
rect -70 -760 -60 -735
rect -40 -760 -20 -735
rect 0 -760 20 -735
rect 40 -760 60 -735
rect 85 -760 105 -735
rect -70 -770 105 -760
rect 2605 -770 2620 -725
rect -70 -830 105 -820
rect -70 -855 -60 -830
rect -40 -855 -20 -830
rect 0 -855 20 -830
rect 40 -855 60 -830
rect 85 -855 105 -830
rect -70 -865 105 -855
rect 2605 -865 2620 -820
rect -70 -925 105 -915
rect -70 -950 -60 -925
rect -40 -950 -20 -925
rect 0 -950 20 -925
rect 40 -950 60 -925
rect 85 -950 105 -925
rect -70 -960 105 -950
rect 2605 -960 2620 -915
rect -70 -1020 105 -1010
rect -70 -1045 -60 -1020
rect -40 -1045 -20 -1020
rect 0 -1045 20 -1020
rect 40 -1045 60 -1020
rect 85 -1045 105 -1020
rect -70 -1055 105 -1045
rect 2605 -1055 2620 -1010
rect -70 -1115 105 -1105
rect -70 -1140 -60 -1115
rect -40 -1140 -20 -1115
rect 0 -1140 20 -1115
rect 40 -1140 60 -1115
rect 85 -1140 105 -1115
rect -70 -1150 105 -1140
rect 2605 -1150 2620 -1105
rect -70 -1210 105 -1200
rect -70 -1235 -60 -1210
rect -40 -1235 -20 -1210
rect 0 -1235 20 -1210
rect 40 -1235 60 -1210
rect 85 -1235 105 -1210
rect -70 -1245 105 -1235
rect 2605 -1245 2620 -1200
rect -70 -1305 105 -1295
rect -70 -1330 -60 -1305
rect -40 -1330 -20 -1305
rect 0 -1330 20 -1305
rect 40 -1330 60 -1305
rect 85 -1330 105 -1305
rect -70 -1340 105 -1330
rect 2605 -1340 2620 -1295
rect -70 -1400 105 -1390
rect -70 -1425 -60 -1400
rect -40 -1425 -20 -1400
rect 0 -1425 20 -1400
rect 40 -1425 60 -1400
rect 85 -1425 105 -1400
rect -70 -1435 105 -1425
rect 2605 -1435 2620 -1390
rect -70 -1495 105 -1485
rect -70 -1520 -60 -1495
rect -40 -1520 -20 -1495
rect 0 -1520 20 -1495
rect 40 -1520 60 -1495
rect 85 -1520 105 -1495
rect -70 -1530 105 -1520
rect 2605 -1530 2620 -1485
rect -70 -1590 105 -1580
rect -70 -1615 -60 -1590
rect -40 -1615 -20 -1590
rect 0 -1615 20 -1590
rect 40 -1615 60 -1590
rect 85 -1615 105 -1590
rect -70 -1625 105 -1615
rect 2605 -1625 2620 -1580
rect -70 -1685 105 -1675
rect -70 -1710 -60 -1685
rect -40 -1710 -20 -1685
rect 0 -1710 20 -1685
rect 40 -1710 60 -1685
rect 85 -1710 105 -1685
rect -70 -1720 105 -1710
rect 2605 -1720 2620 -1675
rect -70 -1780 105 -1770
rect -70 -1805 -60 -1780
rect -40 -1805 -20 -1780
rect 0 -1805 20 -1780
rect 40 -1805 60 -1780
rect 85 -1805 105 -1780
rect -70 -1815 105 -1805
rect 2605 -1815 2620 -1770
rect -70 -1875 105 -1865
rect -70 -1900 -60 -1875
rect -40 -1900 -20 -1875
rect 0 -1900 20 -1875
rect 40 -1900 60 -1875
rect 85 -1900 105 -1875
rect -70 -1910 105 -1900
rect 2605 -1910 2620 -1865
rect -70 -1970 105 -1960
rect -70 -1995 -60 -1970
rect -40 -1995 -20 -1970
rect 0 -1995 20 -1970
rect 40 -1995 60 -1970
rect 85 -1995 105 -1970
rect -70 -2005 105 -1995
rect 2605 -2005 2620 -1960
rect -70 -2065 105 -2055
rect -70 -2090 -60 -2065
rect -40 -2090 -20 -2065
rect 0 -2090 20 -2065
rect 40 -2090 60 -2065
rect 85 -2090 105 -2065
rect -70 -2100 105 -2090
rect 2605 -2100 2620 -2055
rect -70 -2160 105 -2150
rect -70 -2185 -60 -2160
rect -40 -2185 -20 -2160
rect 0 -2185 20 -2160
rect 40 -2185 60 -2160
rect 85 -2185 105 -2160
rect -70 -2195 105 -2185
rect 2605 -2195 2620 -2150
rect -70 -2255 105 -2245
rect -70 -2280 -60 -2255
rect -40 -2280 -20 -2255
rect 0 -2280 20 -2255
rect 40 -2280 60 -2255
rect 85 -2280 105 -2255
rect -70 -2290 105 -2280
rect 2605 -2290 2620 -2245
rect -70 -2350 105 -2340
rect -70 -2375 -60 -2350
rect -40 -2375 -20 -2350
rect 0 -2375 20 -2350
rect 40 -2375 60 -2350
rect 85 -2375 105 -2350
rect -70 -2385 105 -2375
rect 2605 -2385 2620 -2340
rect -70 -2445 105 -2435
rect -70 -2470 -60 -2445
rect -40 -2470 -20 -2445
rect 0 -2470 20 -2445
rect 40 -2470 60 -2445
rect 85 -2470 105 -2445
rect -70 -2480 105 -2470
rect 2605 -2480 2620 -2435
rect -70 -2540 105 -2530
rect -70 -2565 -60 -2540
rect -40 -2565 -20 -2540
rect 0 -2565 20 -2540
rect 40 -2565 60 -2540
rect 85 -2565 105 -2540
rect -70 -2575 105 -2565
rect 2605 -2575 2620 -2530
rect -70 -2635 105 -2625
rect -70 -2660 -60 -2635
rect -40 -2660 -20 -2635
rect 0 -2660 20 -2635
rect 40 -2660 60 -2635
rect 85 -2660 105 -2635
rect -70 -2670 105 -2660
rect 2605 -2670 2620 -2625
<< polycont >>
rect 10 2155 30 2175
rect 50 2155 70 2175
rect 90 2155 110 2175
rect 130 2155 155 2175
rect 10 2075 30 2095
rect 50 2075 70 2095
rect 90 2075 110 2095
rect 130 2075 155 2095
rect 10 1990 30 2010
rect 50 1990 70 2010
rect 90 1990 110 2010
rect 130 1990 155 2010
rect 10 1910 30 1930
rect 50 1910 70 1930
rect 90 1910 110 1930
rect 130 1910 155 1930
rect 10 1830 30 1850
rect 50 1830 70 1850
rect 90 1830 110 1850
rect 130 1830 155 1850
rect 10 1745 30 1765
rect 50 1745 70 1765
rect 90 1745 110 1765
rect 130 1745 155 1765
rect 10 1665 30 1685
rect 50 1665 70 1685
rect 90 1665 110 1685
rect 130 1665 155 1685
rect 10 1580 30 1600
rect 50 1580 70 1600
rect 90 1580 110 1600
rect 130 1580 155 1600
rect 10 1500 30 1520
rect 50 1500 70 1520
rect 90 1500 110 1520
rect 130 1500 155 1520
rect 10 1420 30 1440
rect 50 1420 70 1440
rect 90 1420 110 1440
rect 130 1420 155 1440
rect 10 1335 30 1355
rect 50 1335 70 1355
rect 90 1335 110 1355
rect 130 1335 155 1355
rect 10 1255 30 1275
rect 50 1255 70 1275
rect 90 1255 110 1275
rect 130 1255 155 1275
rect 10 1170 30 1190
rect 50 1170 70 1190
rect 90 1170 110 1190
rect 130 1170 155 1190
rect 10 1090 30 1110
rect 50 1090 70 1110
rect 90 1090 110 1110
rect 130 1090 155 1110
rect 10 1010 30 1030
rect 50 1010 70 1030
rect 90 1010 110 1030
rect 130 1010 155 1030
rect 10 925 30 945
rect 50 925 70 945
rect 90 925 110 945
rect 130 925 155 945
rect 10 845 30 865
rect 50 845 70 865
rect 90 845 110 865
rect 130 845 155 865
rect 10 760 30 780
rect 50 760 70 780
rect 90 760 110 780
rect 130 760 155 780
rect 10 680 30 700
rect 50 680 70 700
rect 90 680 110 700
rect 130 680 155 700
rect 10 600 30 620
rect 50 600 70 620
rect 90 600 110 620
rect 130 600 155 620
rect 10 515 30 535
rect 50 515 70 535
rect 90 515 110 535
rect 130 515 155 535
rect 10 435 30 455
rect 50 435 70 455
rect 90 435 110 455
rect 130 435 155 455
rect 10 355 30 375
rect 50 355 70 375
rect 90 355 110 375
rect 130 355 155 375
rect 10 270 30 290
rect 50 270 70 290
rect 90 270 110 290
rect 130 270 155 290
rect 10 190 30 210
rect 50 190 70 210
rect 90 190 110 210
rect 130 190 155 210
rect 10 110 30 130
rect 50 110 70 130
rect 90 110 110 130
rect 130 110 155 130
rect -60 -285 -40 -260
rect -20 -285 0 -260
rect 20 -285 40 -260
rect 60 -285 85 -260
rect -60 -380 -40 -355
rect -20 -380 0 -355
rect 20 -380 40 -355
rect 60 -380 85 -355
rect -60 -475 -40 -450
rect -20 -475 0 -450
rect 20 -475 40 -450
rect 60 -475 85 -450
rect -60 -570 -40 -545
rect -20 -570 0 -545
rect 20 -570 40 -545
rect 60 -570 85 -545
rect -60 -665 -40 -640
rect -20 -665 0 -640
rect 20 -665 40 -640
rect 60 -665 85 -640
rect -60 -760 -40 -735
rect -20 -760 0 -735
rect 20 -760 40 -735
rect 60 -760 85 -735
rect -60 -855 -40 -830
rect -20 -855 0 -830
rect 20 -855 40 -830
rect 60 -855 85 -830
rect -60 -950 -40 -925
rect -20 -950 0 -925
rect 20 -950 40 -925
rect 60 -950 85 -925
rect -60 -1045 -40 -1020
rect -20 -1045 0 -1020
rect 20 -1045 40 -1020
rect 60 -1045 85 -1020
rect -60 -1140 -40 -1115
rect -20 -1140 0 -1115
rect 20 -1140 40 -1115
rect 60 -1140 85 -1115
rect -60 -1235 -40 -1210
rect -20 -1235 0 -1210
rect 20 -1235 40 -1210
rect 60 -1235 85 -1210
rect -60 -1330 -40 -1305
rect -20 -1330 0 -1305
rect 20 -1330 40 -1305
rect 60 -1330 85 -1305
rect -60 -1425 -40 -1400
rect -20 -1425 0 -1400
rect 20 -1425 40 -1400
rect 60 -1425 85 -1400
rect -60 -1520 -40 -1495
rect -20 -1520 0 -1495
rect 20 -1520 40 -1495
rect 60 -1520 85 -1495
rect -60 -1615 -40 -1590
rect -20 -1615 0 -1590
rect 20 -1615 40 -1590
rect 60 -1615 85 -1590
rect -60 -1710 -40 -1685
rect -20 -1710 0 -1685
rect 20 -1710 40 -1685
rect 60 -1710 85 -1685
rect -60 -1805 -40 -1780
rect -20 -1805 0 -1780
rect 20 -1805 40 -1780
rect 60 -1805 85 -1780
rect -60 -1900 -40 -1875
rect -20 -1900 0 -1875
rect 20 -1900 40 -1875
rect 60 -1900 85 -1875
rect -60 -1995 -40 -1970
rect -20 -1995 0 -1970
rect 20 -1995 40 -1970
rect 60 -1995 85 -1970
rect -60 -2090 -40 -2065
rect -20 -2090 0 -2065
rect 20 -2090 40 -2065
rect 60 -2090 85 -2065
rect -60 -2185 -40 -2160
rect -20 -2185 0 -2160
rect 20 -2185 40 -2160
rect 60 -2185 85 -2160
rect -60 -2280 -40 -2255
rect -20 -2280 0 -2255
rect 20 -2280 40 -2255
rect 60 -2280 85 -2255
rect -60 -2375 -40 -2350
rect -20 -2375 0 -2350
rect 20 -2375 40 -2350
rect 60 -2375 85 -2350
rect -60 -2470 -40 -2445
rect -20 -2470 0 -2445
rect 20 -2470 40 -2445
rect 60 -2470 85 -2445
rect -60 -2565 -40 -2540
rect -20 -2565 0 -2540
rect 20 -2565 40 -2540
rect 60 -2565 85 -2540
rect -60 -2660 -40 -2635
rect -20 -2660 0 -2635
rect 20 -2660 40 -2635
rect 60 -2660 85 -2635
<< locali >>
rect -75 2345 2785 2360
rect -75 2325 -20 2345
rect 0 2325 20 2345
rect 40 2325 60 2345
rect 80 2325 100 2345
rect 120 2325 140 2345
rect 160 2325 180 2345
rect 200 2325 220 2345
rect 240 2325 260 2345
rect 280 2325 300 2345
rect 320 2325 340 2345
rect 360 2325 380 2345
rect 400 2325 420 2345
rect 440 2325 460 2345
rect 480 2325 500 2345
rect 520 2325 540 2345
rect 560 2325 580 2345
rect 600 2325 620 2345
rect 640 2325 660 2345
rect 680 2325 700 2345
rect 720 2325 740 2345
rect 760 2325 780 2345
rect 800 2325 820 2345
rect 840 2325 860 2345
rect 880 2325 900 2345
rect 920 2325 940 2345
rect 960 2325 980 2345
rect 1000 2325 1020 2345
rect 1040 2325 1060 2345
rect 1080 2325 1100 2345
rect 1120 2325 1140 2345
rect 1160 2325 1180 2345
rect 1200 2325 1220 2345
rect 1240 2325 1260 2345
rect 1280 2325 1300 2345
rect 1320 2325 1340 2345
rect 1360 2325 1380 2345
rect 1400 2325 1420 2345
rect 1440 2325 1460 2345
rect 1480 2325 1500 2345
rect 1520 2325 1540 2345
rect 1560 2325 1580 2345
rect 1600 2325 1620 2345
rect 1640 2325 1660 2345
rect 1680 2325 1700 2345
rect 1720 2325 1740 2345
rect 1760 2325 1780 2345
rect 1800 2325 1820 2345
rect 1840 2325 1860 2345
rect 1880 2325 1900 2345
rect 1920 2325 1940 2345
rect 1960 2325 1980 2345
rect 2000 2325 2020 2345
rect 2040 2325 2060 2345
rect 2080 2325 2100 2345
rect 2120 2325 2140 2345
rect 2160 2325 2180 2345
rect 2200 2325 2220 2345
rect 2240 2325 2260 2345
rect 2280 2325 2300 2345
rect 2320 2325 2340 2345
rect 2360 2325 2380 2345
rect 2400 2325 2420 2345
rect 2440 2325 2460 2345
rect 2480 2325 2500 2345
rect 2520 2325 2540 2345
rect 2560 2325 2580 2345
rect 2600 2325 2620 2345
rect 2640 2325 2660 2345
rect 2680 2325 2700 2345
rect 2720 2325 2785 2345
rect -75 2310 2785 2325
rect -75 2290 -60 2310
rect -40 2290 -25 2310
rect -75 2270 -25 2290
rect 2735 2290 2750 2310
rect 2770 2290 2785 2310
rect 2735 2270 2785 2290
rect -75 2250 -60 2270
rect -40 2250 -25 2270
rect -75 2230 -25 2250
rect -75 2210 -60 2230
rect -40 2210 -25 2230
rect -75 2190 -25 2210
rect -75 2170 -60 2190
rect -40 2170 -25 2190
rect 175 2260 2675 2270
rect 175 2240 200 2260
rect 220 2240 240 2260
rect 260 2240 280 2260
rect 300 2240 320 2260
rect 340 2240 360 2260
rect 380 2240 400 2260
rect 420 2240 440 2260
rect 460 2240 480 2260
rect 500 2240 520 2260
rect 540 2240 560 2260
rect 580 2240 600 2260
rect 620 2240 640 2260
rect 660 2240 680 2260
rect 700 2240 720 2260
rect 740 2240 760 2260
rect 780 2240 800 2260
rect 820 2240 840 2260
rect 860 2240 880 2260
rect 900 2240 920 2260
rect 940 2240 960 2260
rect 980 2240 1000 2260
rect 1020 2240 1040 2260
rect 1060 2240 1080 2260
rect 1100 2240 1120 2260
rect 1140 2240 1160 2260
rect 1180 2240 1200 2260
rect 1220 2240 1240 2260
rect 1260 2240 1280 2260
rect 1300 2240 1320 2260
rect 1340 2240 1360 2260
rect 1380 2240 1400 2260
rect 1420 2240 1440 2260
rect 1460 2240 1480 2260
rect 1500 2240 1520 2260
rect 1540 2240 1560 2260
rect 1580 2240 1600 2260
rect 1620 2240 1640 2260
rect 1660 2240 1680 2260
rect 1700 2240 1720 2260
rect 1740 2240 1760 2260
rect 1780 2240 1800 2260
rect 1820 2240 1840 2260
rect 1860 2240 1880 2260
rect 1900 2240 1920 2260
rect 1940 2240 1960 2260
rect 1980 2240 2000 2260
rect 2020 2240 2040 2260
rect 2060 2240 2080 2260
rect 2100 2240 2120 2260
rect 2140 2240 2160 2260
rect 2180 2240 2200 2260
rect 2220 2240 2240 2260
rect 2260 2240 2280 2260
rect 2300 2240 2320 2260
rect 2340 2240 2360 2260
rect 2380 2240 2400 2260
rect 2420 2240 2440 2260
rect 2460 2240 2480 2260
rect 2500 2240 2520 2260
rect 2540 2240 2560 2260
rect 2580 2240 2600 2260
rect 2620 2240 2640 2260
rect 2660 2240 2675 2260
rect 175 2217 2675 2240
rect 175 2197 200 2217
rect 220 2197 240 2217
rect 260 2197 280 2217
rect 300 2197 320 2217
rect 340 2197 360 2217
rect 380 2197 400 2217
rect 420 2197 440 2217
rect 460 2197 480 2217
rect 500 2197 520 2217
rect 540 2197 560 2217
rect 580 2197 600 2217
rect 620 2197 640 2217
rect 660 2197 680 2217
rect 700 2197 720 2217
rect 740 2197 760 2217
rect 780 2197 800 2217
rect 820 2197 840 2217
rect 860 2197 880 2217
rect 900 2197 920 2217
rect 940 2197 960 2217
rect 980 2197 1000 2217
rect 1020 2197 1040 2217
rect 1060 2197 1080 2217
rect 1100 2197 1120 2217
rect 1140 2197 1160 2217
rect 1180 2197 1200 2217
rect 1220 2197 1240 2217
rect 1260 2197 1280 2217
rect 1300 2197 1320 2217
rect 1340 2197 1360 2217
rect 1380 2197 1400 2217
rect 1420 2197 1440 2217
rect 1460 2197 1480 2217
rect 1500 2197 1520 2217
rect 1540 2197 1560 2217
rect 1580 2197 1600 2217
rect 1620 2197 1640 2217
rect 1660 2197 1680 2217
rect 1700 2197 1720 2217
rect 1740 2197 1760 2217
rect 1780 2197 1800 2217
rect 1820 2197 1840 2217
rect 1860 2197 1880 2217
rect 1900 2197 1920 2217
rect 1940 2197 1960 2217
rect 1980 2197 2000 2217
rect 2020 2197 2040 2217
rect 2060 2197 2080 2217
rect 2100 2197 2120 2217
rect 2140 2197 2160 2217
rect 2180 2197 2200 2217
rect 2220 2197 2240 2217
rect 2260 2197 2280 2217
rect 2300 2197 2320 2217
rect 2340 2197 2360 2217
rect 2380 2197 2400 2217
rect 2420 2197 2440 2217
rect 2460 2197 2480 2217
rect 2500 2197 2520 2217
rect 2540 2197 2560 2217
rect 2580 2197 2600 2217
rect 2620 2197 2640 2217
rect 2660 2197 2675 2217
rect 175 2187 2675 2197
rect 2735 2250 2750 2270
rect 2770 2250 2785 2270
rect 2735 2230 2785 2250
rect 2735 2210 2750 2230
rect 2770 2210 2785 2230
rect 2735 2190 2785 2210
rect -75 2150 -25 2170
rect -75 2130 -60 2150
rect -40 2130 -25 2150
rect 0 2175 155 2185
rect 0 2155 10 2175
rect 30 2155 50 2175
rect 70 2155 90 2175
rect 110 2155 130 2175
rect 0 2145 155 2155
rect 2735 2170 2750 2190
rect 2770 2170 2785 2190
rect 2735 2150 2785 2170
rect -75 2110 -25 2130
rect -75 2090 -60 2110
rect -40 2090 -25 2110
rect 175 2135 2675 2145
rect 175 2115 200 2135
rect 220 2115 240 2135
rect 260 2115 280 2135
rect 300 2115 320 2135
rect 340 2115 360 2135
rect 380 2115 400 2135
rect 420 2115 440 2135
rect 460 2115 480 2135
rect 500 2115 520 2135
rect 540 2115 560 2135
rect 580 2115 600 2135
rect 620 2115 640 2135
rect 660 2115 680 2135
rect 700 2115 720 2135
rect 740 2115 760 2135
rect 780 2115 800 2135
rect 820 2115 840 2135
rect 860 2115 880 2135
rect 900 2115 920 2135
rect 940 2115 960 2135
rect 980 2115 1000 2135
rect 1020 2115 1040 2135
rect 1060 2115 1080 2135
rect 1100 2115 1120 2135
rect 1140 2115 1160 2135
rect 1180 2115 1200 2135
rect 1220 2115 1240 2135
rect 1260 2115 1280 2135
rect 1300 2115 1320 2135
rect 1340 2115 1360 2135
rect 1380 2115 1400 2135
rect 1420 2115 1440 2135
rect 1460 2115 1480 2135
rect 1500 2115 1520 2135
rect 1540 2115 1560 2135
rect 1580 2115 1600 2135
rect 1620 2115 1640 2135
rect 1660 2115 1680 2135
rect 1700 2115 1720 2135
rect 1740 2115 1760 2135
rect 1780 2115 1800 2135
rect 1820 2115 1840 2135
rect 1860 2115 1880 2135
rect 1900 2115 1920 2135
rect 1940 2115 1960 2135
rect 1980 2115 2000 2135
rect 2020 2115 2040 2135
rect 2060 2115 2080 2135
rect 2100 2115 2120 2135
rect 2140 2115 2160 2135
rect 2180 2115 2200 2135
rect 2220 2115 2240 2135
rect 2260 2115 2280 2135
rect 2300 2115 2320 2135
rect 2340 2115 2360 2135
rect 2380 2115 2400 2135
rect 2420 2115 2440 2135
rect 2460 2115 2480 2135
rect 2500 2115 2520 2135
rect 2540 2115 2560 2135
rect 2580 2115 2600 2135
rect 2620 2115 2640 2135
rect 2660 2115 2675 2135
rect 175 2105 2675 2115
rect 2735 2130 2750 2150
rect 2770 2130 2785 2150
rect 2735 2110 2785 2130
rect -75 2070 -25 2090
rect -75 2050 -60 2070
rect -40 2050 -25 2070
rect 0 2095 155 2105
rect 0 2075 10 2095
rect 30 2075 50 2095
rect 70 2075 90 2095
rect 110 2075 130 2095
rect 0 2065 155 2075
rect 2735 2090 2750 2110
rect 2770 2090 2785 2110
rect 2735 2070 2785 2090
rect -75 2030 -25 2050
rect -75 2010 -60 2030
rect -40 2010 -25 2030
rect 175 2053 2675 2063
rect 175 2033 200 2053
rect 220 2033 240 2053
rect 260 2033 280 2053
rect 300 2033 320 2053
rect 340 2033 360 2053
rect 380 2033 400 2053
rect 420 2033 440 2053
rect 460 2033 480 2053
rect 500 2033 520 2053
rect 540 2033 560 2053
rect 580 2033 600 2053
rect 620 2033 640 2053
rect 660 2033 680 2053
rect 700 2033 720 2053
rect 740 2033 760 2053
rect 780 2033 800 2053
rect 820 2033 840 2053
rect 860 2033 880 2053
rect 900 2033 920 2053
rect 940 2033 960 2053
rect 980 2033 1000 2053
rect 1020 2033 1040 2053
rect 1060 2033 1080 2053
rect 1100 2033 1120 2053
rect 1140 2033 1160 2053
rect 1180 2033 1200 2053
rect 1220 2033 1240 2053
rect 1260 2033 1280 2053
rect 1300 2033 1320 2053
rect 1340 2033 1360 2053
rect 1380 2033 1400 2053
rect 1420 2033 1440 2053
rect 1460 2033 1480 2053
rect 1500 2033 1520 2053
rect 1540 2033 1560 2053
rect 1580 2033 1600 2053
rect 1620 2033 1640 2053
rect 1660 2033 1680 2053
rect 1700 2033 1720 2053
rect 1740 2033 1760 2053
rect 1780 2033 1800 2053
rect 1820 2033 1840 2053
rect 1860 2033 1880 2053
rect 1900 2033 1920 2053
rect 1940 2033 1960 2053
rect 1980 2033 2000 2053
rect 2020 2033 2040 2053
rect 2060 2033 2080 2053
rect 2100 2033 2120 2053
rect 2140 2033 2160 2053
rect 2180 2033 2200 2053
rect 2220 2033 2240 2053
rect 2260 2033 2280 2053
rect 2300 2033 2320 2053
rect 2340 2033 2360 2053
rect 2380 2033 2400 2053
rect 2420 2033 2440 2053
rect 2460 2033 2480 2053
rect 2500 2033 2520 2053
rect 2540 2033 2560 2053
rect 2580 2033 2600 2053
rect 2620 2033 2640 2053
rect 2660 2033 2675 2053
rect 175 2023 2675 2033
rect 2735 2050 2750 2070
rect 2770 2050 2785 2070
rect 2735 2030 2785 2050
rect -75 1990 -25 2010
rect -75 1970 -60 1990
rect -40 1970 -25 1990
rect 0 2010 155 2020
rect 0 1990 10 2010
rect 30 1990 50 2010
rect 70 1990 90 2010
rect 110 1990 130 2010
rect 0 1980 155 1990
rect 2735 2010 2750 2030
rect 2770 2010 2785 2030
rect 2735 1990 2785 2010
rect -75 1950 -25 1970
rect -75 1930 -60 1950
rect -40 1930 -25 1950
rect 175 1971 2675 1981
rect 175 1951 200 1971
rect 220 1951 240 1971
rect 260 1951 280 1971
rect 300 1951 320 1971
rect 340 1951 360 1971
rect 380 1951 400 1971
rect 420 1951 440 1971
rect 460 1951 480 1971
rect 500 1951 520 1971
rect 540 1951 560 1971
rect 580 1951 600 1971
rect 620 1951 640 1971
rect 660 1951 680 1971
rect 700 1951 720 1971
rect 740 1951 760 1971
rect 780 1951 800 1971
rect 820 1951 840 1971
rect 860 1951 880 1971
rect 900 1951 920 1971
rect 940 1951 960 1971
rect 980 1951 1000 1971
rect 1020 1951 1040 1971
rect 1060 1951 1080 1971
rect 1100 1951 1120 1971
rect 1140 1951 1160 1971
rect 1180 1951 1200 1971
rect 1220 1951 1240 1971
rect 1260 1951 1280 1971
rect 1300 1951 1320 1971
rect 1340 1951 1360 1971
rect 1380 1951 1400 1971
rect 1420 1951 1440 1971
rect 1460 1951 1480 1971
rect 1500 1951 1520 1971
rect 1540 1951 1560 1971
rect 1580 1951 1600 1971
rect 1620 1951 1640 1971
rect 1660 1951 1680 1971
rect 1700 1951 1720 1971
rect 1740 1951 1760 1971
rect 1780 1951 1800 1971
rect 1820 1951 1840 1971
rect 1860 1951 1880 1971
rect 1900 1951 1920 1971
rect 1940 1951 1960 1971
rect 1980 1951 2000 1971
rect 2020 1951 2040 1971
rect 2060 1951 2080 1971
rect 2100 1951 2120 1971
rect 2140 1951 2160 1971
rect 2180 1951 2200 1971
rect 2220 1951 2240 1971
rect 2260 1951 2280 1971
rect 2300 1951 2320 1971
rect 2340 1951 2360 1971
rect 2380 1951 2400 1971
rect 2420 1951 2440 1971
rect 2460 1951 2480 1971
rect 2500 1951 2520 1971
rect 2540 1951 2560 1971
rect 2580 1951 2600 1971
rect 2620 1951 2640 1971
rect 2660 1951 2675 1971
rect 175 1941 2675 1951
rect 2735 1970 2750 1990
rect 2770 1970 2785 1990
rect 2735 1950 2785 1970
rect -75 1910 -25 1930
rect -75 1890 -60 1910
rect -40 1890 -25 1910
rect 0 1930 155 1940
rect 0 1910 10 1930
rect 30 1910 50 1930
rect 70 1910 90 1930
rect 110 1910 130 1930
rect 0 1900 155 1910
rect 2735 1930 2750 1950
rect 2770 1930 2785 1950
rect 2735 1910 2785 1930
rect -75 1870 -25 1890
rect -75 1850 -60 1870
rect -40 1850 -25 1870
rect 175 1889 2675 1899
rect 175 1869 200 1889
rect 220 1869 240 1889
rect 260 1869 280 1889
rect 300 1869 320 1889
rect 340 1869 360 1889
rect 380 1869 400 1889
rect 420 1869 440 1889
rect 460 1869 480 1889
rect 500 1869 520 1889
rect 540 1869 560 1889
rect 580 1869 600 1889
rect 620 1869 640 1889
rect 660 1869 680 1889
rect 700 1869 720 1889
rect 740 1869 760 1889
rect 780 1869 800 1889
rect 820 1869 840 1889
rect 860 1869 880 1889
rect 900 1869 920 1889
rect 940 1869 960 1889
rect 980 1869 1000 1889
rect 1020 1869 1040 1889
rect 1060 1869 1080 1889
rect 1100 1869 1120 1889
rect 1140 1869 1160 1889
rect 1180 1869 1200 1889
rect 1220 1869 1240 1889
rect 1260 1869 1280 1889
rect 1300 1869 1320 1889
rect 1340 1869 1360 1889
rect 1380 1869 1400 1889
rect 1420 1869 1440 1889
rect 1460 1869 1480 1889
rect 1500 1869 1520 1889
rect 1540 1869 1560 1889
rect 1580 1869 1600 1889
rect 1620 1869 1640 1889
rect 1660 1869 1680 1889
rect 1700 1869 1720 1889
rect 1740 1869 1760 1889
rect 1780 1869 1800 1889
rect 1820 1869 1840 1889
rect 1860 1869 1880 1889
rect 1900 1869 1920 1889
rect 1940 1869 1960 1889
rect 1980 1869 2000 1889
rect 2020 1869 2040 1889
rect 2060 1869 2080 1889
rect 2100 1869 2120 1889
rect 2140 1869 2160 1889
rect 2180 1869 2200 1889
rect 2220 1869 2240 1889
rect 2260 1869 2280 1889
rect 2300 1869 2320 1889
rect 2340 1869 2360 1889
rect 2380 1869 2400 1889
rect 2420 1869 2440 1889
rect 2460 1869 2480 1889
rect 2500 1869 2520 1889
rect 2540 1869 2560 1889
rect 2580 1869 2600 1889
rect 2620 1869 2640 1889
rect 2660 1869 2675 1889
rect -75 1830 -25 1850
rect -75 1810 -60 1830
rect -40 1810 -25 1830
rect 0 1850 155 1860
rect 175 1859 2675 1869
rect 2735 1890 2750 1910
rect 2770 1890 2785 1910
rect 2735 1870 2785 1890
rect 0 1830 10 1850
rect 30 1830 50 1850
rect 70 1830 90 1850
rect 110 1830 130 1850
rect 0 1820 155 1830
rect 2735 1850 2750 1870
rect 2770 1850 2785 1870
rect 2735 1830 2785 1850
rect -75 1790 -25 1810
rect -75 1770 -60 1790
rect -40 1770 -25 1790
rect 175 1807 2675 1817
rect 175 1787 200 1807
rect 220 1787 240 1807
rect 260 1787 280 1807
rect 300 1787 320 1807
rect 340 1787 360 1807
rect 380 1787 400 1807
rect 420 1787 440 1807
rect 460 1787 480 1807
rect 500 1787 520 1807
rect 540 1787 560 1807
rect 580 1787 600 1807
rect 620 1787 640 1807
rect 660 1787 680 1807
rect 700 1787 720 1807
rect 740 1787 760 1807
rect 780 1787 800 1807
rect 820 1787 840 1807
rect 860 1787 880 1807
rect 900 1787 920 1807
rect 940 1787 960 1807
rect 980 1787 1000 1807
rect 1020 1787 1040 1807
rect 1060 1787 1080 1807
rect 1100 1787 1120 1807
rect 1140 1787 1160 1807
rect 1180 1787 1200 1807
rect 1220 1787 1240 1807
rect 1260 1787 1280 1807
rect 1300 1787 1320 1807
rect 1340 1787 1360 1807
rect 1380 1787 1400 1807
rect 1420 1787 1440 1807
rect 1460 1787 1480 1807
rect 1500 1787 1520 1807
rect 1540 1787 1560 1807
rect 1580 1787 1600 1807
rect 1620 1787 1640 1807
rect 1660 1787 1680 1807
rect 1700 1787 1720 1807
rect 1740 1787 1760 1807
rect 1780 1787 1800 1807
rect 1820 1787 1840 1807
rect 1860 1787 1880 1807
rect 1900 1787 1920 1807
rect 1940 1787 1960 1807
rect 1980 1787 2000 1807
rect 2020 1787 2040 1807
rect 2060 1787 2080 1807
rect 2100 1787 2120 1807
rect 2140 1787 2160 1807
rect 2180 1787 2200 1807
rect 2220 1787 2240 1807
rect 2260 1787 2280 1807
rect 2300 1787 2320 1807
rect 2340 1787 2360 1807
rect 2380 1787 2400 1807
rect 2420 1787 2440 1807
rect 2460 1787 2480 1807
rect 2500 1787 2520 1807
rect 2540 1787 2560 1807
rect 2580 1787 2600 1807
rect 2620 1787 2640 1807
rect 2660 1787 2675 1807
rect 175 1777 2675 1787
rect 2735 1810 2750 1830
rect 2770 1810 2785 1830
rect 2735 1790 2785 1810
rect -75 1750 -25 1770
rect -75 1730 -60 1750
rect -40 1730 -25 1750
rect 0 1765 155 1775
rect 0 1745 10 1765
rect 30 1745 50 1765
rect 70 1745 90 1765
rect 110 1745 130 1765
rect 0 1735 155 1745
rect 2735 1770 2750 1790
rect 2770 1770 2785 1790
rect 2735 1750 2785 1770
rect -75 1710 -25 1730
rect -75 1690 -60 1710
rect -40 1690 -25 1710
rect 175 1725 2675 1735
rect 175 1705 200 1725
rect 220 1705 240 1725
rect 260 1705 280 1725
rect 300 1705 320 1725
rect 340 1705 360 1725
rect 380 1705 400 1725
rect 420 1705 440 1725
rect 460 1705 480 1725
rect 500 1705 520 1725
rect 540 1705 560 1725
rect 580 1705 600 1725
rect 620 1705 640 1725
rect 660 1705 680 1725
rect 700 1705 720 1725
rect 740 1705 760 1725
rect 780 1705 800 1725
rect 820 1705 840 1725
rect 860 1705 880 1725
rect 900 1705 920 1725
rect 940 1705 960 1725
rect 980 1705 1000 1725
rect 1020 1705 1040 1725
rect 1060 1705 1080 1725
rect 1100 1705 1120 1725
rect 1140 1705 1160 1725
rect 1180 1705 1200 1725
rect 1220 1705 1240 1725
rect 1260 1705 1280 1725
rect 1300 1705 1320 1725
rect 1340 1705 1360 1725
rect 1380 1705 1400 1725
rect 1420 1705 1440 1725
rect 1460 1705 1480 1725
rect 1500 1705 1520 1725
rect 1540 1705 1560 1725
rect 1580 1705 1600 1725
rect 1620 1705 1640 1725
rect 1660 1705 1680 1725
rect 1700 1705 1720 1725
rect 1740 1705 1760 1725
rect 1780 1705 1800 1725
rect 1820 1705 1840 1725
rect 1860 1705 1880 1725
rect 1900 1705 1920 1725
rect 1940 1705 1960 1725
rect 1980 1705 2000 1725
rect 2020 1705 2040 1725
rect 2060 1705 2080 1725
rect 2100 1705 2120 1725
rect 2140 1705 2160 1725
rect 2180 1705 2200 1725
rect 2220 1705 2240 1725
rect 2260 1705 2280 1725
rect 2300 1705 2320 1725
rect 2340 1705 2360 1725
rect 2380 1705 2400 1725
rect 2420 1705 2440 1725
rect 2460 1705 2480 1725
rect 2500 1705 2520 1725
rect 2540 1705 2560 1725
rect 2580 1705 2600 1725
rect 2620 1705 2640 1725
rect 2660 1705 2675 1725
rect 175 1695 2675 1705
rect 2735 1730 2750 1750
rect 2770 1730 2785 1750
rect 2735 1710 2785 1730
rect -75 1670 -25 1690
rect -75 1650 -60 1670
rect -40 1650 -25 1670
rect 0 1685 155 1695
rect 0 1665 10 1685
rect 30 1665 50 1685
rect 70 1665 90 1685
rect 110 1665 130 1685
rect 0 1655 155 1665
rect 2735 1690 2750 1710
rect 2770 1690 2785 1710
rect 2735 1670 2785 1690
rect -75 1630 -25 1650
rect -75 1610 -60 1630
rect -40 1610 -25 1630
rect 175 1643 2675 1653
rect 175 1623 200 1643
rect 220 1623 240 1643
rect 260 1623 280 1643
rect 300 1623 320 1643
rect 340 1623 360 1643
rect 380 1623 400 1643
rect 420 1623 440 1643
rect 460 1623 480 1643
rect 500 1623 520 1643
rect 540 1623 560 1643
rect 580 1623 600 1643
rect 620 1623 640 1643
rect 660 1623 680 1643
rect 700 1623 720 1643
rect 740 1623 760 1643
rect 780 1623 800 1643
rect 820 1623 840 1643
rect 860 1623 880 1643
rect 900 1623 920 1643
rect 940 1623 960 1643
rect 980 1623 1000 1643
rect 1020 1623 1040 1643
rect 1060 1623 1080 1643
rect 1100 1623 1120 1643
rect 1140 1623 1160 1643
rect 1180 1623 1200 1643
rect 1220 1623 1240 1643
rect 1260 1623 1280 1643
rect 1300 1623 1320 1643
rect 1340 1623 1360 1643
rect 1380 1623 1400 1643
rect 1420 1623 1440 1643
rect 1460 1623 1480 1643
rect 1500 1623 1520 1643
rect 1540 1623 1560 1643
rect 1580 1623 1600 1643
rect 1620 1623 1640 1643
rect 1660 1623 1680 1643
rect 1700 1623 1720 1643
rect 1740 1623 1760 1643
rect 1780 1623 1800 1643
rect 1820 1623 1840 1643
rect 1860 1623 1880 1643
rect 1900 1623 1920 1643
rect 1940 1623 1960 1643
rect 1980 1623 2000 1643
rect 2020 1623 2040 1643
rect 2060 1623 2080 1643
rect 2100 1623 2120 1643
rect 2140 1623 2160 1643
rect 2180 1623 2200 1643
rect 2220 1623 2240 1643
rect 2260 1623 2280 1643
rect 2300 1623 2320 1643
rect 2340 1623 2360 1643
rect 2380 1623 2400 1643
rect 2420 1623 2440 1643
rect 2460 1623 2480 1643
rect 2500 1623 2520 1643
rect 2540 1623 2560 1643
rect 2580 1623 2600 1643
rect 2620 1623 2640 1643
rect 2660 1623 2675 1643
rect 175 1613 2675 1623
rect 2735 1650 2750 1670
rect 2770 1650 2785 1670
rect 2735 1630 2785 1650
rect 2735 1610 2750 1630
rect 2770 1610 2785 1630
rect -75 1590 -25 1610
rect -75 1570 -60 1590
rect -40 1570 -25 1590
rect 0 1600 155 1610
rect 0 1580 10 1600
rect 30 1580 50 1600
rect 70 1580 90 1600
rect 110 1580 130 1600
rect 0 1570 155 1580
rect 2735 1590 2785 1610
rect -75 1550 -25 1570
rect -75 1530 -60 1550
rect -40 1530 -25 1550
rect 175 1561 2675 1571
rect 175 1541 200 1561
rect 220 1541 240 1561
rect 260 1541 280 1561
rect 300 1541 320 1561
rect 340 1541 360 1561
rect 380 1541 400 1561
rect 420 1541 440 1561
rect 460 1541 480 1561
rect 500 1541 520 1561
rect 540 1541 560 1561
rect 580 1541 600 1561
rect 620 1541 640 1561
rect 660 1541 680 1561
rect 700 1541 720 1561
rect 740 1541 760 1561
rect 780 1541 800 1561
rect 820 1541 840 1561
rect 860 1541 880 1561
rect 900 1541 920 1561
rect 940 1541 960 1561
rect 980 1541 1000 1561
rect 1020 1541 1040 1561
rect 1060 1541 1080 1561
rect 1100 1541 1120 1561
rect 1140 1541 1160 1561
rect 1180 1541 1200 1561
rect 1220 1541 1240 1561
rect 1260 1541 1280 1561
rect 1300 1541 1320 1561
rect 1340 1541 1360 1561
rect 1380 1541 1400 1561
rect 1420 1541 1440 1561
rect 1460 1541 1480 1561
rect 1500 1541 1520 1561
rect 1540 1541 1560 1561
rect 1580 1541 1600 1561
rect 1620 1541 1640 1561
rect 1660 1541 1680 1561
rect 1700 1541 1720 1561
rect 1740 1541 1760 1561
rect 1780 1541 1800 1561
rect 1820 1541 1840 1561
rect 1860 1541 1880 1561
rect 1900 1541 1920 1561
rect 1940 1541 1960 1561
rect 1980 1541 2000 1561
rect 2020 1541 2040 1561
rect 2060 1541 2080 1561
rect 2100 1541 2120 1561
rect 2140 1541 2160 1561
rect 2180 1541 2200 1561
rect 2220 1541 2240 1561
rect 2260 1541 2280 1561
rect 2300 1541 2320 1561
rect 2340 1541 2360 1561
rect 2380 1541 2400 1561
rect 2420 1541 2440 1561
rect 2460 1541 2480 1561
rect 2500 1541 2520 1561
rect 2540 1541 2560 1561
rect 2580 1541 2600 1561
rect 2620 1541 2640 1561
rect 2660 1541 2675 1561
rect 175 1531 2675 1541
rect 2735 1570 2750 1590
rect 2770 1570 2785 1590
rect 2735 1550 2785 1570
rect 2735 1530 2750 1550
rect 2770 1530 2785 1550
rect -75 1510 -25 1530
rect -75 1490 -60 1510
rect -40 1490 -25 1510
rect 0 1520 155 1530
rect 0 1500 10 1520
rect 30 1500 50 1520
rect 70 1500 90 1520
rect 110 1500 130 1520
rect 0 1490 155 1500
rect 2735 1510 2785 1530
rect 2735 1490 2750 1510
rect 2770 1490 2785 1510
rect -75 1470 -25 1490
rect -75 1450 -60 1470
rect -40 1450 -25 1470
rect 175 1479 2675 1489
rect 175 1459 200 1479
rect 220 1459 240 1479
rect 260 1459 280 1479
rect 300 1459 320 1479
rect 340 1459 360 1479
rect 380 1459 400 1479
rect 420 1459 440 1479
rect 460 1459 480 1479
rect 500 1459 520 1479
rect 540 1459 560 1479
rect 580 1459 600 1479
rect 620 1459 640 1479
rect 660 1459 680 1479
rect 700 1459 720 1479
rect 740 1459 760 1479
rect 780 1459 800 1479
rect 820 1459 840 1479
rect 860 1459 880 1479
rect 900 1459 920 1479
rect 940 1459 960 1479
rect 980 1459 1000 1479
rect 1020 1459 1040 1479
rect 1060 1459 1080 1479
rect 1100 1459 1120 1479
rect 1140 1459 1160 1479
rect 1180 1459 1200 1479
rect 1220 1459 1240 1479
rect 1260 1459 1280 1479
rect 1300 1459 1320 1479
rect 1340 1459 1360 1479
rect 1380 1459 1400 1479
rect 1420 1459 1440 1479
rect 1460 1459 1480 1479
rect 1500 1459 1520 1479
rect 1540 1459 1560 1479
rect 1580 1459 1600 1479
rect 1620 1459 1640 1479
rect 1660 1459 1680 1479
rect 1700 1459 1720 1479
rect 1740 1459 1760 1479
rect 1780 1459 1800 1479
rect 1820 1459 1840 1479
rect 1860 1459 1880 1479
rect 1900 1459 1920 1479
rect 1940 1459 1960 1479
rect 1980 1459 2000 1479
rect 2020 1459 2040 1479
rect 2060 1459 2080 1479
rect 2100 1459 2120 1479
rect 2140 1459 2160 1479
rect 2180 1459 2200 1479
rect 2220 1459 2240 1479
rect 2260 1459 2280 1479
rect 2300 1459 2320 1479
rect 2340 1459 2360 1479
rect 2380 1459 2400 1479
rect 2420 1459 2440 1479
rect 2460 1459 2480 1479
rect 2500 1459 2520 1479
rect 2540 1459 2560 1479
rect 2580 1459 2600 1479
rect 2620 1459 2640 1479
rect 2660 1459 2675 1479
rect -75 1430 -25 1450
rect -75 1410 -60 1430
rect -40 1410 -25 1430
rect 0 1440 155 1450
rect 175 1449 2675 1459
rect 2735 1470 2785 1490
rect 2735 1450 2750 1470
rect 2770 1450 2785 1470
rect 0 1420 10 1440
rect 30 1420 50 1440
rect 70 1420 90 1440
rect 110 1420 130 1440
rect 0 1410 155 1420
rect 2735 1430 2785 1450
rect 2735 1410 2750 1430
rect 2770 1410 2785 1430
rect -75 1390 -25 1410
rect -75 1370 -60 1390
rect -40 1370 -25 1390
rect -75 1350 -25 1370
rect 175 1397 2675 1407
rect 175 1377 200 1397
rect 220 1377 240 1397
rect 260 1377 280 1397
rect 300 1377 320 1397
rect 340 1377 360 1397
rect 380 1377 400 1397
rect 420 1377 440 1397
rect 460 1377 480 1397
rect 500 1377 520 1397
rect 540 1377 560 1397
rect 580 1377 600 1397
rect 620 1377 640 1397
rect 660 1377 680 1397
rect 700 1377 720 1397
rect 740 1377 760 1397
rect 780 1377 800 1397
rect 820 1377 840 1397
rect 860 1377 880 1397
rect 900 1377 920 1397
rect 940 1377 960 1397
rect 980 1377 1000 1397
rect 1020 1377 1040 1397
rect 1060 1377 1080 1397
rect 1100 1377 1120 1397
rect 1140 1377 1160 1397
rect 1180 1377 1200 1397
rect 1220 1377 1240 1397
rect 1260 1377 1280 1397
rect 1300 1377 1320 1397
rect 1340 1377 1360 1397
rect 1380 1377 1400 1397
rect 1420 1377 1440 1397
rect 1460 1377 1480 1397
rect 1500 1377 1520 1397
rect 1540 1377 1560 1397
rect 1580 1377 1600 1397
rect 1620 1377 1640 1397
rect 1660 1377 1680 1397
rect 1700 1377 1720 1397
rect 1740 1377 1760 1397
rect 1780 1377 1800 1397
rect 1820 1377 1840 1397
rect 1860 1377 1880 1397
rect 1900 1377 1920 1397
rect 1940 1377 1960 1397
rect 1980 1377 2000 1397
rect 2020 1377 2040 1397
rect 2060 1377 2080 1397
rect 2100 1377 2120 1397
rect 2140 1377 2160 1397
rect 2180 1377 2200 1397
rect 2220 1377 2240 1397
rect 2260 1377 2280 1397
rect 2300 1377 2320 1397
rect 2340 1377 2360 1397
rect 2380 1377 2400 1397
rect 2420 1377 2440 1397
rect 2460 1377 2480 1397
rect 2500 1377 2520 1397
rect 2540 1377 2560 1397
rect 2580 1377 2600 1397
rect 2620 1377 2640 1397
rect 2660 1377 2675 1397
rect 175 1367 2675 1377
rect 2735 1390 2785 1410
rect 2735 1370 2750 1390
rect 2770 1370 2785 1390
rect -75 1330 -60 1350
rect -40 1330 -25 1350
rect -75 1310 -25 1330
rect 0 1355 155 1365
rect 0 1335 10 1355
rect 30 1335 50 1355
rect 70 1335 90 1355
rect 110 1335 130 1355
rect 0 1325 155 1335
rect 2735 1350 2785 1370
rect 2735 1330 2750 1350
rect 2770 1330 2785 1350
rect -75 1290 -60 1310
rect -40 1290 -25 1310
rect -75 1270 -25 1290
rect 175 1315 2675 1325
rect 175 1295 200 1315
rect 220 1295 240 1315
rect 260 1295 280 1315
rect 300 1295 320 1315
rect 340 1295 360 1315
rect 380 1295 400 1315
rect 420 1295 440 1315
rect 460 1295 480 1315
rect 500 1295 520 1315
rect 540 1295 560 1315
rect 580 1295 600 1315
rect 620 1295 640 1315
rect 660 1295 680 1315
rect 700 1295 720 1315
rect 740 1295 760 1315
rect 780 1295 800 1315
rect 820 1295 840 1315
rect 860 1295 880 1315
rect 900 1295 920 1315
rect 940 1295 960 1315
rect 980 1295 1000 1315
rect 1020 1295 1040 1315
rect 1060 1295 1080 1315
rect 1100 1295 1120 1315
rect 1140 1295 1160 1315
rect 1180 1295 1200 1315
rect 1220 1295 1240 1315
rect 1260 1295 1280 1315
rect 1300 1295 1320 1315
rect 1340 1295 1360 1315
rect 1380 1295 1400 1315
rect 1420 1295 1440 1315
rect 1460 1295 1480 1315
rect 1500 1295 1520 1315
rect 1540 1295 1560 1315
rect 1580 1295 1600 1315
rect 1620 1295 1640 1315
rect 1660 1295 1680 1315
rect 1700 1295 1720 1315
rect 1740 1295 1760 1315
rect 1780 1295 1800 1315
rect 1820 1295 1840 1315
rect 1860 1295 1880 1315
rect 1900 1295 1920 1315
rect 1940 1295 1960 1315
rect 1980 1295 2000 1315
rect 2020 1295 2040 1315
rect 2060 1295 2080 1315
rect 2100 1295 2120 1315
rect 2140 1295 2160 1315
rect 2180 1295 2200 1315
rect 2220 1295 2240 1315
rect 2260 1295 2280 1315
rect 2300 1295 2320 1315
rect 2340 1295 2360 1315
rect 2380 1295 2400 1315
rect 2420 1295 2440 1315
rect 2460 1295 2480 1315
rect 2500 1295 2520 1315
rect 2540 1295 2560 1315
rect 2580 1295 2600 1315
rect 2620 1295 2640 1315
rect 2660 1295 2675 1315
rect 175 1285 2675 1295
rect 2735 1310 2785 1330
rect 2735 1290 2750 1310
rect 2770 1290 2785 1310
rect -75 1250 -60 1270
rect -40 1250 -25 1270
rect -75 1230 -25 1250
rect 0 1275 155 1285
rect 0 1255 10 1275
rect 30 1255 50 1275
rect 70 1255 90 1275
rect 110 1255 130 1275
rect 0 1245 155 1255
rect 2735 1270 2785 1290
rect 2735 1250 2750 1270
rect 2770 1250 2785 1270
rect -75 1210 -60 1230
rect -40 1210 -25 1230
rect -75 1190 -25 1210
rect 175 1233 2675 1243
rect 175 1213 200 1233
rect 220 1213 240 1233
rect 260 1213 280 1233
rect 300 1213 320 1233
rect 340 1213 360 1233
rect 380 1213 400 1233
rect 420 1213 440 1233
rect 460 1213 480 1233
rect 500 1213 520 1233
rect 540 1213 560 1233
rect 580 1213 600 1233
rect 620 1213 640 1233
rect 660 1213 680 1233
rect 700 1213 720 1233
rect 740 1213 760 1233
rect 780 1213 800 1233
rect 820 1213 840 1233
rect 860 1213 880 1233
rect 900 1213 920 1233
rect 940 1213 960 1233
rect 980 1213 1000 1233
rect 1020 1213 1040 1233
rect 1060 1213 1080 1233
rect 1100 1213 1120 1233
rect 1140 1213 1160 1233
rect 1180 1213 1200 1233
rect 1220 1213 1240 1233
rect 1260 1213 1280 1233
rect 1300 1213 1320 1233
rect 1340 1213 1360 1233
rect 1380 1213 1400 1233
rect 1420 1213 1440 1233
rect 1460 1213 1480 1233
rect 1500 1213 1520 1233
rect 1540 1213 1560 1233
rect 1580 1213 1600 1233
rect 1620 1213 1640 1233
rect 1660 1213 1680 1233
rect 1700 1213 1720 1233
rect 1740 1213 1760 1233
rect 1780 1213 1800 1233
rect 1820 1213 1840 1233
rect 1860 1213 1880 1233
rect 1900 1213 1920 1233
rect 1940 1213 1960 1233
rect 1980 1213 2000 1233
rect 2020 1213 2040 1233
rect 2060 1213 2080 1233
rect 2100 1213 2120 1233
rect 2140 1213 2160 1233
rect 2180 1213 2200 1233
rect 2220 1213 2240 1233
rect 2260 1213 2280 1233
rect 2300 1213 2320 1233
rect 2340 1213 2360 1233
rect 2380 1213 2400 1233
rect 2420 1213 2440 1233
rect 2460 1213 2480 1233
rect 2500 1213 2520 1233
rect 2540 1213 2560 1233
rect 2580 1213 2600 1233
rect 2620 1213 2640 1233
rect 2660 1213 2675 1233
rect 175 1203 2675 1213
rect 2735 1230 2785 1250
rect 2735 1210 2750 1230
rect 2770 1210 2785 1230
rect -75 1170 -60 1190
rect -40 1170 -25 1190
rect -75 1150 -25 1170
rect 0 1190 155 1200
rect 0 1170 10 1190
rect 30 1170 50 1190
rect 70 1170 90 1190
rect 110 1170 130 1190
rect 0 1160 155 1170
rect 2735 1190 2785 1210
rect 2735 1170 2750 1190
rect 2770 1170 2785 1190
rect -75 1130 -60 1150
rect -40 1130 -25 1150
rect -75 1110 -25 1130
rect 175 1151 2675 1161
rect 175 1131 200 1151
rect 220 1131 240 1151
rect 260 1131 280 1151
rect 300 1131 320 1151
rect 340 1131 360 1151
rect 380 1131 400 1151
rect 420 1131 440 1151
rect 460 1131 480 1151
rect 500 1131 520 1151
rect 540 1131 560 1151
rect 580 1131 600 1151
rect 620 1131 640 1151
rect 660 1131 680 1151
rect 700 1131 720 1151
rect 740 1131 760 1151
rect 780 1131 800 1151
rect 820 1131 840 1151
rect 860 1131 880 1151
rect 900 1131 920 1151
rect 940 1131 960 1151
rect 980 1131 1000 1151
rect 1020 1131 1040 1151
rect 1060 1131 1080 1151
rect 1100 1131 1120 1151
rect 1140 1131 1160 1151
rect 1180 1131 1200 1151
rect 1220 1131 1240 1151
rect 1260 1131 1280 1151
rect 1300 1131 1320 1151
rect 1340 1131 1360 1151
rect 1380 1131 1400 1151
rect 1420 1131 1440 1151
rect 1460 1131 1480 1151
rect 1500 1131 1520 1151
rect 1540 1131 1560 1151
rect 1580 1131 1600 1151
rect 1620 1131 1640 1151
rect 1660 1131 1680 1151
rect 1700 1131 1720 1151
rect 1740 1131 1760 1151
rect 1780 1131 1800 1151
rect 1820 1131 1840 1151
rect 1860 1131 1880 1151
rect 1900 1131 1920 1151
rect 1940 1131 1960 1151
rect 1980 1131 2000 1151
rect 2020 1131 2040 1151
rect 2060 1131 2080 1151
rect 2100 1131 2120 1151
rect 2140 1131 2160 1151
rect 2180 1131 2200 1151
rect 2220 1131 2240 1151
rect 2260 1131 2280 1151
rect 2300 1131 2320 1151
rect 2340 1131 2360 1151
rect 2380 1131 2400 1151
rect 2420 1131 2440 1151
rect 2460 1131 2480 1151
rect 2500 1131 2520 1151
rect 2540 1131 2560 1151
rect 2580 1131 2600 1151
rect 2620 1131 2640 1151
rect 2660 1131 2675 1151
rect 175 1121 2675 1131
rect 2735 1150 2785 1170
rect 2735 1130 2750 1150
rect 2770 1130 2785 1150
rect -75 1090 -60 1110
rect -40 1090 -25 1110
rect -75 1070 -25 1090
rect 0 1110 155 1120
rect 0 1090 10 1110
rect 30 1090 50 1110
rect 70 1090 90 1110
rect 110 1090 130 1110
rect 0 1080 155 1090
rect 2735 1110 2785 1130
rect 2735 1090 2750 1110
rect 2770 1090 2785 1110
rect -75 1050 -60 1070
rect -40 1050 -25 1070
rect -75 1030 -25 1050
rect 175 1069 2675 1079
rect 175 1049 200 1069
rect 220 1049 240 1069
rect 260 1049 280 1069
rect 300 1049 320 1069
rect 340 1049 360 1069
rect 380 1049 400 1069
rect 420 1049 440 1069
rect 460 1049 480 1069
rect 500 1049 520 1069
rect 540 1049 560 1069
rect 580 1049 600 1069
rect 620 1049 640 1069
rect 660 1049 680 1069
rect 700 1049 720 1069
rect 740 1049 760 1069
rect 780 1049 800 1069
rect 820 1049 840 1069
rect 860 1049 880 1069
rect 900 1049 920 1069
rect 940 1049 960 1069
rect 980 1049 1000 1069
rect 1020 1049 1040 1069
rect 1060 1049 1080 1069
rect 1100 1049 1120 1069
rect 1140 1049 1160 1069
rect 1180 1049 1200 1069
rect 1220 1049 1240 1069
rect 1260 1049 1280 1069
rect 1300 1049 1320 1069
rect 1340 1049 1360 1069
rect 1380 1049 1400 1069
rect 1420 1049 1440 1069
rect 1460 1049 1480 1069
rect 1500 1049 1520 1069
rect 1540 1049 1560 1069
rect 1580 1049 1600 1069
rect 1620 1049 1640 1069
rect 1660 1049 1680 1069
rect 1700 1049 1720 1069
rect 1740 1049 1760 1069
rect 1780 1049 1800 1069
rect 1820 1049 1840 1069
rect 1860 1049 1880 1069
rect 1900 1049 1920 1069
rect 1940 1049 1960 1069
rect 1980 1049 2000 1069
rect 2020 1049 2040 1069
rect 2060 1049 2080 1069
rect 2100 1049 2120 1069
rect 2140 1049 2160 1069
rect 2180 1049 2200 1069
rect 2220 1049 2240 1069
rect 2260 1049 2280 1069
rect 2300 1049 2320 1069
rect 2340 1049 2360 1069
rect 2380 1049 2400 1069
rect 2420 1049 2440 1069
rect 2460 1049 2480 1069
rect 2500 1049 2520 1069
rect 2540 1049 2560 1069
rect 2580 1049 2600 1069
rect 2620 1049 2640 1069
rect 2660 1049 2675 1069
rect -75 1010 -60 1030
rect -40 1010 -25 1030
rect -75 990 -25 1010
rect 0 1030 155 1040
rect 175 1039 2675 1049
rect 2735 1070 2785 1090
rect 2735 1050 2750 1070
rect 2770 1050 2785 1070
rect 0 1010 10 1030
rect 30 1010 50 1030
rect 70 1010 90 1030
rect 110 1010 130 1030
rect 0 1000 155 1010
rect 2735 1030 2785 1050
rect 2735 1010 2750 1030
rect 2770 1010 2785 1030
rect -75 970 -60 990
rect -40 970 -25 990
rect -75 950 -25 970
rect 175 987 2675 997
rect 175 967 200 987
rect 220 967 240 987
rect 260 967 280 987
rect 300 967 320 987
rect 340 967 360 987
rect 380 967 400 987
rect 420 967 440 987
rect 460 967 480 987
rect 500 967 520 987
rect 540 967 560 987
rect 580 967 600 987
rect 620 967 640 987
rect 660 967 680 987
rect 700 967 720 987
rect 740 967 760 987
rect 780 967 800 987
rect 820 967 840 987
rect 860 967 880 987
rect 900 967 920 987
rect 940 967 960 987
rect 980 967 1000 987
rect 1020 967 1040 987
rect 1060 967 1080 987
rect 1100 967 1120 987
rect 1140 967 1160 987
rect 1180 967 1200 987
rect 1220 967 1240 987
rect 1260 967 1280 987
rect 1300 967 1320 987
rect 1340 967 1360 987
rect 1380 967 1400 987
rect 1420 967 1440 987
rect 1460 967 1480 987
rect 1500 967 1520 987
rect 1540 967 1560 987
rect 1580 967 1600 987
rect 1620 967 1640 987
rect 1660 967 1680 987
rect 1700 967 1720 987
rect 1740 967 1760 987
rect 1780 967 1800 987
rect 1820 967 1840 987
rect 1860 967 1880 987
rect 1900 967 1920 987
rect 1940 967 1960 987
rect 1980 967 2000 987
rect 2020 967 2040 987
rect 2060 967 2080 987
rect 2100 967 2120 987
rect 2140 967 2160 987
rect 2180 967 2200 987
rect 2220 967 2240 987
rect 2260 967 2280 987
rect 2300 967 2320 987
rect 2340 967 2360 987
rect 2380 967 2400 987
rect 2420 967 2440 987
rect 2460 967 2480 987
rect 2500 967 2520 987
rect 2540 967 2560 987
rect 2580 967 2600 987
rect 2620 967 2640 987
rect 2660 967 2675 987
rect 175 957 2675 967
rect 2735 990 2785 1010
rect 2735 970 2750 990
rect 2770 970 2785 990
rect -75 930 -60 950
rect -40 930 -25 950
rect -75 910 -25 930
rect 0 945 155 955
rect 0 925 10 945
rect 30 925 50 945
rect 70 925 90 945
rect 110 925 130 945
rect 0 915 155 925
rect 2735 950 2785 970
rect 2735 930 2750 950
rect 2770 930 2785 950
rect -75 890 -60 910
rect -40 890 -25 910
rect -75 870 -25 890
rect 175 905 2675 915
rect 175 885 200 905
rect 220 885 240 905
rect 260 885 280 905
rect 300 885 320 905
rect 340 885 360 905
rect 380 885 400 905
rect 420 885 440 905
rect 460 885 480 905
rect 500 885 520 905
rect 540 885 560 905
rect 580 885 600 905
rect 620 885 640 905
rect 660 885 680 905
rect 700 885 720 905
rect 740 885 760 905
rect 780 885 800 905
rect 820 885 840 905
rect 860 885 880 905
rect 900 885 920 905
rect 940 885 960 905
rect 980 885 1000 905
rect 1020 885 1040 905
rect 1060 885 1080 905
rect 1100 885 1120 905
rect 1140 885 1160 905
rect 1180 885 1200 905
rect 1220 885 1240 905
rect 1260 885 1280 905
rect 1300 885 1320 905
rect 1340 885 1360 905
rect 1380 885 1400 905
rect 1420 885 1440 905
rect 1460 885 1480 905
rect 1500 885 1520 905
rect 1540 885 1560 905
rect 1580 885 1600 905
rect 1620 885 1640 905
rect 1660 885 1680 905
rect 1700 885 1720 905
rect 1740 885 1760 905
rect 1780 885 1800 905
rect 1820 885 1840 905
rect 1860 885 1880 905
rect 1900 885 1920 905
rect 1940 885 1960 905
rect 1980 885 2000 905
rect 2020 885 2040 905
rect 2060 885 2080 905
rect 2100 885 2120 905
rect 2140 885 2160 905
rect 2180 885 2200 905
rect 2220 885 2240 905
rect 2260 885 2280 905
rect 2300 885 2320 905
rect 2340 885 2360 905
rect 2380 885 2400 905
rect 2420 885 2440 905
rect 2460 885 2480 905
rect 2500 885 2520 905
rect 2540 885 2560 905
rect 2580 885 2600 905
rect 2620 885 2640 905
rect 2660 885 2675 905
rect 175 875 2675 885
rect 2735 910 2785 930
rect 2735 890 2750 910
rect 2770 890 2785 910
rect -75 850 -60 870
rect -40 850 -25 870
rect -75 830 -25 850
rect 0 865 155 875
rect 0 845 10 865
rect 30 845 50 865
rect 70 845 90 865
rect 110 845 130 865
rect 0 835 155 845
rect 2735 870 2785 890
rect 2735 850 2750 870
rect 2770 850 2785 870
rect -75 810 -60 830
rect -40 810 -25 830
rect -75 790 -25 810
rect 175 823 2675 833
rect 175 803 200 823
rect 220 803 240 823
rect 260 803 280 823
rect 300 803 320 823
rect 340 803 360 823
rect 380 803 400 823
rect 420 803 440 823
rect 460 803 480 823
rect 500 803 520 823
rect 540 803 560 823
rect 580 803 600 823
rect 620 803 640 823
rect 660 803 680 823
rect 700 803 720 823
rect 740 803 760 823
rect 780 803 800 823
rect 820 803 840 823
rect 860 803 880 823
rect 900 803 920 823
rect 940 803 960 823
rect 980 803 1000 823
rect 1020 803 1040 823
rect 1060 803 1080 823
rect 1100 803 1120 823
rect 1140 803 1160 823
rect 1180 803 1200 823
rect 1220 803 1240 823
rect 1260 803 1280 823
rect 1300 803 1320 823
rect 1340 803 1360 823
rect 1380 803 1400 823
rect 1420 803 1440 823
rect 1460 803 1480 823
rect 1500 803 1520 823
rect 1540 803 1560 823
rect 1580 803 1600 823
rect 1620 803 1640 823
rect 1660 803 1680 823
rect 1700 803 1720 823
rect 1740 803 1760 823
rect 1780 803 1800 823
rect 1820 803 1840 823
rect 1860 803 1880 823
rect 1900 803 1920 823
rect 1940 803 1960 823
rect 1980 803 2000 823
rect 2020 803 2040 823
rect 2060 803 2080 823
rect 2100 803 2120 823
rect 2140 803 2160 823
rect 2180 803 2200 823
rect 2220 803 2240 823
rect 2260 803 2280 823
rect 2300 803 2320 823
rect 2340 803 2360 823
rect 2380 803 2400 823
rect 2420 803 2440 823
rect 2460 803 2480 823
rect 2500 803 2520 823
rect 2540 803 2560 823
rect 2580 803 2600 823
rect 2620 803 2640 823
rect 2660 803 2675 823
rect 175 793 2675 803
rect 2735 830 2785 850
rect 2735 810 2750 830
rect 2770 810 2785 830
rect 2735 790 2785 810
rect -75 770 -60 790
rect -40 770 -25 790
rect -75 750 -25 770
rect 0 780 155 790
rect 0 760 10 780
rect 30 760 50 780
rect 70 760 90 780
rect 110 760 130 780
rect 0 750 155 760
rect 2735 770 2750 790
rect 2770 770 2785 790
rect -75 730 -60 750
rect -40 730 -25 750
rect -75 710 -25 730
rect 175 741 2675 751
rect 175 721 200 741
rect 220 721 240 741
rect 260 721 280 741
rect 300 721 320 741
rect 340 721 360 741
rect 380 721 400 741
rect 420 721 440 741
rect 460 721 480 741
rect 500 721 520 741
rect 540 721 560 741
rect 580 721 600 741
rect 620 721 640 741
rect 660 721 680 741
rect 700 721 720 741
rect 740 721 760 741
rect 780 721 800 741
rect 820 721 840 741
rect 860 721 880 741
rect 900 721 920 741
rect 940 721 960 741
rect 980 721 1000 741
rect 1020 721 1040 741
rect 1060 721 1080 741
rect 1100 721 1120 741
rect 1140 721 1160 741
rect 1180 721 1200 741
rect 1220 721 1240 741
rect 1260 721 1280 741
rect 1300 721 1320 741
rect 1340 721 1360 741
rect 1380 721 1400 741
rect 1420 721 1440 741
rect 1460 721 1480 741
rect 1500 721 1520 741
rect 1540 721 1560 741
rect 1580 721 1600 741
rect 1620 721 1640 741
rect 1660 721 1680 741
rect 1700 721 1720 741
rect 1740 721 1760 741
rect 1780 721 1800 741
rect 1820 721 1840 741
rect 1860 721 1880 741
rect 1900 721 1920 741
rect 1940 721 1960 741
rect 1980 721 2000 741
rect 2020 721 2040 741
rect 2060 721 2080 741
rect 2100 721 2120 741
rect 2140 721 2160 741
rect 2180 721 2200 741
rect 2220 721 2240 741
rect 2260 721 2280 741
rect 2300 721 2320 741
rect 2340 721 2360 741
rect 2380 721 2400 741
rect 2420 721 2440 741
rect 2460 721 2480 741
rect 2500 721 2520 741
rect 2540 721 2560 741
rect 2580 721 2600 741
rect 2620 721 2640 741
rect 2660 721 2675 741
rect 175 711 2675 721
rect 2735 750 2785 770
rect 2735 730 2750 750
rect 2770 730 2785 750
rect 2735 710 2785 730
rect -75 690 -60 710
rect -40 690 -25 710
rect -75 670 -25 690
rect 0 700 155 710
rect 0 680 10 700
rect 30 680 50 700
rect 70 680 90 700
rect 110 680 130 700
rect 0 670 155 680
rect 2735 690 2750 710
rect 2770 690 2785 710
rect 2735 670 2785 690
rect -75 650 -60 670
rect -40 650 -25 670
rect -75 630 -25 650
rect 175 659 2675 669
rect 175 639 200 659
rect 220 639 240 659
rect 260 639 280 659
rect 300 639 320 659
rect 340 639 360 659
rect 380 639 400 659
rect 420 639 440 659
rect 460 639 480 659
rect 500 639 520 659
rect 540 639 560 659
rect 580 639 600 659
rect 620 639 640 659
rect 660 639 680 659
rect 700 639 720 659
rect 740 639 760 659
rect 780 639 800 659
rect 820 639 840 659
rect 860 639 880 659
rect 900 639 920 659
rect 940 639 960 659
rect 980 639 1000 659
rect 1020 639 1040 659
rect 1060 639 1080 659
rect 1100 639 1120 659
rect 1140 639 1160 659
rect 1180 639 1200 659
rect 1220 639 1240 659
rect 1260 639 1280 659
rect 1300 639 1320 659
rect 1340 639 1360 659
rect 1380 639 1400 659
rect 1420 639 1440 659
rect 1460 639 1480 659
rect 1500 639 1520 659
rect 1540 639 1560 659
rect 1580 639 1600 659
rect 1620 639 1640 659
rect 1660 639 1680 659
rect 1700 639 1720 659
rect 1740 639 1760 659
rect 1780 639 1800 659
rect 1820 639 1840 659
rect 1860 639 1880 659
rect 1900 639 1920 659
rect 1940 639 1960 659
rect 1980 639 2000 659
rect 2020 639 2040 659
rect 2060 639 2080 659
rect 2100 639 2120 659
rect 2140 639 2160 659
rect 2180 639 2200 659
rect 2220 639 2240 659
rect 2260 639 2280 659
rect 2300 639 2320 659
rect 2340 639 2360 659
rect 2380 639 2400 659
rect 2420 639 2440 659
rect 2460 639 2480 659
rect 2500 639 2520 659
rect 2540 639 2560 659
rect 2580 639 2600 659
rect 2620 639 2640 659
rect 2660 639 2675 659
rect -75 610 -60 630
rect -40 610 -25 630
rect -75 590 -25 610
rect 0 620 155 630
rect 175 629 2675 639
rect 2735 650 2750 670
rect 2770 650 2785 670
rect 2735 630 2785 650
rect 0 600 10 620
rect 30 600 50 620
rect 70 600 90 620
rect 110 600 130 620
rect 0 590 155 600
rect 2735 610 2750 630
rect 2770 610 2785 630
rect 2735 590 2785 610
rect -75 570 -60 590
rect -40 570 -25 590
rect -75 550 -25 570
rect -75 530 -60 550
rect -40 530 -25 550
rect 175 577 2675 587
rect 175 557 200 577
rect 220 557 240 577
rect 260 557 280 577
rect 300 557 320 577
rect 340 557 360 577
rect 380 557 400 577
rect 420 557 440 577
rect 460 557 480 577
rect 500 557 520 577
rect 540 557 560 577
rect 580 557 600 577
rect 620 557 640 577
rect 660 557 680 577
rect 700 557 720 577
rect 740 557 760 577
rect 780 557 800 577
rect 820 557 840 577
rect 860 557 880 577
rect 900 557 920 577
rect 940 557 960 577
rect 980 557 1000 577
rect 1020 557 1040 577
rect 1060 557 1080 577
rect 1100 557 1120 577
rect 1140 557 1160 577
rect 1180 557 1200 577
rect 1220 557 1240 577
rect 1260 557 1280 577
rect 1300 557 1320 577
rect 1340 557 1360 577
rect 1380 557 1400 577
rect 1420 557 1440 577
rect 1460 557 1480 577
rect 1500 557 1520 577
rect 1540 557 1560 577
rect 1580 557 1600 577
rect 1620 557 1640 577
rect 1660 557 1680 577
rect 1700 557 1720 577
rect 1740 557 1760 577
rect 1780 557 1800 577
rect 1820 557 1840 577
rect 1860 557 1880 577
rect 1900 557 1920 577
rect 1940 557 1960 577
rect 1980 557 2000 577
rect 2020 557 2040 577
rect 2060 557 2080 577
rect 2100 557 2120 577
rect 2140 557 2160 577
rect 2180 557 2200 577
rect 2220 557 2240 577
rect 2260 557 2280 577
rect 2300 557 2320 577
rect 2340 557 2360 577
rect 2380 557 2400 577
rect 2420 557 2440 577
rect 2460 557 2480 577
rect 2500 557 2520 577
rect 2540 557 2560 577
rect 2580 557 2600 577
rect 2620 557 2640 577
rect 2660 557 2675 577
rect 175 547 2675 557
rect 2735 570 2750 590
rect 2770 570 2785 590
rect 2735 550 2785 570
rect -75 510 -25 530
rect -75 490 -60 510
rect -40 490 -25 510
rect 0 535 155 545
rect 0 515 10 535
rect 30 515 50 535
rect 70 515 90 535
rect 110 515 130 535
rect 0 505 155 515
rect 2735 530 2750 550
rect 2770 530 2785 550
rect 2735 510 2785 530
rect -75 470 -25 490
rect -75 450 -60 470
rect -40 450 -25 470
rect 175 495 2675 505
rect 175 475 200 495
rect 220 475 240 495
rect 260 475 280 495
rect 300 475 320 495
rect 340 475 360 495
rect 380 475 400 495
rect 420 475 440 495
rect 460 475 480 495
rect 500 475 520 495
rect 540 475 560 495
rect 580 475 600 495
rect 620 475 640 495
rect 660 475 680 495
rect 700 475 720 495
rect 740 475 760 495
rect 780 475 800 495
rect 820 475 840 495
rect 860 475 880 495
rect 900 475 920 495
rect 940 475 960 495
rect 980 475 1000 495
rect 1020 475 1040 495
rect 1060 475 1080 495
rect 1100 475 1120 495
rect 1140 475 1160 495
rect 1180 475 1200 495
rect 1220 475 1240 495
rect 1260 475 1280 495
rect 1300 475 1320 495
rect 1340 475 1360 495
rect 1380 475 1400 495
rect 1420 475 1440 495
rect 1460 475 1480 495
rect 1500 475 1520 495
rect 1540 475 1560 495
rect 1580 475 1600 495
rect 1620 475 1640 495
rect 1660 475 1680 495
rect 1700 475 1720 495
rect 1740 475 1760 495
rect 1780 475 1800 495
rect 1820 475 1840 495
rect 1860 475 1880 495
rect 1900 475 1920 495
rect 1940 475 1960 495
rect 1980 475 2000 495
rect 2020 475 2040 495
rect 2060 475 2080 495
rect 2100 475 2120 495
rect 2140 475 2160 495
rect 2180 475 2200 495
rect 2220 475 2240 495
rect 2260 475 2280 495
rect 2300 475 2320 495
rect 2340 475 2360 495
rect 2380 475 2400 495
rect 2420 475 2440 495
rect 2460 475 2480 495
rect 2500 475 2520 495
rect 2540 475 2560 495
rect 2580 475 2600 495
rect 2620 475 2640 495
rect 2660 475 2675 495
rect 175 465 2675 475
rect 2735 490 2750 510
rect 2770 490 2785 510
rect 2735 470 2785 490
rect -75 430 -25 450
rect -75 410 -60 430
rect -40 410 -25 430
rect 0 455 155 465
rect 0 435 10 455
rect 30 435 50 455
rect 70 435 90 455
rect 110 435 130 455
rect 0 425 155 435
rect 2735 450 2750 470
rect 2770 450 2785 470
rect 2735 430 2785 450
rect -75 390 -25 410
rect -75 370 -60 390
rect -40 370 -25 390
rect 175 413 2675 423
rect 175 393 200 413
rect 220 393 240 413
rect 260 393 280 413
rect 300 393 320 413
rect 340 393 360 413
rect 380 393 400 413
rect 420 393 440 413
rect 460 393 480 413
rect 500 393 520 413
rect 540 393 560 413
rect 580 393 600 413
rect 620 393 640 413
rect 660 393 680 413
rect 700 393 720 413
rect 740 393 760 413
rect 780 393 800 413
rect 820 393 840 413
rect 860 393 880 413
rect 900 393 920 413
rect 940 393 960 413
rect 980 393 1000 413
rect 1020 393 1040 413
rect 1060 393 1080 413
rect 1100 393 1120 413
rect 1140 393 1160 413
rect 1180 393 1200 413
rect 1220 393 1240 413
rect 1260 393 1280 413
rect 1300 393 1320 413
rect 1340 393 1360 413
rect 1380 393 1400 413
rect 1420 393 1440 413
rect 1460 393 1480 413
rect 1500 393 1520 413
rect 1540 393 1560 413
rect 1580 393 1600 413
rect 1620 393 1640 413
rect 1660 393 1680 413
rect 1700 393 1720 413
rect 1740 393 1760 413
rect 1780 393 1800 413
rect 1820 393 1840 413
rect 1860 393 1880 413
rect 1900 393 1920 413
rect 1940 393 1960 413
rect 1980 393 2000 413
rect 2020 393 2040 413
rect 2060 393 2080 413
rect 2100 393 2120 413
rect 2140 393 2160 413
rect 2180 393 2200 413
rect 2220 393 2240 413
rect 2260 393 2280 413
rect 2300 393 2320 413
rect 2340 393 2360 413
rect 2380 393 2400 413
rect 2420 393 2440 413
rect 2460 393 2480 413
rect 2500 393 2520 413
rect 2540 393 2560 413
rect 2580 393 2600 413
rect 2620 393 2640 413
rect 2660 393 2675 413
rect -75 350 -25 370
rect -75 330 -60 350
rect -40 330 -25 350
rect 0 375 155 385
rect 175 383 2675 393
rect 2735 410 2750 430
rect 2770 410 2785 430
rect 2735 390 2785 410
rect 0 355 10 375
rect 30 355 50 375
rect 70 355 90 375
rect 110 355 130 375
rect 0 345 155 355
rect 2735 370 2750 390
rect 2770 370 2785 390
rect 2735 350 2785 370
rect -75 310 -25 330
rect -75 290 -60 310
rect -40 290 -25 310
rect 175 331 2675 341
rect 175 311 200 331
rect 220 311 240 331
rect 260 311 280 331
rect 300 311 320 331
rect 340 311 360 331
rect 380 311 400 331
rect 420 311 440 331
rect 460 311 480 331
rect 500 311 520 331
rect 540 311 560 331
rect 580 311 600 331
rect 620 311 640 331
rect 660 311 680 331
rect 700 311 720 331
rect 740 311 760 331
rect 780 311 800 331
rect 820 311 840 331
rect 860 311 880 331
rect 900 311 920 331
rect 940 311 960 331
rect 980 311 1000 331
rect 1020 311 1040 331
rect 1060 311 1080 331
rect 1100 311 1120 331
rect 1140 311 1160 331
rect 1180 311 1200 331
rect 1220 311 1240 331
rect 1260 311 1280 331
rect 1300 311 1320 331
rect 1340 311 1360 331
rect 1380 311 1400 331
rect 1420 311 1440 331
rect 1460 311 1480 331
rect 1500 311 1520 331
rect 1540 311 1560 331
rect 1580 311 1600 331
rect 1620 311 1640 331
rect 1660 311 1680 331
rect 1700 311 1720 331
rect 1740 311 1760 331
rect 1780 311 1800 331
rect 1820 311 1840 331
rect 1860 311 1880 331
rect 1900 311 1920 331
rect 1940 311 1960 331
rect 1980 311 2000 331
rect 2020 311 2040 331
rect 2060 311 2080 331
rect 2100 311 2120 331
rect 2140 311 2160 331
rect 2180 311 2200 331
rect 2220 311 2240 331
rect 2260 311 2280 331
rect 2300 311 2320 331
rect 2340 311 2360 331
rect 2380 311 2400 331
rect 2420 311 2440 331
rect 2460 311 2480 331
rect 2500 311 2520 331
rect 2540 311 2560 331
rect 2580 311 2600 331
rect 2620 311 2640 331
rect 2660 311 2675 331
rect 175 301 2675 311
rect 2735 330 2750 350
rect 2770 330 2785 350
rect 2735 310 2785 330
rect -75 270 -25 290
rect -75 250 -60 270
rect -40 250 -25 270
rect 0 290 155 300
rect 0 270 10 290
rect 30 270 50 290
rect 70 270 90 290
rect 110 270 130 290
rect 0 260 155 270
rect 2735 290 2750 310
rect 2770 290 2785 310
rect 2735 270 2785 290
rect -75 230 -25 250
rect -75 210 -60 230
rect -40 210 -25 230
rect 175 249 2675 259
rect 175 229 200 249
rect 220 229 240 249
rect 260 229 280 249
rect 300 229 320 249
rect 340 229 360 249
rect 380 229 400 249
rect 420 229 440 249
rect 460 229 480 249
rect 500 229 520 249
rect 540 229 560 249
rect 580 229 600 249
rect 620 229 640 249
rect 660 229 680 249
rect 700 229 720 249
rect 740 229 760 249
rect 780 229 800 249
rect 820 229 840 249
rect 860 229 880 249
rect 900 229 920 249
rect 940 229 960 249
rect 980 229 1000 249
rect 1020 229 1040 249
rect 1060 229 1080 249
rect 1100 229 1120 249
rect 1140 229 1160 249
rect 1180 229 1200 249
rect 1220 229 1240 249
rect 1260 229 1280 249
rect 1300 229 1320 249
rect 1340 229 1360 249
rect 1380 229 1400 249
rect 1420 229 1440 249
rect 1460 229 1480 249
rect 1500 229 1520 249
rect 1540 229 1560 249
rect 1580 229 1600 249
rect 1620 229 1640 249
rect 1660 229 1680 249
rect 1700 229 1720 249
rect 1740 229 1760 249
rect 1780 229 1800 249
rect 1820 229 1840 249
rect 1860 229 1880 249
rect 1900 229 1920 249
rect 1940 229 1960 249
rect 1980 229 2000 249
rect 2020 229 2040 249
rect 2060 229 2080 249
rect 2100 229 2120 249
rect 2140 229 2160 249
rect 2180 229 2200 249
rect 2220 229 2240 249
rect 2260 229 2280 249
rect 2300 229 2320 249
rect 2340 229 2360 249
rect 2380 229 2400 249
rect 2420 229 2440 249
rect 2460 229 2480 249
rect 2500 229 2520 249
rect 2540 229 2560 249
rect 2580 229 2600 249
rect 2620 229 2640 249
rect 2660 229 2675 249
rect -75 190 -25 210
rect -75 170 -60 190
rect -40 170 -25 190
rect 0 210 155 220
rect 175 219 2675 229
rect 2735 250 2750 270
rect 2770 250 2785 270
rect 2735 230 2785 250
rect 0 190 10 210
rect 30 190 50 210
rect 70 190 90 210
rect 110 190 130 210
rect 0 180 155 190
rect 2735 210 2750 230
rect 2770 210 2785 230
rect 2735 190 2785 210
rect -75 150 -25 170
rect -75 130 -60 150
rect -40 130 -25 150
rect 175 167 2675 177
rect 175 147 200 167
rect 220 147 240 167
rect 260 147 280 167
rect 300 147 320 167
rect 340 147 360 167
rect 380 147 400 167
rect 420 147 440 167
rect 460 147 480 167
rect 500 147 520 167
rect 540 147 560 167
rect 580 147 600 167
rect 620 147 640 167
rect 660 147 680 167
rect 700 147 720 167
rect 740 147 760 167
rect 780 147 800 167
rect 820 147 840 167
rect 860 147 880 167
rect 900 147 920 167
rect 940 147 960 167
rect 980 147 1000 167
rect 1020 147 1040 167
rect 1060 147 1080 167
rect 1100 147 1120 167
rect 1140 147 1160 167
rect 1180 147 1200 167
rect 1220 147 1240 167
rect 1260 147 1280 167
rect 1300 147 1320 167
rect 1340 147 1360 167
rect 1380 147 1400 167
rect 1420 147 1440 167
rect 1460 147 1480 167
rect 1500 147 1520 167
rect 1540 147 1560 167
rect 1580 147 1600 167
rect 1620 147 1640 167
rect 1660 147 1680 167
rect 1700 147 1720 167
rect 1740 147 1760 167
rect 1780 147 1800 167
rect 1820 147 1840 167
rect 1860 147 1880 167
rect 1900 147 1920 167
rect 1940 147 1960 167
rect 1980 147 2000 167
rect 2020 147 2040 167
rect 2060 147 2080 167
rect 2100 147 2120 167
rect 2140 147 2160 167
rect 2180 147 2200 167
rect 2220 147 2240 167
rect 2260 147 2280 167
rect 2300 147 2320 167
rect 2340 147 2360 167
rect 2380 147 2400 167
rect 2420 147 2440 167
rect 2460 147 2480 167
rect 2500 147 2520 167
rect 2540 147 2560 167
rect 2580 147 2600 167
rect 2620 147 2640 167
rect 2660 147 2675 167
rect -75 110 -25 130
rect -75 90 -60 110
rect -40 90 -25 110
rect 0 130 155 140
rect 175 137 2675 147
rect 2735 170 2750 190
rect 2770 170 2785 190
rect 2735 150 2785 170
rect 0 110 10 130
rect 30 110 50 130
rect 70 110 90 130
rect 110 110 130 130
rect 0 100 155 110
rect 2735 130 2750 150
rect 2770 130 2785 150
rect 2735 110 2785 130
rect -75 70 -25 90
rect -75 50 -60 70
rect -40 50 -25 70
rect -75 30 -25 50
rect -75 10 -60 30
rect -40 10 -25 30
rect 175 85 2675 95
rect 175 65 200 85
rect 220 65 240 85
rect 260 65 280 85
rect 300 65 320 85
rect 340 65 360 85
rect 380 65 400 85
rect 420 65 440 85
rect 460 65 480 85
rect 500 65 520 85
rect 540 65 560 85
rect 580 65 600 85
rect 620 65 640 85
rect 660 65 680 85
rect 700 65 720 85
rect 740 65 760 85
rect 780 65 800 85
rect 820 65 840 85
rect 860 65 880 85
rect 900 65 920 85
rect 940 65 960 85
rect 980 65 1000 85
rect 1020 65 1040 85
rect 1060 65 1080 85
rect 1100 65 1120 85
rect 1140 65 1160 85
rect 1180 65 1200 85
rect 1220 65 1240 85
rect 1260 65 1280 85
rect 1300 65 1320 85
rect 1340 65 1360 85
rect 1380 65 1400 85
rect 1420 65 1440 85
rect 1460 65 1480 85
rect 1500 65 1520 85
rect 1540 65 1560 85
rect 1580 65 1600 85
rect 1620 65 1640 85
rect 1660 65 1680 85
rect 1700 65 1720 85
rect 1740 65 1760 85
rect 1780 65 1800 85
rect 1820 65 1840 85
rect 1860 65 1880 85
rect 1900 65 1920 85
rect 1940 65 1960 85
rect 1980 65 2000 85
rect 2020 65 2040 85
rect 2060 65 2080 85
rect 2100 65 2120 85
rect 2140 65 2160 85
rect 2180 65 2200 85
rect 2220 65 2240 85
rect 2260 65 2280 85
rect 2300 65 2320 85
rect 2340 65 2360 85
rect 2380 65 2400 85
rect 2420 65 2440 85
rect 2460 65 2480 85
rect 2500 65 2520 85
rect 2540 65 2560 85
rect 2580 65 2600 85
rect 2620 65 2640 85
rect 2660 65 2675 85
rect 175 45 2675 65
rect 175 25 200 45
rect 220 25 240 45
rect 260 25 280 45
rect 300 25 320 45
rect 340 25 360 45
rect 380 25 400 45
rect 420 25 440 45
rect 460 25 480 45
rect 500 25 520 45
rect 540 25 560 45
rect 580 25 600 45
rect 620 25 640 45
rect 660 25 680 45
rect 700 25 720 45
rect 740 25 760 45
rect 780 25 800 45
rect 820 25 840 45
rect 860 25 880 45
rect 900 25 920 45
rect 940 25 960 45
rect 980 25 1000 45
rect 1020 25 1040 45
rect 1060 25 1080 45
rect 1100 25 1120 45
rect 1140 25 1160 45
rect 1180 25 1200 45
rect 1220 25 1240 45
rect 1260 25 1280 45
rect 1300 25 1320 45
rect 1340 25 1360 45
rect 1380 25 1400 45
rect 1420 25 1440 45
rect 1460 25 1480 45
rect 1500 25 1520 45
rect 1540 25 1560 45
rect 1580 25 1600 45
rect 1620 25 1640 45
rect 1660 25 1680 45
rect 1700 25 1720 45
rect 1740 25 1760 45
rect 1780 25 1800 45
rect 1820 25 1840 45
rect 1860 25 1880 45
rect 1900 25 1920 45
rect 1940 25 1960 45
rect 1980 25 2000 45
rect 2020 25 2040 45
rect 2060 25 2080 45
rect 2100 25 2120 45
rect 2140 25 2160 45
rect 2180 25 2200 45
rect 2220 25 2240 45
rect 2260 25 2280 45
rect 2300 25 2320 45
rect 2340 25 2360 45
rect 2380 25 2400 45
rect 2420 25 2440 45
rect 2460 25 2480 45
rect 2500 25 2520 45
rect 2540 25 2560 45
rect 2580 25 2600 45
rect 2620 25 2640 45
rect 2660 25 2675 45
rect 175 15 2675 25
rect 2735 90 2750 110
rect 2770 90 2785 110
rect 2735 70 2785 90
rect 2735 50 2750 70
rect 2770 50 2785 70
rect 2735 30 2785 50
rect -75 -10 -25 10
rect -75 -30 -60 -10
rect -40 -25 -25 -10
rect 2735 10 2750 30
rect 2770 10 2785 30
rect 2735 -10 2785 10
rect 2735 -25 2750 -10
rect -40 -30 2750 -25
rect 2770 -30 2785 -10
rect -75 -40 2785 -30
rect -75 -60 -20 -40
rect 0 -60 20 -40
rect 40 -60 60 -40
rect 80 -60 100 -40
rect 120 -60 140 -40
rect 160 -60 180 -40
rect 200 -60 220 -40
rect 240 -60 260 -40
rect 280 -60 300 -40
rect 320 -60 340 -40
rect 360 -60 380 -40
rect 400 -60 420 -40
rect 440 -60 460 -40
rect 480 -60 500 -40
rect 520 -60 540 -40
rect 560 -60 580 -40
rect 600 -60 620 -40
rect 640 -60 660 -40
rect 680 -60 700 -40
rect 720 -60 740 -40
rect 760 -60 780 -40
rect 800 -60 820 -40
rect 840 -60 860 -40
rect 880 -60 900 -40
rect 920 -60 940 -40
rect 960 -60 980 -40
rect 1000 -60 1020 -40
rect 1040 -60 1060 -40
rect 1080 -60 1100 -40
rect 1120 -60 1140 -40
rect 1160 -60 1180 -40
rect 1200 -60 1220 -40
rect 1240 -60 1260 -40
rect 1280 -60 1300 -40
rect 1320 -60 1340 -40
rect 1360 -60 1380 -40
rect 1400 -60 1420 -40
rect 1440 -60 1460 -40
rect 1480 -60 1500 -40
rect 1520 -60 1540 -40
rect 1560 -60 1580 -40
rect 1600 -60 1620 -40
rect 1640 -60 1660 -40
rect 1680 -60 1700 -40
rect 1720 -60 1740 -40
rect 1760 -60 1780 -40
rect 1800 -60 1820 -40
rect 1840 -60 1860 -40
rect 1880 -60 1900 -40
rect 1920 -60 1940 -40
rect 1960 -60 1980 -40
rect 2000 -60 2020 -40
rect 2040 -60 2060 -40
rect 2080 -60 2100 -40
rect 2120 -60 2140 -40
rect 2160 -60 2180 -40
rect 2200 -60 2220 -40
rect 2240 -60 2260 -40
rect 2280 -60 2300 -40
rect 2320 -60 2340 -40
rect 2360 -60 2380 -40
rect 2400 -60 2420 -40
rect 2440 -60 2460 -40
rect 2480 -60 2500 -40
rect 2520 -60 2540 -40
rect 2560 -60 2580 -40
rect 2600 -60 2620 -40
rect 2640 -60 2660 -40
rect 2680 -60 2700 -40
rect 2720 -60 2785 -40
rect -75 -75 2785 -60
rect 105 -175 2605 -165
rect 105 -195 120 -175
rect 140 -195 160 -175
rect 180 -195 200 -175
rect 220 -195 240 -175
rect 260 -195 280 -175
rect 300 -195 320 -175
rect 340 -195 360 -175
rect 380 -195 400 -175
rect 420 -195 440 -175
rect 460 -195 480 -175
rect 500 -195 520 -175
rect 540 -195 560 -175
rect 580 -195 600 -175
rect 620 -195 640 -175
rect 660 -195 680 -175
rect 700 -195 720 -175
rect 740 -195 760 -175
rect 780 -195 800 -175
rect 820 -195 840 -175
rect 860 -195 880 -175
rect 900 -195 920 -175
rect 940 -195 960 -175
rect 980 -195 1000 -175
rect 1020 -195 1040 -175
rect 1060 -195 1080 -175
rect 1100 -195 1120 -175
rect 1140 -195 1160 -175
rect 1180 -195 1200 -175
rect 1220 -195 1240 -175
rect 1260 -195 1280 -175
rect 1300 -195 1320 -175
rect 1340 -195 1360 -175
rect 1380 -195 1400 -175
rect 1420 -195 1440 -175
rect 1460 -195 1480 -175
rect 1500 -195 1520 -175
rect 1540 -195 1560 -175
rect 1580 -195 1600 -175
rect 1620 -195 1640 -175
rect 1660 -195 1680 -175
rect 1700 -195 1720 -175
rect 1740 -195 1760 -175
rect 1780 -195 1800 -175
rect 1820 -195 1840 -175
rect 1860 -195 1880 -175
rect 1900 -195 1920 -175
rect 1940 -195 1960 -175
rect 1980 -195 2000 -175
rect 2020 -195 2040 -175
rect 2060 -195 2080 -175
rect 2100 -195 2120 -175
rect 2140 -195 2160 -175
rect 2180 -195 2200 -175
rect 2220 -195 2240 -175
rect 2260 -195 2280 -175
rect 2300 -195 2320 -175
rect 2340 -195 2360 -175
rect 2380 -195 2400 -175
rect 2420 -195 2440 -175
rect 2460 -195 2480 -175
rect 2500 -195 2520 -175
rect 2540 -195 2560 -175
rect 2590 -195 2605 -175
rect 105 -215 2605 -195
rect 105 -235 120 -215
rect 140 -235 160 -215
rect 180 -235 200 -215
rect 220 -235 240 -215
rect 260 -235 280 -215
rect 300 -235 320 -215
rect 340 -235 360 -215
rect 380 -235 400 -215
rect 420 -235 440 -215
rect 460 -235 480 -215
rect 500 -235 520 -215
rect 540 -235 560 -215
rect 580 -235 600 -215
rect 620 -235 640 -215
rect 660 -235 680 -215
rect 700 -235 720 -215
rect 740 -235 760 -215
rect 780 -235 800 -215
rect 820 -235 840 -215
rect 860 -235 880 -215
rect 900 -235 920 -215
rect 940 -235 960 -215
rect 980 -235 1000 -215
rect 1020 -235 1040 -215
rect 1060 -235 1080 -215
rect 1100 -235 1120 -215
rect 1140 -235 1160 -215
rect 1180 -235 1200 -215
rect 1220 -235 1240 -215
rect 1260 -235 1280 -215
rect 1300 -235 1320 -215
rect 1340 -235 1360 -215
rect 1380 -235 1400 -215
rect 1420 -235 1440 -215
rect 1460 -235 1480 -215
rect 1500 -235 1520 -215
rect 1540 -235 1560 -215
rect 1580 -235 1600 -215
rect 1620 -235 1640 -215
rect 1660 -235 1680 -215
rect 1700 -235 1720 -215
rect 1740 -235 1760 -215
rect 1780 -235 1800 -215
rect 1820 -235 1840 -215
rect 1860 -235 1880 -215
rect 1900 -235 1920 -215
rect 1940 -235 1960 -215
rect 1980 -235 2000 -215
rect 2020 -235 2040 -215
rect 2060 -235 2080 -215
rect 2100 -235 2120 -215
rect 2140 -235 2160 -215
rect 2180 -235 2200 -215
rect 2220 -235 2240 -215
rect 2260 -235 2280 -215
rect 2300 -235 2320 -215
rect 2340 -235 2360 -215
rect 2380 -235 2400 -215
rect 2420 -235 2440 -215
rect 2460 -235 2480 -215
rect 2500 -235 2520 -215
rect 2540 -235 2560 -215
rect 2590 -235 2605 -215
rect 105 -245 2605 -235
rect -70 -260 85 -250
rect -70 -285 -60 -260
rect -40 -285 -20 -260
rect 0 -285 20 -260
rect 40 -285 60 -260
rect -70 -295 85 -285
rect 105 -310 2605 -300
rect 105 -330 120 -310
rect 140 -330 160 -310
rect 180 -330 200 -310
rect 220 -330 240 -310
rect 260 -330 280 -310
rect 300 -330 320 -310
rect 340 -330 360 -310
rect 380 -330 400 -310
rect 420 -330 440 -310
rect 460 -330 480 -310
rect 500 -330 520 -310
rect 540 -330 560 -310
rect 580 -330 600 -310
rect 620 -330 640 -310
rect 660 -330 680 -310
rect 700 -330 720 -310
rect 740 -330 760 -310
rect 780 -330 800 -310
rect 820 -330 840 -310
rect 860 -330 880 -310
rect 900 -330 920 -310
rect 940 -330 960 -310
rect 980 -330 1000 -310
rect 1020 -330 1040 -310
rect 1060 -330 1080 -310
rect 1100 -330 1120 -310
rect 1140 -330 1160 -310
rect 1180 -330 1200 -310
rect 1220 -330 1240 -310
rect 1260 -330 1280 -310
rect 1300 -330 1320 -310
rect 1340 -330 1360 -310
rect 1380 -330 1400 -310
rect 1420 -330 1440 -310
rect 1460 -330 1480 -310
rect 1500 -330 1520 -310
rect 1540 -330 1560 -310
rect 1580 -330 1600 -310
rect 1620 -330 1640 -310
rect 1660 -330 1680 -310
rect 1700 -330 1720 -310
rect 1740 -330 1760 -310
rect 1780 -330 1800 -310
rect 1820 -330 1840 -310
rect 1860 -330 1880 -310
rect 1900 -330 1920 -310
rect 1940 -330 1960 -310
rect 1980 -330 2000 -310
rect 2020 -330 2040 -310
rect 2060 -330 2080 -310
rect 2100 -330 2120 -310
rect 2140 -330 2160 -310
rect 2180 -330 2200 -310
rect 2220 -330 2240 -310
rect 2260 -330 2280 -310
rect 2300 -330 2320 -310
rect 2340 -330 2360 -310
rect 2380 -330 2400 -310
rect 2420 -330 2440 -310
rect 2460 -330 2480 -310
rect 2500 -330 2520 -310
rect 2540 -330 2560 -310
rect 2590 -330 2605 -310
rect 105 -340 2605 -330
rect -70 -355 85 -345
rect -70 -380 -60 -355
rect -40 -380 -20 -355
rect 0 -380 20 -355
rect 40 -380 60 -355
rect -70 -390 85 -380
rect 105 -405 2605 -395
rect 105 -425 120 -405
rect 140 -425 160 -405
rect 180 -425 200 -405
rect 220 -425 240 -405
rect 260 -425 280 -405
rect 300 -425 320 -405
rect 340 -425 360 -405
rect 380 -425 400 -405
rect 420 -425 440 -405
rect 460 -425 480 -405
rect 500 -425 520 -405
rect 540 -425 560 -405
rect 580 -425 600 -405
rect 620 -425 640 -405
rect 660 -425 680 -405
rect 700 -425 720 -405
rect 740 -425 760 -405
rect 780 -425 800 -405
rect 820 -425 840 -405
rect 860 -425 880 -405
rect 900 -425 920 -405
rect 940 -425 960 -405
rect 980 -425 1000 -405
rect 1020 -425 1040 -405
rect 1060 -425 1080 -405
rect 1100 -425 1120 -405
rect 1140 -425 1160 -405
rect 1180 -425 1200 -405
rect 1220 -425 1240 -405
rect 1260 -425 1280 -405
rect 1300 -425 1320 -405
rect 1340 -425 1360 -405
rect 1380 -425 1400 -405
rect 1420 -425 1440 -405
rect 1460 -425 1480 -405
rect 1500 -425 1520 -405
rect 1540 -425 1560 -405
rect 1580 -425 1600 -405
rect 1620 -425 1640 -405
rect 1660 -425 1680 -405
rect 1700 -425 1720 -405
rect 1740 -425 1760 -405
rect 1780 -425 1800 -405
rect 1820 -425 1840 -405
rect 1860 -425 1880 -405
rect 1900 -425 1920 -405
rect 1940 -425 1960 -405
rect 1980 -425 2000 -405
rect 2020 -425 2040 -405
rect 2060 -425 2080 -405
rect 2100 -425 2120 -405
rect 2140 -425 2160 -405
rect 2180 -425 2200 -405
rect 2220 -425 2240 -405
rect 2260 -425 2280 -405
rect 2300 -425 2320 -405
rect 2340 -425 2360 -405
rect 2380 -425 2400 -405
rect 2420 -425 2440 -405
rect 2460 -425 2480 -405
rect 2500 -425 2520 -405
rect 2540 -425 2560 -405
rect 2590 -425 2605 -405
rect 105 -435 2605 -425
rect -70 -450 85 -440
rect -70 -475 -60 -450
rect -40 -475 -20 -450
rect 0 -475 20 -450
rect 40 -475 60 -450
rect -70 -485 85 -475
rect 105 -500 2605 -490
rect 105 -520 120 -500
rect 140 -520 160 -500
rect 180 -520 200 -500
rect 220 -520 240 -500
rect 260 -520 280 -500
rect 300 -520 320 -500
rect 340 -520 360 -500
rect 380 -520 400 -500
rect 420 -520 440 -500
rect 460 -520 480 -500
rect 500 -520 520 -500
rect 540 -520 560 -500
rect 580 -520 600 -500
rect 620 -520 640 -500
rect 660 -520 680 -500
rect 700 -520 720 -500
rect 740 -520 760 -500
rect 780 -520 800 -500
rect 820 -520 840 -500
rect 860 -520 880 -500
rect 900 -520 920 -500
rect 940 -520 960 -500
rect 980 -520 1000 -500
rect 1020 -520 1040 -500
rect 1060 -520 1080 -500
rect 1100 -520 1120 -500
rect 1140 -520 1160 -500
rect 1180 -520 1200 -500
rect 1220 -520 1240 -500
rect 1260 -520 1280 -500
rect 1300 -520 1320 -500
rect 1340 -520 1360 -500
rect 1380 -520 1400 -500
rect 1420 -520 1440 -500
rect 1460 -520 1480 -500
rect 1500 -520 1520 -500
rect 1540 -520 1560 -500
rect 1580 -520 1600 -500
rect 1620 -520 1640 -500
rect 1660 -520 1680 -500
rect 1700 -520 1720 -500
rect 1740 -520 1760 -500
rect 1780 -520 1800 -500
rect 1820 -520 1840 -500
rect 1860 -520 1880 -500
rect 1900 -520 1920 -500
rect 1940 -520 1960 -500
rect 1980 -520 2000 -500
rect 2020 -520 2040 -500
rect 2060 -520 2080 -500
rect 2100 -520 2120 -500
rect 2140 -520 2160 -500
rect 2180 -520 2200 -500
rect 2220 -520 2240 -500
rect 2260 -520 2280 -500
rect 2300 -520 2320 -500
rect 2340 -520 2360 -500
rect 2380 -520 2400 -500
rect 2420 -520 2440 -500
rect 2460 -520 2480 -500
rect 2500 -520 2520 -500
rect 2540 -520 2560 -500
rect 2590 -520 2605 -500
rect 105 -530 2605 -520
rect -70 -545 85 -535
rect -70 -570 -60 -545
rect -40 -570 -20 -545
rect 0 -570 20 -545
rect 40 -570 60 -545
rect -70 -580 85 -570
rect 105 -595 2605 -585
rect 105 -615 120 -595
rect 140 -615 160 -595
rect 180 -615 200 -595
rect 220 -615 240 -595
rect 260 -615 280 -595
rect 300 -615 320 -595
rect 340 -615 360 -595
rect 380 -615 400 -595
rect 420 -615 440 -595
rect 460 -615 480 -595
rect 500 -615 520 -595
rect 540 -615 560 -595
rect 580 -615 600 -595
rect 620 -615 640 -595
rect 660 -615 680 -595
rect 700 -615 720 -595
rect 740 -615 760 -595
rect 780 -615 800 -595
rect 820 -615 840 -595
rect 860 -615 880 -595
rect 900 -615 920 -595
rect 940 -615 960 -595
rect 980 -615 1000 -595
rect 1020 -615 1040 -595
rect 1060 -615 1080 -595
rect 1100 -615 1120 -595
rect 1140 -615 1160 -595
rect 1180 -615 1200 -595
rect 1220 -615 1240 -595
rect 1260 -615 1280 -595
rect 1300 -615 1320 -595
rect 1340 -615 1360 -595
rect 1380 -615 1400 -595
rect 1420 -615 1440 -595
rect 1460 -615 1480 -595
rect 1500 -615 1520 -595
rect 1540 -615 1560 -595
rect 1580 -615 1600 -595
rect 1620 -615 1640 -595
rect 1660 -615 1680 -595
rect 1700 -615 1720 -595
rect 1740 -615 1760 -595
rect 1780 -615 1800 -595
rect 1820 -615 1840 -595
rect 1860 -615 1880 -595
rect 1900 -615 1920 -595
rect 1940 -615 1960 -595
rect 1980 -615 2000 -595
rect 2020 -615 2040 -595
rect 2060 -615 2080 -595
rect 2100 -615 2120 -595
rect 2140 -615 2160 -595
rect 2180 -615 2200 -595
rect 2220 -615 2240 -595
rect 2260 -615 2280 -595
rect 2300 -615 2320 -595
rect 2340 -615 2360 -595
rect 2380 -615 2400 -595
rect 2420 -615 2440 -595
rect 2460 -615 2480 -595
rect 2500 -615 2520 -595
rect 2540 -615 2560 -595
rect 2590 -615 2605 -595
rect 105 -625 2605 -615
rect -70 -640 85 -630
rect -70 -665 -60 -640
rect -40 -665 -20 -640
rect 0 -665 20 -640
rect 40 -665 60 -640
rect -70 -675 85 -665
rect 105 -690 2605 -680
rect 105 -710 120 -690
rect 140 -710 160 -690
rect 180 -710 200 -690
rect 220 -710 240 -690
rect 260 -710 280 -690
rect 300 -710 320 -690
rect 340 -710 360 -690
rect 380 -710 400 -690
rect 420 -710 440 -690
rect 460 -710 480 -690
rect 500 -710 520 -690
rect 540 -710 560 -690
rect 580 -710 600 -690
rect 620 -710 640 -690
rect 660 -710 680 -690
rect 700 -710 720 -690
rect 740 -710 760 -690
rect 780 -710 800 -690
rect 820 -710 840 -690
rect 860 -710 880 -690
rect 900 -710 920 -690
rect 940 -710 960 -690
rect 980 -710 1000 -690
rect 1020 -710 1040 -690
rect 1060 -710 1080 -690
rect 1100 -710 1120 -690
rect 1140 -710 1160 -690
rect 1180 -710 1200 -690
rect 1220 -710 1240 -690
rect 1260 -710 1280 -690
rect 1300 -710 1320 -690
rect 1340 -710 1360 -690
rect 1380 -710 1400 -690
rect 1420 -710 1440 -690
rect 1460 -710 1480 -690
rect 1500 -710 1520 -690
rect 1540 -710 1560 -690
rect 1580 -710 1600 -690
rect 1620 -710 1640 -690
rect 1660 -710 1680 -690
rect 1700 -710 1720 -690
rect 1740 -710 1760 -690
rect 1780 -710 1800 -690
rect 1820 -710 1840 -690
rect 1860 -710 1880 -690
rect 1900 -710 1920 -690
rect 1940 -710 1960 -690
rect 1980 -710 2000 -690
rect 2020 -710 2040 -690
rect 2060 -710 2080 -690
rect 2100 -710 2120 -690
rect 2140 -710 2160 -690
rect 2180 -710 2200 -690
rect 2220 -710 2240 -690
rect 2260 -710 2280 -690
rect 2300 -710 2320 -690
rect 2340 -710 2360 -690
rect 2380 -710 2400 -690
rect 2420 -710 2440 -690
rect 2460 -710 2480 -690
rect 2500 -710 2520 -690
rect 2540 -710 2560 -690
rect 2590 -710 2605 -690
rect 105 -720 2605 -710
rect -70 -735 85 -725
rect -70 -760 -60 -735
rect -40 -760 -20 -735
rect 0 -760 20 -735
rect 40 -760 60 -735
rect -70 -770 85 -760
rect 105 -785 2605 -775
rect 105 -805 120 -785
rect 140 -805 160 -785
rect 180 -805 200 -785
rect 220 -805 240 -785
rect 260 -805 280 -785
rect 300 -805 320 -785
rect 340 -805 360 -785
rect 380 -805 400 -785
rect 420 -805 440 -785
rect 460 -805 480 -785
rect 500 -805 520 -785
rect 540 -805 560 -785
rect 580 -805 600 -785
rect 620 -805 640 -785
rect 660 -805 680 -785
rect 700 -805 720 -785
rect 740 -805 760 -785
rect 780 -805 800 -785
rect 820 -805 840 -785
rect 860 -805 880 -785
rect 900 -805 920 -785
rect 940 -805 960 -785
rect 980 -805 1000 -785
rect 1020 -805 1040 -785
rect 1060 -805 1080 -785
rect 1100 -805 1120 -785
rect 1140 -805 1160 -785
rect 1180 -805 1200 -785
rect 1220 -805 1240 -785
rect 1260 -805 1280 -785
rect 1300 -805 1320 -785
rect 1340 -805 1360 -785
rect 1380 -805 1400 -785
rect 1420 -805 1440 -785
rect 1460 -805 1480 -785
rect 1500 -805 1520 -785
rect 1540 -805 1560 -785
rect 1580 -805 1600 -785
rect 1620 -805 1640 -785
rect 1660 -805 1680 -785
rect 1700 -805 1720 -785
rect 1740 -805 1760 -785
rect 1780 -805 1800 -785
rect 1820 -805 1840 -785
rect 1860 -805 1880 -785
rect 1900 -805 1920 -785
rect 1940 -805 1960 -785
rect 1980 -805 2000 -785
rect 2020 -805 2040 -785
rect 2060 -805 2080 -785
rect 2100 -805 2120 -785
rect 2140 -805 2160 -785
rect 2180 -805 2200 -785
rect 2220 -805 2240 -785
rect 2260 -805 2280 -785
rect 2300 -805 2320 -785
rect 2340 -805 2360 -785
rect 2380 -805 2400 -785
rect 2420 -805 2440 -785
rect 2460 -805 2480 -785
rect 2500 -805 2520 -785
rect 2540 -805 2560 -785
rect 2590 -805 2605 -785
rect 105 -815 2605 -805
rect -70 -830 85 -820
rect -70 -855 -60 -830
rect -40 -855 -20 -830
rect 0 -855 20 -830
rect 40 -855 60 -830
rect -70 -865 85 -855
rect 105 -880 2605 -870
rect 105 -900 120 -880
rect 140 -900 160 -880
rect 180 -900 200 -880
rect 220 -900 240 -880
rect 260 -900 280 -880
rect 300 -900 320 -880
rect 340 -900 360 -880
rect 380 -900 400 -880
rect 420 -900 440 -880
rect 460 -900 480 -880
rect 500 -900 520 -880
rect 540 -900 560 -880
rect 580 -900 600 -880
rect 620 -900 640 -880
rect 660 -900 680 -880
rect 700 -900 720 -880
rect 740 -900 760 -880
rect 780 -900 800 -880
rect 820 -900 840 -880
rect 860 -900 880 -880
rect 900 -900 920 -880
rect 940 -900 960 -880
rect 980 -900 1000 -880
rect 1020 -900 1040 -880
rect 1060 -900 1080 -880
rect 1100 -900 1120 -880
rect 1140 -900 1160 -880
rect 1180 -900 1200 -880
rect 1220 -900 1240 -880
rect 1260 -900 1280 -880
rect 1300 -900 1320 -880
rect 1340 -900 1360 -880
rect 1380 -900 1400 -880
rect 1420 -900 1440 -880
rect 1460 -900 1480 -880
rect 1500 -900 1520 -880
rect 1540 -900 1560 -880
rect 1580 -900 1600 -880
rect 1620 -900 1640 -880
rect 1660 -900 1680 -880
rect 1700 -900 1720 -880
rect 1740 -900 1760 -880
rect 1780 -900 1800 -880
rect 1820 -900 1840 -880
rect 1860 -900 1880 -880
rect 1900 -900 1920 -880
rect 1940 -900 1960 -880
rect 1980 -900 2000 -880
rect 2020 -900 2040 -880
rect 2060 -900 2080 -880
rect 2100 -900 2120 -880
rect 2140 -900 2160 -880
rect 2180 -900 2200 -880
rect 2220 -900 2240 -880
rect 2260 -900 2280 -880
rect 2300 -900 2320 -880
rect 2340 -900 2360 -880
rect 2380 -900 2400 -880
rect 2420 -900 2440 -880
rect 2460 -900 2480 -880
rect 2500 -900 2520 -880
rect 2540 -900 2560 -880
rect 2590 -900 2605 -880
rect 105 -910 2605 -900
rect -70 -925 85 -915
rect -70 -950 -60 -925
rect -40 -950 -20 -925
rect 0 -950 20 -925
rect 40 -950 60 -925
rect -70 -960 85 -950
rect 105 -975 2605 -965
rect 105 -995 120 -975
rect 140 -995 160 -975
rect 180 -995 200 -975
rect 220 -995 240 -975
rect 260 -995 280 -975
rect 300 -995 320 -975
rect 340 -995 360 -975
rect 380 -995 400 -975
rect 420 -995 440 -975
rect 460 -995 480 -975
rect 500 -995 520 -975
rect 540 -995 560 -975
rect 580 -995 600 -975
rect 620 -995 640 -975
rect 660 -995 680 -975
rect 700 -995 720 -975
rect 740 -995 760 -975
rect 780 -995 800 -975
rect 820 -995 840 -975
rect 860 -995 880 -975
rect 900 -995 920 -975
rect 940 -995 960 -975
rect 980 -995 1000 -975
rect 1020 -995 1040 -975
rect 1060 -995 1080 -975
rect 1100 -995 1120 -975
rect 1140 -995 1160 -975
rect 1180 -995 1200 -975
rect 1220 -995 1240 -975
rect 1260 -995 1280 -975
rect 1300 -995 1320 -975
rect 1340 -995 1360 -975
rect 1380 -995 1400 -975
rect 1420 -995 1440 -975
rect 1460 -995 1480 -975
rect 1500 -995 1520 -975
rect 1540 -995 1560 -975
rect 1580 -995 1600 -975
rect 1620 -995 1640 -975
rect 1660 -995 1680 -975
rect 1700 -995 1720 -975
rect 1740 -995 1760 -975
rect 1780 -995 1800 -975
rect 1820 -995 1840 -975
rect 1860 -995 1880 -975
rect 1900 -995 1920 -975
rect 1940 -995 1960 -975
rect 1980 -995 2000 -975
rect 2020 -995 2040 -975
rect 2060 -995 2080 -975
rect 2100 -995 2120 -975
rect 2140 -995 2160 -975
rect 2180 -995 2200 -975
rect 2220 -995 2240 -975
rect 2260 -995 2280 -975
rect 2300 -995 2320 -975
rect 2340 -995 2360 -975
rect 2380 -995 2400 -975
rect 2420 -995 2440 -975
rect 2460 -995 2480 -975
rect 2500 -995 2520 -975
rect 2540 -995 2560 -975
rect 2590 -995 2605 -975
rect 105 -1005 2605 -995
rect -70 -1020 85 -1010
rect -70 -1045 -60 -1020
rect -40 -1045 -20 -1020
rect 0 -1045 20 -1020
rect 40 -1045 60 -1020
rect -70 -1055 85 -1045
rect 105 -1070 2605 -1060
rect 105 -1090 120 -1070
rect 140 -1090 160 -1070
rect 180 -1090 200 -1070
rect 220 -1090 240 -1070
rect 260 -1090 280 -1070
rect 300 -1090 320 -1070
rect 340 -1090 360 -1070
rect 380 -1090 400 -1070
rect 420 -1090 440 -1070
rect 460 -1090 480 -1070
rect 500 -1090 520 -1070
rect 540 -1090 560 -1070
rect 580 -1090 600 -1070
rect 620 -1090 640 -1070
rect 660 -1090 680 -1070
rect 700 -1090 720 -1070
rect 740 -1090 760 -1070
rect 780 -1090 800 -1070
rect 820 -1090 840 -1070
rect 860 -1090 880 -1070
rect 900 -1090 920 -1070
rect 940 -1090 960 -1070
rect 980 -1090 1000 -1070
rect 1020 -1090 1040 -1070
rect 1060 -1090 1080 -1070
rect 1100 -1090 1120 -1070
rect 1140 -1090 1160 -1070
rect 1180 -1090 1200 -1070
rect 1220 -1090 1240 -1070
rect 1260 -1090 1280 -1070
rect 1300 -1090 1320 -1070
rect 1340 -1090 1360 -1070
rect 1380 -1090 1400 -1070
rect 1420 -1090 1440 -1070
rect 1460 -1090 1480 -1070
rect 1500 -1090 1520 -1070
rect 1540 -1090 1560 -1070
rect 1580 -1090 1600 -1070
rect 1620 -1090 1640 -1070
rect 1660 -1090 1680 -1070
rect 1700 -1090 1720 -1070
rect 1740 -1090 1760 -1070
rect 1780 -1090 1800 -1070
rect 1820 -1090 1840 -1070
rect 1860 -1090 1880 -1070
rect 1900 -1090 1920 -1070
rect 1940 -1090 1960 -1070
rect 1980 -1090 2000 -1070
rect 2020 -1090 2040 -1070
rect 2060 -1090 2080 -1070
rect 2100 -1090 2120 -1070
rect 2140 -1090 2160 -1070
rect 2180 -1090 2200 -1070
rect 2220 -1090 2240 -1070
rect 2260 -1090 2280 -1070
rect 2300 -1090 2320 -1070
rect 2340 -1090 2360 -1070
rect 2380 -1090 2400 -1070
rect 2420 -1090 2440 -1070
rect 2460 -1090 2480 -1070
rect 2500 -1090 2520 -1070
rect 2540 -1090 2560 -1070
rect 2590 -1090 2605 -1070
rect 105 -1100 2605 -1090
rect -70 -1115 85 -1105
rect -70 -1140 -60 -1115
rect -40 -1140 -20 -1115
rect 0 -1140 20 -1115
rect 40 -1140 60 -1115
rect -70 -1150 85 -1140
rect 105 -1165 2605 -1155
rect 105 -1185 120 -1165
rect 140 -1185 160 -1165
rect 180 -1185 200 -1165
rect 220 -1185 240 -1165
rect 260 -1185 280 -1165
rect 300 -1185 320 -1165
rect 340 -1185 360 -1165
rect 380 -1185 400 -1165
rect 420 -1185 440 -1165
rect 460 -1185 480 -1165
rect 500 -1185 520 -1165
rect 540 -1185 560 -1165
rect 580 -1185 600 -1165
rect 620 -1185 640 -1165
rect 660 -1185 680 -1165
rect 700 -1185 720 -1165
rect 740 -1185 760 -1165
rect 780 -1185 800 -1165
rect 820 -1185 840 -1165
rect 860 -1185 880 -1165
rect 900 -1185 920 -1165
rect 940 -1185 960 -1165
rect 980 -1185 1000 -1165
rect 1020 -1185 1040 -1165
rect 1060 -1185 1080 -1165
rect 1100 -1185 1120 -1165
rect 1140 -1185 1160 -1165
rect 1180 -1185 1200 -1165
rect 1220 -1185 1240 -1165
rect 1260 -1185 1280 -1165
rect 1300 -1185 1320 -1165
rect 1340 -1185 1360 -1165
rect 1380 -1185 1400 -1165
rect 1420 -1185 1440 -1165
rect 1460 -1185 1480 -1165
rect 1500 -1185 1520 -1165
rect 1540 -1185 1560 -1165
rect 1580 -1185 1600 -1165
rect 1620 -1185 1640 -1165
rect 1660 -1185 1680 -1165
rect 1700 -1185 1720 -1165
rect 1740 -1185 1760 -1165
rect 1780 -1185 1800 -1165
rect 1820 -1185 1840 -1165
rect 1860 -1185 1880 -1165
rect 1900 -1185 1920 -1165
rect 1940 -1185 1960 -1165
rect 1980 -1185 2000 -1165
rect 2020 -1185 2040 -1165
rect 2060 -1185 2080 -1165
rect 2100 -1185 2120 -1165
rect 2140 -1185 2160 -1165
rect 2180 -1185 2200 -1165
rect 2220 -1185 2240 -1165
rect 2260 -1185 2280 -1165
rect 2300 -1185 2320 -1165
rect 2340 -1185 2360 -1165
rect 2380 -1185 2400 -1165
rect 2420 -1185 2440 -1165
rect 2460 -1185 2480 -1165
rect 2500 -1185 2520 -1165
rect 2540 -1185 2560 -1165
rect 2590 -1185 2605 -1165
rect 105 -1195 2605 -1185
rect -70 -1210 85 -1200
rect -70 -1235 -60 -1210
rect -40 -1235 -20 -1210
rect 0 -1235 20 -1210
rect 40 -1235 60 -1210
rect -70 -1245 85 -1235
rect 105 -1260 2605 -1250
rect 105 -1280 120 -1260
rect 140 -1280 160 -1260
rect 180 -1280 200 -1260
rect 220 -1280 240 -1260
rect 260 -1280 280 -1260
rect 300 -1280 320 -1260
rect 340 -1280 360 -1260
rect 380 -1280 400 -1260
rect 420 -1280 440 -1260
rect 460 -1280 480 -1260
rect 500 -1280 520 -1260
rect 540 -1280 560 -1260
rect 580 -1280 600 -1260
rect 620 -1280 640 -1260
rect 660 -1280 680 -1260
rect 700 -1280 720 -1260
rect 740 -1280 760 -1260
rect 780 -1280 800 -1260
rect 820 -1280 840 -1260
rect 860 -1280 880 -1260
rect 900 -1280 920 -1260
rect 940 -1280 960 -1260
rect 980 -1280 1000 -1260
rect 1020 -1280 1040 -1260
rect 1060 -1280 1080 -1260
rect 1100 -1280 1120 -1260
rect 1140 -1280 1160 -1260
rect 1180 -1280 1200 -1260
rect 1220 -1280 1240 -1260
rect 1260 -1280 1280 -1260
rect 1300 -1280 1320 -1260
rect 1340 -1280 1360 -1260
rect 1380 -1280 1400 -1260
rect 1420 -1280 1440 -1260
rect 1460 -1280 1480 -1260
rect 1500 -1280 1520 -1260
rect 1540 -1280 1560 -1260
rect 1580 -1280 1600 -1260
rect 1620 -1280 1640 -1260
rect 1660 -1280 1680 -1260
rect 1700 -1280 1720 -1260
rect 1740 -1280 1760 -1260
rect 1780 -1280 1800 -1260
rect 1820 -1280 1840 -1260
rect 1860 -1280 1880 -1260
rect 1900 -1280 1920 -1260
rect 1940 -1280 1960 -1260
rect 1980 -1280 2000 -1260
rect 2020 -1280 2040 -1260
rect 2060 -1280 2080 -1260
rect 2100 -1280 2120 -1260
rect 2140 -1280 2160 -1260
rect 2180 -1280 2200 -1260
rect 2220 -1280 2240 -1260
rect 2260 -1280 2280 -1260
rect 2300 -1280 2320 -1260
rect 2340 -1280 2360 -1260
rect 2380 -1280 2400 -1260
rect 2420 -1280 2440 -1260
rect 2460 -1280 2480 -1260
rect 2500 -1280 2520 -1260
rect 2540 -1280 2560 -1260
rect 2590 -1280 2605 -1260
rect 105 -1290 2605 -1280
rect -70 -1305 85 -1295
rect -70 -1330 -60 -1305
rect -40 -1330 -20 -1305
rect 0 -1330 20 -1305
rect 40 -1330 60 -1305
rect -70 -1340 85 -1330
rect 105 -1355 2605 -1345
rect 105 -1375 120 -1355
rect 140 -1375 160 -1355
rect 180 -1375 200 -1355
rect 220 -1375 240 -1355
rect 260 -1375 280 -1355
rect 300 -1375 320 -1355
rect 340 -1375 360 -1355
rect 380 -1375 400 -1355
rect 420 -1375 440 -1355
rect 460 -1375 480 -1355
rect 500 -1375 520 -1355
rect 540 -1375 560 -1355
rect 580 -1375 600 -1355
rect 620 -1375 640 -1355
rect 660 -1375 680 -1355
rect 700 -1375 720 -1355
rect 740 -1375 760 -1355
rect 780 -1375 800 -1355
rect 820 -1375 840 -1355
rect 860 -1375 880 -1355
rect 900 -1375 920 -1355
rect 940 -1375 960 -1355
rect 980 -1375 1000 -1355
rect 1020 -1375 1040 -1355
rect 1060 -1375 1080 -1355
rect 1100 -1375 1120 -1355
rect 1140 -1375 1160 -1355
rect 1180 -1375 1200 -1355
rect 1220 -1375 1240 -1355
rect 1260 -1375 1280 -1355
rect 1300 -1375 1320 -1355
rect 1340 -1375 1360 -1355
rect 1380 -1375 1400 -1355
rect 1420 -1375 1440 -1355
rect 1460 -1375 1480 -1355
rect 1500 -1375 1520 -1355
rect 1540 -1375 1560 -1355
rect 1580 -1375 1600 -1355
rect 1620 -1375 1640 -1355
rect 1660 -1375 1680 -1355
rect 1700 -1375 1720 -1355
rect 1740 -1375 1760 -1355
rect 1780 -1375 1800 -1355
rect 1820 -1375 1840 -1355
rect 1860 -1375 1880 -1355
rect 1900 -1375 1920 -1355
rect 1940 -1375 1960 -1355
rect 1980 -1375 2000 -1355
rect 2020 -1375 2040 -1355
rect 2060 -1375 2080 -1355
rect 2100 -1375 2120 -1355
rect 2140 -1375 2160 -1355
rect 2180 -1375 2200 -1355
rect 2220 -1375 2240 -1355
rect 2260 -1375 2280 -1355
rect 2300 -1375 2320 -1355
rect 2340 -1375 2360 -1355
rect 2380 -1375 2400 -1355
rect 2420 -1375 2440 -1355
rect 2460 -1375 2480 -1355
rect 2500 -1375 2520 -1355
rect 2540 -1375 2560 -1355
rect 2590 -1375 2605 -1355
rect 105 -1385 2605 -1375
rect -70 -1400 85 -1390
rect -70 -1425 -60 -1400
rect -40 -1425 -20 -1400
rect 0 -1425 20 -1400
rect 40 -1425 60 -1400
rect -70 -1435 85 -1425
rect 105 -1450 2605 -1440
rect 105 -1470 120 -1450
rect 140 -1470 160 -1450
rect 180 -1470 200 -1450
rect 220 -1470 240 -1450
rect 260 -1470 280 -1450
rect 300 -1470 320 -1450
rect 340 -1470 360 -1450
rect 380 -1470 400 -1450
rect 420 -1470 440 -1450
rect 460 -1470 480 -1450
rect 500 -1470 520 -1450
rect 540 -1470 560 -1450
rect 580 -1470 600 -1450
rect 620 -1470 640 -1450
rect 660 -1470 680 -1450
rect 700 -1470 720 -1450
rect 740 -1470 760 -1450
rect 780 -1470 800 -1450
rect 820 -1470 840 -1450
rect 860 -1470 880 -1450
rect 900 -1470 920 -1450
rect 940 -1470 960 -1450
rect 980 -1470 1000 -1450
rect 1020 -1470 1040 -1450
rect 1060 -1470 1080 -1450
rect 1100 -1470 1120 -1450
rect 1140 -1470 1160 -1450
rect 1180 -1470 1200 -1450
rect 1220 -1470 1240 -1450
rect 1260 -1470 1280 -1450
rect 1300 -1470 1320 -1450
rect 1340 -1470 1360 -1450
rect 1380 -1470 1400 -1450
rect 1420 -1470 1440 -1450
rect 1460 -1470 1480 -1450
rect 1500 -1470 1520 -1450
rect 1540 -1470 1560 -1450
rect 1580 -1470 1600 -1450
rect 1620 -1470 1640 -1450
rect 1660 -1470 1680 -1450
rect 1700 -1470 1720 -1450
rect 1740 -1470 1760 -1450
rect 1780 -1470 1800 -1450
rect 1820 -1470 1840 -1450
rect 1860 -1470 1880 -1450
rect 1900 -1470 1920 -1450
rect 1940 -1470 1960 -1450
rect 1980 -1470 2000 -1450
rect 2020 -1470 2040 -1450
rect 2060 -1470 2080 -1450
rect 2100 -1470 2120 -1450
rect 2140 -1470 2160 -1450
rect 2180 -1470 2200 -1450
rect 2220 -1470 2240 -1450
rect 2260 -1470 2280 -1450
rect 2300 -1470 2320 -1450
rect 2340 -1470 2360 -1450
rect 2380 -1470 2400 -1450
rect 2420 -1470 2440 -1450
rect 2460 -1470 2480 -1450
rect 2500 -1470 2520 -1450
rect 2540 -1470 2560 -1450
rect 2590 -1470 2605 -1450
rect 105 -1480 2605 -1470
rect -70 -1495 85 -1485
rect -70 -1520 -60 -1495
rect -40 -1520 -20 -1495
rect 0 -1520 20 -1495
rect 40 -1520 60 -1495
rect -70 -1530 85 -1520
rect 105 -1545 2605 -1535
rect 105 -1565 120 -1545
rect 140 -1565 160 -1545
rect 180 -1565 200 -1545
rect 220 -1565 240 -1545
rect 260 -1565 280 -1545
rect 300 -1565 320 -1545
rect 340 -1565 360 -1545
rect 380 -1565 400 -1545
rect 420 -1565 440 -1545
rect 460 -1565 480 -1545
rect 500 -1565 520 -1545
rect 540 -1565 560 -1545
rect 580 -1565 600 -1545
rect 620 -1565 640 -1545
rect 660 -1565 680 -1545
rect 700 -1565 720 -1545
rect 740 -1565 760 -1545
rect 780 -1565 800 -1545
rect 820 -1565 840 -1545
rect 860 -1565 880 -1545
rect 900 -1565 920 -1545
rect 940 -1565 960 -1545
rect 980 -1565 1000 -1545
rect 1020 -1565 1040 -1545
rect 1060 -1565 1080 -1545
rect 1100 -1565 1120 -1545
rect 1140 -1565 1160 -1545
rect 1180 -1565 1200 -1545
rect 1220 -1565 1240 -1545
rect 1260 -1565 1280 -1545
rect 1300 -1565 1320 -1545
rect 1340 -1565 1360 -1545
rect 1380 -1565 1400 -1545
rect 1420 -1565 1440 -1545
rect 1460 -1565 1480 -1545
rect 1500 -1565 1520 -1545
rect 1540 -1565 1560 -1545
rect 1580 -1565 1600 -1545
rect 1620 -1565 1640 -1545
rect 1660 -1565 1680 -1545
rect 1700 -1565 1720 -1545
rect 1740 -1565 1760 -1545
rect 1780 -1565 1800 -1545
rect 1820 -1565 1840 -1545
rect 1860 -1565 1880 -1545
rect 1900 -1565 1920 -1545
rect 1940 -1565 1960 -1545
rect 1980 -1565 2000 -1545
rect 2020 -1565 2040 -1545
rect 2060 -1565 2080 -1545
rect 2100 -1565 2120 -1545
rect 2140 -1565 2160 -1545
rect 2180 -1565 2200 -1545
rect 2220 -1565 2240 -1545
rect 2260 -1565 2280 -1545
rect 2300 -1565 2320 -1545
rect 2340 -1565 2360 -1545
rect 2380 -1565 2400 -1545
rect 2420 -1565 2440 -1545
rect 2460 -1565 2480 -1545
rect 2500 -1565 2520 -1545
rect 2540 -1565 2560 -1545
rect 2590 -1565 2605 -1545
rect 105 -1575 2605 -1565
rect -70 -1590 85 -1580
rect -70 -1615 -60 -1590
rect -40 -1615 -20 -1590
rect 0 -1615 20 -1590
rect 40 -1615 60 -1590
rect -70 -1625 85 -1615
rect 105 -1640 2605 -1630
rect 105 -1660 120 -1640
rect 140 -1660 160 -1640
rect 180 -1660 200 -1640
rect 220 -1660 240 -1640
rect 260 -1660 280 -1640
rect 300 -1660 320 -1640
rect 340 -1660 360 -1640
rect 380 -1660 400 -1640
rect 420 -1660 440 -1640
rect 460 -1660 480 -1640
rect 500 -1660 520 -1640
rect 540 -1660 560 -1640
rect 580 -1660 600 -1640
rect 620 -1660 640 -1640
rect 660 -1660 680 -1640
rect 700 -1660 720 -1640
rect 740 -1660 760 -1640
rect 780 -1660 800 -1640
rect 820 -1660 840 -1640
rect 860 -1660 880 -1640
rect 900 -1660 920 -1640
rect 940 -1660 960 -1640
rect 980 -1660 1000 -1640
rect 1020 -1660 1040 -1640
rect 1060 -1660 1080 -1640
rect 1100 -1660 1120 -1640
rect 1140 -1660 1160 -1640
rect 1180 -1660 1200 -1640
rect 1220 -1660 1240 -1640
rect 1260 -1660 1280 -1640
rect 1300 -1660 1320 -1640
rect 1340 -1660 1360 -1640
rect 1380 -1660 1400 -1640
rect 1420 -1660 1440 -1640
rect 1460 -1660 1480 -1640
rect 1500 -1660 1520 -1640
rect 1540 -1660 1560 -1640
rect 1580 -1660 1600 -1640
rect 1620 -1660 1640 -1640
rect 1660 -1660 1680 -1640
rect 1700 -1660 1720 -1640
rect 1740 -1660 1760 -1640
rect 1780 -1660 1800 -1640
rect 1820 -1660 1840 -1640
rect 1860 -1660 1880 -1640
rect 1900 -1660 1920 -1640
rect 1940 -1660 1960 -1640
rect 1980 -1660 2000 -1640
rect 2020 -1660 2040 -1640
rect 2060 -1660 2080 -1640
rect 2100 -1660 2120 -1640
rect 2140 -1660 2160 -1640
rect 2180 -1660 2200 -1640
rect 2220 -1660 2240 -1640
rect 2260 -1660 2280 -1640
rect 2300 -1660 2320 -1640
rect 2340 -1660 2360 -1640
rect 2380 -1660 2400 -1640
rect 2420 -1660 2440 -1640
rect 2460 -1660 2480 -1640
rect 2500 -1660 2520 -1640
rect 2540 -1660 2560 -1640
rect 2590 -1660 2605 -1640
rect 105 -1670 2605 -1660
rect -70 -1685 85 -1675
rect -70 -1710 -60 -1685
rect -40 -1710 -20 -1685
rect 0 -1710 20 -1685
rect 40 -1710 60 -1685
rect -70 -1720 85 -1710
rect 105 -1735 2605 -1725
rect 105 -1755 120 -1735
rect 140 -1755 160 -1735
rect 180 -1755 200 -1735
rect 220 -1755 240 -1735
rect 260 -1755 280 -1735
rect 300 -1755 320 -1735
rect 340 -1755 360 -1735
rect 380 -1755 400 -1735
rect 420 -1755 440 -1735
rect 460 -1755 480 -1735
rect 500 -1755 520 -1735
rect 540 -1755 560 -1735
rect 580 -1755 600 -1735
rect 620 -1755 640 -1735
rect 660 -1755 680 -1735
rect 700 -1755 720 -1735
rect 740 -1755 760 -1735
rect 780 -1755 800 -1735
rect 820 -1755 840 -1735
rect 860 -1755 880 -1735
rect 900 -1755 920 -1735
rect 940 -1755 960 -1735
rect 980 -1755 1000 -1735
rect 1020 -1755 1040 -1735
rect 1060 -1755 1080 -1735
rect 1100 -1755 1120 -1735
rect 1140 -1755 1160 -1735
rect 1180 -1755 1200 -1735
rect 1220 -1755 1240 -1735
rect 1260 -1755 1280 -1735
rect 1300 -1755 1320 -1735
rect 1340 -1755 1360 -1735
rect 1380 -1755 1400 -1735
rect 1420 -1755 1440 -1735
rect 1460 -1755 1480 -1735
rect 1500 -1755 1520 -1735
rect 1540 -1755 1560 -1735
rect 1580 -1755 1600 -1735
rect 1620 -1755 1640 -1735
rect 1660 -1755 1680 -1735
rect 1700 -1755 1720 -1735
rect 1740 -1755 1760 -1735
rect 1780 -1755 1800 -1735
rect 1820 -1755 1840 -1735
rect 1860 -1755 1880 -1735
rect 1900 -1755 1920 -1735
rect 1940 -1755 1960 -1735
rect 1980 -1755 2000 -1735
rect 2020 -1755 2040 -1735
rect 2060 -1755 2080 -1735
rect 2100 -1755 2120 -1735
rect 2140 -1755 2160 -1735
rect 2180 -1755 2200 -1735
rect 2220 -1755 2240 -1735
rect 2260 -1755 2280 -1735
rect 2300 -1755 2320 -1735
rect 2340 -1755 2360 -1735
rect 2380 -1755 2400 -1735
rect 2420 -1755 2440 -1735
rect 2460 -1755 2480 -1735
rect 2500 -1755 2520 -1735
rect 2540 -1755 2560 -1735
rect 2590 -1755 2605 -1735
rect 105 -1765 2605 -1755
rect -70 -1780 85 -1770
rect -70 -1805 -60 -1780
rect -40 -1805 -20 -1780
rect 0 -1805 20 -1780
rect 40 -1805 60 -1780
rect -70 -1815 85 -1805
rect 105 -1830 2605 -1820
rect 105 -1850 120 -1830
rect 140 -1850 160 -1830
rect 180 -1850 200 -1830
rect 220 -1850 240 -1830
rect 260 -1850 280 -1830
rect 300 -1850 320 -1830
rect 340 -1850 360 -1830
rect 380 -1850 400 -1830
rect 420 -1850 440 -1830
rect 460 -1850 480 -1830
rect 500 -1850 520 -1830
rect 540 -1850 560 -1830
rect 580 -1850 600 -1830
rect 620 -1850 640 -1830
rect 660 -1850 680 -1830
rect 700 -1850 720 -1830
rect 740 -1850 760 -1830
rect 780 -1850 800 -1830
rect 820 -1850 840 -1830
rect 860 -1850 880 -1830
rect 900 -1850 920 -1830
rect 940 -1850 960 -1830
rect 980 -1850 1000 -1830
rect 1020 -1850 1040 -1830
rect 1060 -1850 1080 -1830
rect 1100 -1850 1120 -1830
rect 1140 -1850 1160 -1830
rect 1180 -1850 1200 -1830
rect 1220 -1850 1240 -1830
rect 1260 -1850 1280 -1830
rect 1300 -1850 1320 -1830
rect 1340 -1850 1360 -1830
rect 1380 -1850 1400 -1830
rect 1420 -1850 1440 -1830
rect 1460 -1850 1480 -1830
rect 1500 -1850 1520 -1830
rect 1540 -1850 1560 -1830
rect 1580 -1850 1600 -1830
rect 1620 -1850 1640 -1830
rect 1660 -1850 1680 -1830
rect 1700 -1850 1720 -1830
rect 1740 -1850 1760 -1830
rect 1780 -1850 1800 -1830
rect 1820 -1850 1840 -1830
rect 1860 -1850 1880 -1830
rect 1900 -1850 1920 -1830
rect 1940 -1850 1960 -1830
rect 1980 -1850 2000 -1830
rect 2020 -1850 2040 -1830
rect 2060 -1850 2080 -1830
rect 2100 -1850 2120 -1830
rect 2140 -1850 2160 -1830
rect 2180 -1850 2200 -1830
rect 2220 -1850 2240 -1830
rect 2260 -1850 2280 -1830
rect 2300 -1850 2320 -1830
rect 2340 -1850 2360 -1830
rect 2380 -1850 2400 -1830
rect 2420 -1850 2440 -1830
rect 2460 -1850 2480 -1830
rect 2500 -1850 2520 -1830
rect 2540 -1850 2560 -1830
rect 2590 -1850 2605 -1830
rect 105 -1860 2605 -1850
rect -70 -1875 85 -1865
rect -70 -1900 -60 -1875
rect -40 -1900 -20 -1875
rect 0 -1900 20 -1875
rect 40 -1900 60 -1875
rect -70 -1910 85 -1900
rect 105 -1925 2605 -1915
rect 105 -1945 120 -1925
rect 140 -1945 160 -1925
rect 180 -1945 200 -1925
rect 220 -1945 240 -1925
rect 260 -1945 280 -1925
rect 300 -1945 320 -1925
rect 340 -1945 360 -1925
rect 380 -1945 400 -1925
rect 420 -1945 440 -1925
rect 460 -1945 480 -1925
rect 500 -1945 520 -1925
rect 540 -1945 560 -1925
rect 580 -1945 600 -1925
rect 620 -1945 640 -1925
rect 660 -1945 680 -1925
rect 700 -1945 720 -1925
rect 740 -1945 760 -1925
rect 780 -1945 800 -1925
rect 820 -1945 840 -1925
rect 860 -1945 880 -1925
rect 900 -1945 920 -1925
rect 940 -1945 960 -1925
rect 980 -1945 1000 -1925
rect 1020 -1945 1040 -1925
rect 1060 -1945 1080 -1925
rect 1100 -1945 1120 -1925
rect 1140 -1945 1160 -1925
rect 1180 -1945 1200 -1925
rect 1220 -1945 1240 -1925
rect 1260 -1945 1280 -1925
rect 1300 -1945 1320 -1925
rect 1340 -1945 1360 -1925
rect 1380 -1945 1400 -1925
rect 1420 -1945 1440 -1925
rect 1460 -1945 1480 -1925
rect 1500 -1945 1520 -1925
rect 1540 -1945 1560 -1925
rect 1580 -1945 1600 -1925
rect 1620 -1945 1640 -1925
rect 1660 -1945 1680 -1925
rect 1700 -1945 1720 -1925
rect 1740 -1945 1760 -1925
rect 1780 -1945 1800 -1925
rect 1820 -1945 1840 -1925
rect 1860 -1945 1880 -1925
rect 1900 -1945 1920 -1925
rect 1940 -1945 1960 -1925
rect 1980 -1945 2000 -1925
rect 2020 -1945 2040 -1925
rect 2060 -1945 2080 -1925
rect 2100 -1945 2120 -1925
rect 2140 -1945 2160 -1925
rect 2180 -1945 2200 -1925
rect 2220 -1945 2240 -1925
rect 2260 -1945 2280 -1925
rect 2300 -1945 2320 -1925
rect 2340 -1945 2360 -1925
rect 2380 -1945 2400 -1925
rect 2420 -1945 2440 -1925
rect 2460 -1945 2480 -1925
rect 2500 -1945 2520 -1925
rect 2540 -1945 2560 -1925
rect 2590 -1945 2605 -1925
rect 105 -1955 2605 -1945
rect -70 -1970 85 -1960
rect -70 -1995 -60 -1970
rect -40 -1995 -20 -1970
rect 0 -1995 20 -1970
rect 40 -1995 60 -1970
rect -70 -2005 85 -1995
rect 105 -2020 2605 -2010
rect 105 -2040 120 -2020
rect 140 -2040 160 -2020
rect 180 -2040 200 -2020
rect 220 -2040 240 -2020
rect 260 -2040 280 -2020
rect 300 -2040 320 -2020
rect 340 -2040 360 -2020
rect 380 -2040 400 -2020
rect 420 -2040 440 -2020
rect 460 -2040 480 -2020
rect 500 -2040 520 -2020
rect 540 -2040 560 -2020
rect 580 -2040 600 -2020
rect 620 -2040 640 -2020
rect 660 -2040 680 -2020
rect 700 -2040 720 -2020
rect 740 -2040 760 -2020
rect 780 -2040 800 -2020
rect 820 -2040 840 -2020
rect 860 -2040 880 -2020
rect 900 -2040 920 -2020
rect 940 -2040 960 -2020
rect 980 -2040 1000 -2020
rect 1020 -2040 1040 -2020
rect 1060 -2040 1080 -2020
rect 1100 -2040 1120 -2020
rect 1140 -2040 1160 -2020
rect 1180 -2040 1200 -2020
rect 1220 -2040 1240 -2020
rect 1260 -2040 1280 -2020
rect 1300 -2040 1320 -2020
rect 1340 -2040 1360 -2020
rect 1380 -2040 1400 -2020
rect 1420 -2040 1440 -2020
rect 1460 -2040 1480 -2020
rect 1500 -2040 1520 -2020
rect 1540 -2040 1560 -2020
rect 1580 -2040 1600 -2020
rect 1620 -2040 1640 -2020
rect 1660 -2040 1680 -2020
rect 1700 -2040 1720 -2020
rect 1740 -2040 1760 -2020
rect 1780 -2040 1800 -2020
rect 1820 -2040 1840 -2020
rect 1860 -2040 1880 -2020
rect 1900 -2040 1920 -2020
rect 1940 -2040 1960 -2020
rect 1980 -2040 2000 -2020
rect 2020 -2040 2040 -2020
rect 2060 -2040 2080 -2020
rect 2100 -2040 2120 -2020
rect 2140 -2040 2160 -2020
rect 2180 -2040 2200 -2020
rect 2220 -2040 2240 -2020
rect 2260 -2040 2280 -2020
rect 2300 -2040 2320 -2020
rect 2340 -2040 2360 -2020
rect 2380 -2040 2400 -2020
rect 2420 -2040 2440 -2020
rect 2460 -2040 2480 -2020
rect 2500 -2040 2520 -2020
rect 2540 -2040 2560 -2020
rect 2590 -2040 2605 -2020
rect 105 -2050 2605 -2040
rect -70 -2065 85 -2055
rect -70 -2090 -60 -2065
rect -40 -2090 -20 -2065
rect 0 -2090 20 -2065
rect 40 -2090 60 -2065
rect -70 -2100 85 -2090
rect 105 -2115 2605 -2105
rect 105 -2135 120 -2115
rect 140 -2135 160 -2115
rect 180 -2135 200 -2115
rect 220 -2135 240 -2115
rect 260 -2135 280 -2115
rect 300 -2135 320 -2115
rect 340 -2135 360 -2115
rect 380 -2135 400 -2115
rect 420 -2135 440 -2115
rect 460 -2135 480 -2115
rect 500 -2135 520 -2115
rect 540 -2135 560 -2115
rect 580 -2135 600 -2115
rect 620 -2135 640 -2115
rect 660 -2135 680 -2115
rect 700 -2135 720 -2115
rect 740 -2135 760 -2115
rect 780 -2135 800 -2115
rect 820 -2135 840 -2115
rect 860 -2135 880 -2115
rect 900 -2135 920 -2115
rect 940 -2135 960 -2115
rect 980 -2135 1000 -2115
rect 1020 -2135 1040 -2115
rect 1060 -2135 1080 -2115
rect 1100 -2135 1120 -2115
rect 1140 -2135 1160 -2115
rect 1180 -2135 1200 -2115
rect 1220 -2135 1240 -2115
rect 1260 -2135 1280 -2115
rect 1300 -2135 1320 -2115
rect 1340 -2135 1360 -2115
rect 1380 -2135 1400 -2115
rect 1420 -2135 1440 -2115
rect 1460 -2135 1480 -2115
rect 1500 -2135 1520 -2115
rect 1540 -2135 1560 -2115
rect 1580 -2135 1600 -2115
rect 1620 -2135 1640 -2115
rect 1660 -2135 1680 -2115
rect 1700 -2135 1720 -2115
rect 1740 -2135 1760 -2115
rect 1780 -2135 1800 -2115
rect 1820 -2135 1840 -2115
rect 1860 -2135 1880 -2115
rect 1900 -2135 1920 -2115
rect 1940 -2135 1960 -2115
rect 1980 -2135 2000 -2115
rect 2020 -2135 2040 -2115
rect 2060 -2135 2080 -2115
rect 2100 -2135 2120 -2115
rect 2140 -2135 2160 -2115
rect 2180 -2135 2200 -2115
rect 2220 -2135 2240 -2115
rect 2260 -2135 2280 -2115
rect 2300 -2135 2320 -2115
rect 2340 -2135 2360 -2115
rect 2380 -2135 2400 -2115
rect 2420 -2135 2440 -2115
rect 2460 -2135 2480 -2115
rect 2500 -2135 2520 -2115
rect 2540 -2135 2560 -2115
rect 2590 -2135 2605 -2115
rect 105 -2145 2605 -2135
rect -70 -2160 85 -2150
rect -70 -2185 -60 -2160
rect -40 -2185 -20 -2160
rect 0 -2185 20 -2160
rect 40 -2185 60 -2160
rect -70 -2195 85 -2185
rect 105 -2210 2605 -2200
rect 105 -2230 120 -2210
rect 140 -2230 160 -2210
rect 180 -2230 200 -2210
rect 220 -2230 240 -2210
rect 260 -2230 280 -2210
rect 300 -2230 320 -2210
rect 340 -2230 360 -2210
rect 380 -2230 400 -2210
rect 420 -2230 440 -2210
rect 460 -2230 480 -2210
rect 500 -2230 520 -2210
rect 540 -2230 560 -2210
rect 580 -2230 600 -2210
rect 620 -2230 640 -2210
rect 660 -2230 680 -2210
rect 700 -2230 720 -2210
rect 740 -2230 760 -2210
rect 780 -2230 800 -2210
rect 820 -2230 840 -2210
rect 860 -2230 880 -2210
rect 900 -2230 920 -2210
rect 940 -2230 960 -2210
rect 980 -2230 1000 -2210
rect 1020 -2230 1040 -2210
rect 1060 -2230 1080 -2210
rect 1100 -2230 1120 -2210
rect 1140 -2230 1160 -2210
rect 1180 -2230 1200 -2210
rect 1220 -2230 1240 -2210
rect 1260 -2230 1280 -2210
rect 1300 -2230 1320 -2210
rect 1340 -2230 1360 -2210
rect 1380 -2230 1400 -2210
rect 1420 -2230 1440 -2210
rect 1460 -2230 1480 -2210
rect 1500 -2230 1520 -2210
rect 1540 -2230 1560 -2210
rect 1580 -2230 1600 -2210
rect 1620 -2230 1640 -2210
rect 1660 -2230 1680 -2210
rect 1700 -2230 1720 -2210
rect 1740 -2230 1760 -2210
rect 1780 -2230 1800 -2210
rect 1820 -2230 1840 -2210
rect 1860 -2230 1880 -2210
rect 1900 -2230 1920 -2210
rect 1940 -2230 1960 -2210
rect 1980 -2230 2000 -2210
rect 2020 -2230 2040 -2210
rect 2060 -2230 2080 -2210
rect 2100 -2230 2120 -2210
rect 2140 -2230 2160 -2210
rect 2180 -2230 2200 -2210
rect 2220 -2230 2240 -2210
rect 2260 -2230 2280 -2210
rect 2300 -2230 2320 -2210
rect 2340 -2230 2360 -2210
rect 2380 -2230 2400 -2210
rect 2420 -2230 2440 -2210
rect 2460 -2230 2480 -2210
rect 2500 -2230 2520 -2210
rect 2540 -2230 2560 -2210
rect 2590 -2230 2605 -2210
rect 105 -2240 2605 -2230
rect -70 -2255 85 -2245
rect -70 -2280 -60 -2255
rect -40 -2280 -20 -2255
rect 0 -2280 20 -2255
rect 40 -2280 60 -2255
rect -70 -2290 85 -2280
rect 105 -2305 2605 -2295
rect 105 -2325 120 -2305
rect 140 -2325 160 -2305
rect 180 -2325 200 -2305
rect 220 -2325 240 -2305
rect 260 -2325 280 -2305
rect 300 -2325 320 -2305
rect 340 -2325 360 -2305
rect 380 -2325 400 -2305
rect 420 -2325 440 -2305
rect 460 -2325 480 -2305
rect 500 -2325 520 -2305
rect 540 -2325 560 -2305
rect 580 -2325 600 -2305
rect 620 -2325 640 -2305
rect 660 -2325 680 -2305
rect 700 -2325 720 -2305
rect 740 -2325 760 -2305
rect 780 -2325 800 -2305
rect 820 -2325 840 -2305
rect 860 -2325 880 -2305
rect 900 -2325 920 -2305
rect 940 -2325 960 -2305
rect 980 -2325 1000 -2305
rect 1020 -2325 1040 -2305
rect 1060 -2325 1080 -2305
rect 1100 -2325 1120 -2305
rect 1140 -2325 1160 -2305
rect 1180 -2325 1200 -2305
rect 1220 -2325 1240 -2305
rect 1260 -2325 1280 -2305
rect 1300 -2325 1320 -2305
rect 1340 -2325 1360 -2305
rect 1380 -2325 1400 -2305
rect 1420 -2325 1440 -2305
rect 1460 -2325 1480 -2305
rect 1500 -2325 1520 -2305
rect 1540 -2325 1560 -2305
rect 1580 -2325 1600 -2305
rect 1620 -2325 1640 -2305
rect 1660 -2325 1680 -2305
rect 1700 -2325 1720 -2305
rect 1740 -2325 1760 -2305
rect 1780 -2325 1800 -2305
rect 1820 -2325 1840 -2305
rect 1860 -2325 1880 -2305
rect 1900 -2325 1920 -2305
rect 1940 -2325 1960 -2305
rect 1980 -2325 2000 -2305
rect 2020 -2325 2040 -2305
rect 2060 -2325 2080 -2305
rect 2100 -2325 2120 -2305
rect 2140 -2325 2160 -2305
rect 2180 -2325 2200 -2305
rect 2220 -2325 2240 -2305
rect 2260 -2325 2280 -2305
rect 2300 -2325 2320 -2305
rect 2340 -2325 2360 -2305
rect 2380 -2325 2400 -2305
rect 2420 -2325 2440 -2305
rect 2460 -2325 2480 -2305
rect 2500 -2325 2520 -2305
rect 2540 -2325 2560 -2305
rect 2590 -2325 2605 -2305
rect 105 -2335 2605 -2325
rect -70 -2350 85 -2340
rect -70 -2375 -60 -2350
rect -40 -2375 -20 -2350
rect 0 -2375 20 -2350
rect 40 -2375 60 -2350
rect -70 -2385 85 -2375
rect 105 -2400 2605 -2390
rect 105 -2420 120 -2400
rect 140 -2420 160 -2400
rect 180 -2420 200 -2400
rect 220 -2420 240 -2400
rect 260 -2420 280 -2400
rect 300 -2420 320 -2400
rect 340 -2420 360 -2400
rect 380 -2420 400 -2400
rect 420 -2420 440 -2400
rect 460 -2420 480 -2400
rect 500 -2420 520 -2400
rect 540 -2420 560 -2400
rect 580 -2420 600 -2400
rect 620 -2420 640 -2400
rect 660 -2420 680 -2400
rect 700 -2420 720 -2400
rect 740 -2420 760 -2400
rect 780 -2420 800 -2400
rect 820 -2420 840 -2400
rect 860 -2420 880 -2400
rect 900 -2420 920 -2400
rect 940 -2420 960 -2400
rect 980 -2420 1000 -2400
rect 1020 -2420 1040 -2400
rect 1060 -2420 1080 -2400
rect 1100 -2420 1120 -2400
rect 1140 -2420 1160 -2400
rect 1180 -2420 1200 -2400
rect 1220 -2420 1240 -2400
rect 1260 -2420 1280 -2400
rect 1300 -2420 1320 -2400
rect 1340 -2420 1360 -2400
rect 1380 -2420 1400 -2400
rect 1420 -2420 1440 -2400
rect 1460 -2420 1480 -2400
rect 1500 -2420 1520 -2400
rect 1540 -2420 1560 -2400
rect 1580 -2420 1600 -2400
rect 1620 -2420 1640 -2400
rect 1660 -2420 1680 -2400
rect 1700 -2420 1720 -2400
rect 1740 -2420 1760 -2400
rect 1780 -2420 1800 -2400
rect 1820 -2420 1840 -2400
rect 1860 -2420 1880 -2400
rect 1900 -2420 1920 -2400
rect 1940 -2420 1960 -2400
rect 1980 -2420 2000 -2400
rect 2020 -2420 2040 -2400
rect 2060 -2420 2080 -2400
rect 2100 -2420 2120 -2400
rect 2140 -2420 2160 -2400
rect 2180 -2420 2200 -2400
rect 2220 -2420 2240 -2400
rect 2260 -2420 2280 -2400
rect 2300 -2420 2320 -2400
rect 2340 -2420 2360 -2400
rect 2380 -2420 2400 -2400
rect 2420 -2420 2440 -2400
rect 2460 -2420 2480 -2400
rect 2500 -2420 2520 -2400
rect 2540 -2420 2560 -2400
rect 2590 -2420 2605 -2400
rect 105 -2430 2605 -2420
rect -70 -2445 85 -2435
rect -70 -2470 -60 -2445
rect -40 -2470 -20 -2445
rect 0 -2470 20 -2445
rect 40 -2470 60 -2445
rect -70 -2480 85 -2470
rect 105 -2495 2605 -2485
rect 105 -2515 120 -2495
rect 140 -2515 160 -2495
rect 180 -2515 200 -2495
rect 220 -2515 240 -2495
rect 260 -2515 280 -2495
rect 300 -2515 320 -2495
rect 340 -2515 360 -2495
rect 380 -2515 400 -2495
rect 420 -2515 440 -2495
rect 460 -2515 480 -2495
rect 500 -2515 520 -2495
rect 540 -2515 560 -2495
rect 580 -2515 600 -2495
rect 620 -2515 640 -2495
rect 660 -2515 680 -2495
rect 700 -2515 720 -2495
rect 740 -2515 760 -2495
rect 780 -2515 800 -2495
rect 820 -2515 840 -2495
rect 860 -2515 880 -2495
rect 900 -2515 920 -2495
rect 940 -2515 960 -2495
rect 980 -2515 1000 -2495
rect 1020 -2515 1040 -2495
rect 1060 -2515 1080 -2495
rect 1100 -2515 1120 -2495
rect 1140 -2515 1160 -2495
rect 1180 -2515 1200 -2495
rect 1220 -2515 1240 -2495
rect 1260 -2515 1280 -2495
rect 1300 -2515 1320 -2495
rect 1340 -2515 1360 -2495
rect 1380 -2515 1400 -2495
rect 1420 -2515 1440 -2495
rect 1460 -2515 1480 -2495
rect 1500 -2515 1520 -2495
rect 1540 -2515 1560 -2495
rect 1580 -2515 1600 -2495
rect 1620 -2515 1640 -2495
rect 1660 -2515 1680 -2495
rect 1700 -2515 1720 -2495
rect 1740 -2515 1760 -2495
rect 1780 -2515 1800 -2495
rect 1820 -2515 1840 -2495
rect 1860 -2515 1880 -2495
rect 1900 -2515 1920 -2495
rect 1940 -2515 1960 -2495
rect 1980 -2515 2000 -2495
rect 2020 -2515 2040 -2495
rect 2060 -2515 2080 -2495
rect 2100 -2515 2120 -2495
rect 2140 -2515 2160 -2495
rect 2180 -2515 2200 -2495
rect 2220 -2515 2240 -2495
rect 2260 -2515 2280 -2495
rect 2300 -2515 2320 -2495
rect 2340 -2515 2360 -2495
rect 2380 -2515 2400 -2495
rect 2420 -2515 2440 -2495
rect 2460 -2515 2480 -2495
rect 2500 -2515 2520 -2495
rect 2540 -2515 2560 -2495
rect 2590 -2515 2605 -2495
rect 105 -2525 2605 -2515
rect -70 -2540 85 -2530
rect -70 -2565 -60 -2540
rect -40 -2565 -20 -2540
rect 0 -2565 20 -2540
rect 40 -2565 60 -2540
rect -70 -2575 85 -2565
rect 105 -2590 2605 -2580
rect 105 -2610 120 -2590
rect 140 -2610 160 -2590
rect 180 -2610 200 -2590
rect 220 -2610 240 -2590
rect 260 -2610 280 -2590
rect 300 -2610 320 -2590
rect 340 -2610 360 -2590
rect 380 -2610 400 -2590
rect 420 -2610 440 -2590
rect 460 -2610 480 -2590
rect 500 -2610 520 -2590
rect 540 -2610 560 -2590
rect 580 -2610 600 -2590
rect 620 -2610 640 -2590
rect 660 -2610 680 -2590
rect 700 -2610 720 -2590
rect 740 -2610 760 -2590
rect 780 -2610 800 -2590
rect 820 -2610 840 -2590
rect 860 -2610 880 -2590
rect 900 -2610 920 -2590
rect 940 -2610 960 -2590
rect 980 -2610 1000 -2590
rect 1020 -2610 1040 -2590
rect 1060 -2610 1080 -2590
rect 1100 -2610 1120 -2590
rect 1140 -2610 1160 -2590
rect 1180 -2610 1200 -2590
rect 1220 -2610 1240 -2590
rect 1260 -2610 1280 -2590
rect 1300 -2610 1320 -2590
rect 1340 -2610 1360 -2590
rect 1380 -2610 1400 -2590
rect 1420 -2610 1440 -2590
rect 1460 -2610 1480 -2590
rect 1500 -2610 1520 -2590
rect 1540 -2610 1560 -2590
rect 1580 -2610 1600 -2590
rect 1620 -2610 1640 -2590
rect 1660 -2610 1680 -2590
rect 1700 -2610 1720 -2590
rect 1740 -2610 1760 -2590
rect 1780 -2610 1800 -2590
rect 1820 -2610 1840 -2590
rect 1860 -2610 1880 -2590
rect 1900 -2610 1920 -2590
rect 1940 -2610 1960 -2590
rect 1980 -2610 2000 -2590
rect 2020 -2610 2040 -2590
rect 2060 -2610 2080 -2590
rect 2100 -2610 2120 -2590
rect 2140 -2610 2160 -2590
rect 2180 -2610 2200 -2590
rect 2220 -2610 2240 -2590
rect 2260 -2610 2280 -2590
rect 2300 -2610 2320 -2590
rect 2340 -2610 2360 -2590
rect 2380 -2610 2400 -2590
rect 2420 -2610 2440 -2590
rect 2460 -2610 2480 -2590
rect 2500 -2610 2520 -2590
rect 2540 -2610 2560 -2590
rect 2590 -2610 2605 -2590
rect 105 -2620 2605 -2610
rect -70 -2635 85 -2625
rect -70 -2660 -60 -2635
rect -40 -2660 -20 -2635
rect 0 -2660 20 -2635
rect 40 -2660 60 -2635
rect -70 -2670 85 -2660
rect 105 -2685 2605 -2675
rect 105 -2705 120 -2685
rect 140 -2705 160 -2685
rect 180 -2705 200 -2685
rect 220 -2705 240 -2685
rect 260 -2705 280 -2685
rect 300 -2705 320 -2685
rect 340 -2705 360 -2685
rect 380 -2705 400 -2685
rect 420 -2705 440 -2685
rect 460 -2705 480 -2685
rect 500 -2705 520 -2685
rect 540 -2705 560 -2685
rect 580 -2705 600 -2685
rect 620 -2705 640 -2685
rect 660 -2705 680 -2685
rect 700 -2705 720 -2685
rect 740 -2705 760 -2685
rect 780 -2705 800 -2685
rect 820 -2705 840 -2685
rect 860 -2705 880 -2685
rect 900 -2705 920 -2685
rect 940 -2705 960 -2685
rect 980 -2705 1000 -2685
rect 1020 -2705 1040 -2685
rect 1060 -2705 1080 -2685
rect 1100 -2705 1120 -2685
rect 1140 -2705 1160 -2685
rect 1180 -2705 1200 -2685
rect 1220 -2705 1240 -2685
rect 1260 -2705 1280 -2685
rect 1300 -2705 1320 -2685
rect 1340 -2705 1360 -2685
rect 1380 -2705 1400 -2685
rect 1420 -2705 1440 -2685
rect 1460 -2705 1480 -2685
rect 1500 -2705 1520 -2685
rect 1540 -2705 1560 -2685
rect 1580 -2705 1600 -2685
rect 1620 -2705 1640 -2685
rect 1660 -2705 1680 -2685
rect 1700 -2705 1720 -2685
rect 1740 -2705 1760 -2685
rect 1780 -2705 1800 -2685
rect 1820 -2705 1840 -2685
rect 1860 -2705 1880 -2685
rect 1900 -2705 1920 -2685
rect 1940 -2705 1960 -2685
rect 1980 -2705 2000 -2685
rect 2020 -2705 2040 -2685
rect 2060 -2705 2080 -2685
rect 2100 -2705 2120 -2685
rect 2140 -2705 2160 -2685
rect 2180 -2705 2200 -2685
rect 2220 -2705 2240 -2685
rect 2260 -2705 2280 -2685
rect 2300 -2705 2320 -2685
rect 2340 -2705 2360 -2685
rect 2380 -2705 2400 -2685
rect 2420 -2705 2440 -2685
rect 2460 -2705 2480 -2685
rect 2500 -2705 2520 -2685
rect 2540 -2705 2560 -2685
rect 2590 -2705 2605 -2685
rect 105 -2725 2605 -2705
rect 105 -2745 120 -2725
rect 140 -2745 160 -2725
rect 180 -2745 200 -2725
rect 220 -2745 240 -2725
rect 260 -2745 280 -2725
rect 300 -2745 320 -2725
rect 340 -2745 360 -2725
rect 380 -2745 400 -2725
rect 420 -2745 440 -2725
rect 460 -2745 480 -2725
rect 500 -2745 520 -2725
rect 540 -2745 560 -2725
rect 580 -2745 600 -2725
rect 620 -2745 640 -2725
rect 660 -2745 680 -2725
rect 700 -2745 720 -2725
rect 740 -2745 760 -2725
rect 780 -2745 800 -2725
rect 820 -2745 840 -2725
rect 860 -2745 880 -2725
rect 900 -2745 920 -2725
rect 940 -2745 960 -2725
rect 980 -2745 1000 -2725
rect 1020 -2745 1040 -2725
rect 1060 -2745 1080 -2725
rect 1100 -2745 1120 -2725
rect 1140 -2745 1160 -2725
rect 1180 -2745 1200 -2725
rect 1220 -2745 1240 -2725
rect 1260 -2745 1280 -2725
rect 1300 -2745 1320 -2725
rect 1340 -2745 1360 -2725
rect 1380 -2745 1400 -2725
rect 1420 -2745 1440 -2725
rect 1460 -2745 1480 -2725
rect 1500 -2745 1520 -2725
rect 1540 -2745 1560 -2725
rect 1580 -2745 1600 -2725
rect 1620 -2745 1640 -2725
rect 1660 -2745 1680 -2725
rect 1700 -2745 1720 -2725
rect 1740 -2745 1760 -2725
rect 1780 -2745 1800 -2725
rect 1820 -2745 1840 -2725
rect 1860 -2745 1880 -2725
rect 1900 -2745 1920 -2725
rect 1940 -2745 1960 -2725
rect 1980 -2745 2000 -2725
rect 2020 -2745 2040 -2725
rect 2060 -2745 2080 -2725
rect 2100 -2745 2120 -2725
rect 2140 -2745 2160 -2725
rect 2180 -2745 2200 -2725
rect 2220 -2745 2240 -2725
rect 2260 -2745 2280 -2725
rect 2300 -2745 2320 -2725
rect 2340 -2745 2360 -2725
rect 2380 -2745 2400 -2725
rect 2420 -2745 2440 -2725
rect 2460 -2745 2480 -2725
rect 2500 -2745 2520 -2725
rect 2540 -2745 2560 -2725
rect 2590 -2745 2605 -2725
rect 105 -2755 2605 -2745
<< viali >>
rect 1780 2325 1800 2345
rect 1820 2325 1840 2345
rect 1860 2325 1880 2345
rect 1900 2325 1920 2345
rect 1940 2325 1960 2345
rect 1980 2325 2000 2345
rect 2020 2325 2040 2345
rect 2060 2325 2080 2345
rect 2100 2325 2120 2345
rect 2140 2325 2160 2345
rect 2180 2325 2200 2345
rect 2220 2325 2240 2345
rect 2260 2325 2280 2345
rect 2300 2325 2320 2345
rect 2340 2325 2360 2345
rect 2380 2325 2400 2345
rect 2420 2325 2440 2345
rect 2460 2325 2480 2345
rect 2500 2325 2520 2345
rect 680 2240 700 2260
rect 720 2240 740 2260
rect 760 2240 780 2260
rect 800 2240 820 2260
rect 840 2240 860 2260
rect 880 2240 900 2260
rect 920 2240 940 2260
rect 960 2240 980 2260
rect 1000 2240 1020 2260
rect 1040 2240 1060 2260
rect 1080 2240 1100 2260
rect 1120 2240 1140 2260
rect 1160 2240 1180 2260
rect 1200 2240 1220 2260
rect 1240 2240 1260 2260
rect 1280 2240 1300 2260
rect 1320 2240 1340 2260
rect 1360 2240 1380 2260
rect 1400 2240 1420 2260
rect 1440 2240 1460 2260
rect 680 2197 700 2217
rect 720 2197 740 2217
rect 760 2197 780 2217
rect 800 2197 820 2217
rect 840 2197 860 2217
rect 880 2197 900 2217
rect 920 2197 940 2217
rect 960 2197 980 2217
rect 1000 2197 1020 2217
rect 1040 2197 1060 2217
rect 1080 2197 1100 2217
rect 1120 2197 1140 2217
rect 1160 2197 1180 2217
rect 1200 2197 1220 2217
rect 1240 2197 1260 2217
rect 1280 2197 1300 2217
rect 1320 2197 1340 2217
rect 1360 2197 1380 2217
rect 1400 2197 1420 2217
rect 1440 2197 1460 2217
rect 10 2155 30 2175
rect 50 2155 70 2175
rect 90 2155 110 2175
rect 130 2155 150 2175
rect 1760 2115 1780 2135
rect 1800 2115 1820 2135
rect 1840 2115 1860 2135
rect 1880 2115 1900 2135
rect 1920 2115 1940 2135
rect 1960 2115 1980 2135
rect 2000 2115 2020 2135
rect 2040 2115 2060 2135
rect 2080 2115 2100 2135
rect 2120 2115 2140 2135
rect 2160 2115 2180 2135
rect 2200 2115 2220 2135
rect 2240 2115 2260 2135
rect 2280 2115 2300 2135
rect 2320 2115 2340 2135
rect 2360 2115 2380 2135
rect 2400 2115 2420 2135
rect 2440 2115 2460 2135
rect 2480 2115 2500 2135
rect 2520 2115 2540 2135
rect 10 2075 30 2095
rect 50 2075 70 2095
rect 90 2075 110 2095
rect 130 2075 150 2095
rect 680 2033 700 2053
rect 720 2033 740 2053
rect 760 2033 780 2053
rect 800 2033 820 2053
rect 840 2033 860 2053
rect 880 2033 900 2053
rect 920 2033 940 2053
rect 960 2033 980 2053
rect 1000 2033 1020 2053
rect 1040 2033 1060 2053
rect 1080 2033 1100 2053
rect 1120 2033 1140 2053
rect 1160 2033 1180 2053
rect 1200 2033 1220 2053
rect 1240 2033 1260 2053
rect 1280 2033 1300 2053
rect 1320 2033 1340 2053
rect 1360 2033 1380 2053
rect 1400 2033 1420 2053
rect 1440 2033 1460 2053
rect 10 1990 30 2010
rect 50 1990 70 2010
rect 90 1990 110 2010
rect 130 1990 150 2010
rect 1760 1951 1780 1971
rect 1800 1951 1820 1971
rect 1840 1951 1860 1971
rect 1880 1951 1900 1971
rect 1920 1951 1940 1971
rect 1960 1951 1980 1971
rect 2000 1951 2020 1971
rect 2040 1951 2060 1971
rect 2080 1951 2100 1971
rect 2120 1951 2140 1971
rect 2160 1951 2180 1971
rect 2200 1951 2220 1971
rect 2240 1951 2260 1971
rect 2280 1951 2300 1971
rect 2320 1951 2340 1971
rect 2360 1951 2380 1971
rect 2400 1951 2420 1971
rect 2440 1951 2460 1971
rect 2480 1951 2500 1971
rect 2520 1951 2540 1971
rect 10 1910 30 1930
rect 50 1910 70 1930
rect 90 1910 110 1930
rect 130 1910 150 1930
rect 680 1869 700 1889
rect 720 1869 740 1889
rect 760 1869 780 1889
rect 800 1869 820 1889
rect 840 1869 860 1889
rect 880 1869 900 1889
rect 920 1869 940 1889
rect 960 1869 980 1889
rect 1000 1869 1020 1889
rect 1040 1869 1060 1889
rect 1080 1869 1100 1889
rect 1120 1869 1140 1889
rect 1160 1869 1180 1889
rect 1200 1869 1220 1889
rect 1240 1869 1260 1889
rect 1280 1869 1300 1889
rect 1320 1869 1340 1889
rect 1360 1869 1380 1889
rect 1400 1869 1420 1889
rect 1440 1869 1460 1889
rect 10 1830 30 1850
rect 50 1830 70 1850
rect 90 1830 110 1850
rect 130 1830 150 1850
rect 1760 1787 1780 1807
rect 1800 1787 1820 1807
rect 1840 1787 1860 1807
rect 1880 1787 1900 1807
rect 1920 1787 1940 1807
rect 1960 1787 1980 1807
rect 2000 1787 2020 1807
rect 2040 1787 2060 1807
rect 2080 1787 2100 1807
rect 2120 1787 2140 1807
rect 2160 1787 2180 1807
rect 2200 1787 2220 1807
rect 2240 1787 2260 1807
rect 2280 1787 2300 1807
rect 2320 1787 2340 1807
rect 2360 1787 2380 1807
rect 2400 1787 2420 1807
rect 2440 1787 2460 1807
rect 2480 1787 2500 1807
rect 2520 1787 2540 1807
rect 10 1745 30 1765
rect 50 1745 70 1765
rect 90 1745 110 1765
rect 130 1745 150 1765
rect 680 1705 700 1725
rect 720 1705 740 1725
rect 760 1705 780 1725
rect 800 1705 820 1725
rect 840 1705 860 1725
rect 880 1705 900 1725
rect 920 1705 940 1725
rect 960 1705 980 1725
rect 1000 1705 1020 1725
rect 1040 1705 1060 1725
rect 1080 1705 1100 1725
rect 1120 1705 1140 1725
rect 1160 1705 1180 1725
rect 1200 1705 1220 1725
rect 1240 1705 1260 1725
rect 1280 1705 1300 1725
rect 1320 1705 1340 1725
rect 1360 1705 1380 1725
rect 1400 1705 1420 1725
rect 1440 1705 1460 1725
rect 10 1665 30 1685
rect 50 1665 70 1685
rect 90 1665 110 1685
rect 130 1665 150 1685
rect 1760 1623 1780 1643
rect 1800 1623 1820 1643
rect 1840 1623 1860 1643
rect 1880 1623 1900 1643
rect 1920 1623 1940 1643
rect 1960 1623 1980 1643
rect 2000 1623 2020 1643
rect 2040 1623 2060 1643
rect 2080 1623 2100 1643
rect 2120 1623 2140 1643
rect 2160 1623 2180 1643
rect 2200 1623 2220 1643
rect 2240 1623 2260 1643
rect 2280 1623 2300 1643
rect 2320 1623 2340 1643
rect 2360 1623 2380 1643
rect 2400 1623 2420 1643
rect 2440 1623 2460 1643
rect 2480 1623 2500 1643
rect 2520 1623 2540 1643
rect 10 1580 30 1600
rect 50 1580 70 1600
rect 90 1580 110 1600
rect 130 1580 150 1600
rect 680 1541 700 1561
rect 720 1541 740 1561
rect 760 1541 780 1561
rect 800 1541 820 1561
rect 840 1541 860 1561
rect 880 1541 900 1561
rect 920 1541 940 1561
rect 960 1541 980 1561
rect 1000 1541 1020 1561
rect 1040 1541 1060 1561
rect 1080 1541 1100 1561
rect 1120 1541 1140 1561
rect 1160 1541 1180 1561
rect 1200 1541 1220 1561
rect 1240 1541 1260 1561
rect 1280 1541 1300 1561
rect 1320 1541 1340 1561
rect 1360 1541 1380 1561
rect 1400 1541 1420 1561
rect 1440 1541 1460 1561
rect 10 1500 30 1520
rect 50 1500 70 1520
rect 90 1500 110 1520
rect 130 1500 150 1520
rect 1760 1459 1780 1479
rect 1800 1459 1820 1479
rect 1840 1459 1860 1479
rect 1880 1459 1900 1479
rect 1920 1459 1940 1479
rect 1960 1459 1980 1479
rect 2000 1459 2020 1479
rect 2040 1459 2060 1479
rect 2080 1459 2100 1479
rect 2120 1459 2140 1479
rect 2160 1459 2180 1479
rect 2200 1459 2220 1479
rect 2240 1459 2260 1479
rect 2280 1459 2300 1479
rect 2320 1459 2340 1479
rect 2360 1459 2380 1479
rect 2400 1459 2420 1479
rect 2440 1459 2460 1479
rect 2480 1459 2500 1479
rect 2520 1459 2540 1479
rect 10 1420 30 1440
rect 50 1420 70 1440
rect 90 1420 110 1440
rect 130 1420 150 1440
rect 680 1377 700 1397
rect 720 1377 740 1397
rect 760 1377 780 1397
rect 800 1377 820 1397
rect 840 1377 860 1397
rect 880 1377 900 1397
rect 920 1377 940 1397
rect 960 1377 980 1397
rect 1000 1377 1020 1397
rect 1040 1377 1060 1397
rect 1080 1377 1100 1397
rect 1120 1377 1140 1397
rect 1160 1377 1180 1397
rect 1200 1377 1220 1397
rect 1240 1377 1260 1397
rect 1280 1377 1300 1397
rect 1320 1377 1340 1397
rect 1360 1377 1380 1397
rect 1400 1377 1420 1397
rect 1440 1377 1460 1397
rect 10 1335 30 1355
rect 50 1335 70 1355
rect 90 1335 110 1355
rect 130 1335 150 1355
rect 1760 1295 1780 1315
rect 1800 1295 1820 1315
rect 1840 1295 1860 1315
rect 1880 1295 1900 1315
rect 1920 1295 1940 1315
rect 1960 1295 1980 1315
rect 2000 1295 2020 1315
rect 2040 1295 2060 1315
rect 2080 1295 2100 1315
rect 2120 1295 2140 1315
rect 2160 1295 2180 1315
rect 2200 1295 2220 1315
rect 2240 1295 2260 1315
rect 2280 1295 2300 1315
rect 2320 1295 2340 1315
rect 2360 1295 2380 1315
rect 2400 1295 2420 1315
rect 2440 1295 2460 1315
rect 2480 1295 2500 1315
rect 2520 1295 2540 1315
rect 10 1255 30 1275
rect 50 1255 70 1275
rect 90 1255 110 1275
rect 130 1255 150 1275
rect 680 1213 700 1233
rect 720 1213 740 1233
rect 760 1213 780 1233
rect 800 1213 820 1233
rect 840 1213 860 1233
rect 880 1213 900 1233
rect 920 1213 940 1233
rect 960 1213 980 1233
rect 1000 1213 1020 1233
rect 1040 1213 1060 1233
rect 1080 1213 1100 1233
rect 1120 1213 1140 1233
rect 1160 1213 1180 1233
rect 1200 1213 1220 1233
rect 1240 1213 1260 1233
rect 1280 1213 1300 1233
rect 1320 1213 1340 1233
rect 1360 1213 1380 1233
rect 1400 1213 1420 1233
rect 1440 1213 1460 1233
rect 10 1170 30 1190
rect 50 1170 70 1190
rect 90 1170 110 1190
rect 130 1170 150 1190
rect 1760 1131 1780 1151
rect 1800 1131 1820 1151
rect 1840 1131 1860 1151
rect 1880 1131 1900 1151
rect 1920 1131 1940 1151
rect 1960 1131 1980 1151
rect 2000 1131 2020 1151
rect 2040 1131 2060 1151
rect 2080 1131 2100 1151
rect 2120 1131 2140 1151
rect 2160 1131 2180 1151
rect 2200 1131 2220 1151
rect 2240 1131 2260 1151
rect 2280 1131 2300 1151
rect 2320 1131 2340 1151
rect 2360 1131 2380 1151
rect 2400 1131 2420 1151
rect 2440 1131 2460 1151
rect 2480 1131 2500 1151
rect 2520 1131 2540 1151
rect 10 1090 30 1110
rect 50 1090 70 1110
rect 90 1090 110 1110
rect 130 1090 150 1110
rect 680 1049 700 1069
rect 720 1049 740 1069
rect 760 1049 780 1069
rect 800 1049 820 1069
rect 840 1049 860 1069
rect 880 1049 900 1069
rect 920 1049 940 1069
rect 960 1049 980 1069
rect 1000 1049 1020 1069
rect 1040 1049 1060 1069
rect 1080 1049 1100 1069
rect 1120 1049 1140 1069
rect 1160 1049 1180 1069
rect 1200 1049 1220 1069
rect 1240 1049 1260 1069
rect 1280 1049 1300 1069
rect 1320 1049 1340 1069
rect 1360 1049 1380 1069
rect 1400 1049 1420 1069
rect 1440 1049 1460 1069
rect 10 1010 30 1030
rect 50 1010 70 1030
rect 90 1010 110 1030
rect 130 1010 150 1030
rect 1760 967 1780 987
rect 1800 967 1820 987
rect 1840 967 1860 987
rect 1880 967 1900 987
rect 1920 967 1940 987
rect 1960 967 1980 987
rect 2000 967 2020 987
rect 2040 967 2060 987
rect 2080 967 2100 987
rect 2120 967 2140 987
rect 2160 967 2180 987
rect 2200 967 2220 987
rect 2240 967 2260 987
rect 2280 967 2300 987
rect 2320 967 2340 987
rect 2360 967 2380 987
rect 2400 967 2420 987
rect 2440 967 2460 987
rect 2480 967 2500 987
rect 2520 967 2540 987
rect 10 925 30 945
rect 50 925 70 945
rect 90 925 110 945
rect 130 925 150 945
rect 680 885 700 905
rect 720 885 740 905
rect 760 885 780 905
rect 800 885 820 905
rect 840 885 860 905
rect 880 885 900 905
rect 920 885 940 905
rect 960 885 980 905
rect 1000 885 1020 905
rect 1040 885 1060 905
rect 1080 885 1100 905
rect 1120 885 1140 905
rect 1160 885 1180 905
rect 1200 885 1220 905
rect 1240 885 1260 905
rect 1280 885 1300 905
rect 1320 885 1340 905
rect 1360 885 1380 905
rect 1400 885 1420 905
rect 1440 885 1460 905
rect 10 845 30 865
rect 50 845 70 865
rect 90 845 110 865
rect 130 845 150 865
rect 1760 803 1780 823
rect 1800 803 1820 823
rect 1840 803 1860 823
rect 1880 803 1900 823
rect 1920 803 1940 823
rect 1960 803 1980 823
rect 2000 803 2020 823
rect 2040 803 2060 823
rect 2080 803 2100 823
rect 2120 803 2140 823
rect 2160 803 2180 823
rect 2200 803 2220 823
rect 2240 803 2260 823
rect 2280 803 2300 823
rect 2320 803 2340 823
rect 2360 803 2380 823
rect 2400 803 2420 823
rect 2440 803 2460 823
rect 2480 803 2500 823
rect 2520 803 2540 823
rect 10 760 30 780
rect 50 760 70 780
rect 90 760 110 780
rect 130 760 150 780
rect 680 721 700 741
rect 720 721 740 741
rect 760 721 780 741
rect 800 721 820 741
rect 840 721 860 741
rect 880 721 900 741
rect 920 721 940 741
rect 960 721 980 741
rect 1000 721 1020 741
rect 1040 721 1060 741
rect 1080 721 1100 741
rect 1120 721 1140 741
rect 1160 721 1180 741
rect 1200 721 1220 741
rect 1240 721 1260 741
rect 1280 721 1300 741
rect 1320 721 1340 741
rect 1360 721 1380 741
rect 1400 721 1420 741
rect 1440 721 1460 741
rect 10 680 30 700
rect 50 680 70 700
rect 90 680 110 700
rect 130 680 150 700
rect 1760 639 1780 659
rect 1800 639 1820 659
rect 1840 639 1860 659
rect 1880 639 1900 659
rect 1920 639 1940 659
rect 1960 639 1980 659
rect 2000 639 2020 659
rect 2040 639 2060 659
rect 2080 639 2100 659
rect 2120 639 2140 659
rect 2160 639 2180 659
rect 2200 639 2220 659
rect 2240 639 2260 659
rect 2280 639 2300 659
rect 2320 639 2340 659
rect 2360 639 2380 659
rect 2400 639 2420 659
rect 2440 639 2460 659
rect 2480 639 2500 659
rect 2520 639 2540 659
rect 10 600 30 620
rect 50 600 70 620
rect 90 600 110 620
rect 130 600 150 620
rect 680 557 700 577
rect 720 557 740 577
rect 760 557 780 577
rect 800 557 820 577
rect 840 557 860 577
rect 880 557 900 577
rect 920 557 940 577
rect 960 557 980 577
rect 1000 557 1020 577
rect 1040 557 1060 577
rect 1080 557 1100 577
rect 1120 557 1140 577
rect 1160 557 1180 577
rect 1200 557 1220 577
rect 1240 557 1260 577
rect 1280 557 1300 577
rect 1320 557 1340 577
rect 1360 557 1380 577
rect 1400 557 1420 577
rect 1440 557 1460 577
rect 10 515 30 535
rect 50 515 70 535
rect 90 515 110 535
rect 130 515 150 535
rect 1760 475 1780 495
rect 1800 475 1820 495
rect 1840 475 1860 495
rect 1880 475 1900 495
rect 1920 475 1940 495
rect 1960 475 1980 495
rect 2000 475 2020 495
rect 2040 475 2060 495
rect 2080 475 2100 495
rect 2120 475 2140 495
rect 2160 475 2180 495
rect 2200 475 2220 495
rect 2240 475 2260 495
rect 2280 475 2300 495
rect 2320 475 2340 495
rect 2360 475 2380 495
rect 2400 475 2420 495
rect 2440 475 2460 495
rect 2480 475 2500 495
rect 2520 475 2540 495
rect 10 435 30 455
rect 50 435 70 455
rect 90 435 110 455
rect 130 435 150 455
rect 680 393 700 413
rect 720 393 740 413
rect 760 393 780 413
rect 800 393 820 413
rect 840 393 860 413
rect 880 393 900 413
rect 920 393 940 413
rect 960 393 980 413
rect 1000 393 1020 413
rect 1040 393 1060 413
rect 1080 393 1100 413
rect 1120 393 1140 413
rect 1160 393 1180 413
rect 1200 393 1220 413
rect 1240 393 1260 413
rect 1280 393 1300 413
rect 1320 393 1340 413
rect 1360 393 1380 413
rect 1400 393 1420 413
rect 1440 393 1460 413
rect 10 355 30 375
rect 50 355 70 375
rect 90 355 110 375
rect 130 355 150 375
rect 1760 311 1780 331
rect 1800 311 1820 331
rect 1840 311 1860 331
rect 1880 311 1900 331
rect 1920 311 1940 331
rect 1960 311 1980 331
rect 2000 311 2020 331
rect 2040 311 2060 331
rect 2080 311 2100 331
rect 2120 311 2140 331
rect 2160 311 2180 331
rect 2200 311 2220 331
rect 2240 311 2260 331
rect 2280 311 2300 331
rect 2320 311 2340 331
rect 2360 311 2380 331
rect 2400 311 2420 331
rect 2440 311 2460 331
rect 2480 311 2500 331
rect 2520 311 2540 331
rect 10 270 30 290
rect 50 270 70 290
rect 90 270 110 290
rect 130 270 150 290
rect 680 229 700 249
rect 720 229 740 249
rect 760 229 780 249
rect 800 229 820 249
rect 840 229 860 249
rect 880 229 900 249
rect 920 229 940 249
rect 960 229 980 249
rect 1000 229 1020 249
rect 1040 229 1060 249
rect 1080 229 1100 249
rect 1120 229 1140 249
rect 1160 229 1180 249
rect 1200 229 1220 249
rect 1240 229 1260 249
rect 1280 229 1300 249
rect 1320 229 1340 249
rect 1360 229 1380 249
rect 1400 229 1420 249
rect 1440 229 1460 249
rect 10 190 30 210
rect 50 190 70 210
rect 90 190 110 210
rect 130 190 150 210
rect 1760 147 1780 167
rect 1800 147 1820 167
rect 1840 147 1860 167
rect 1880 147 1900 167
rect 1920 147 1940 167
rect 1960 147 1980 167
rect 2000 147 2020 167
rect 2040 147 2060 167
rect 2080 147 2100 167
rect 2120 147 2140 167
rect 2160 147 2180 167
rect 2200 147 2220 167
rect 2240 147 2260 167
rect 2280 147 2300 167
rect 2320 147 2340 167
rect 2360 147 2380 167
rect 2400 147 2420 167
rect 2440 147 2460 167
rect 2480 147 2500 167
rect 2520 147 2540 167
rect 10 110 30 130
rect 50 110 70 130
rect 90 110 110 130
rect 130 110 150 130
rect 680 65 700 85
rect 720 65 740 85
rect 760 65 780 85
rect 800 65 820 85
rect 840 65 860 85
rect 880 65 900 85
rect 920 65 940 85
rect 960 65 980 85
rect 1000 65 1020 85
rect 1040 65 1060 85
rect 1080 65 1100 85
rect 1120 65 1140 85
rect 1160 65 1180 85
rect 1200 65 1220 85
rect 1240 65 1260 85
rect 1280 65 1300 85
rect 1320 65 1340 85
rect 1360 65 1380 85
rect 1400 65 1420 85
rect 1440 65 1460 85
rect 680 25 700 45
rect 720 25 740 45
rect 760 25 780 45
rect 800 25 820 45
rect 840 25 860 45
rect 880 25 900 45
rect 920 25 940 45
rect 960 25 980 45
rect 1000 25 1020 45
rect 1040 25 1060 45
rect 1080 25 1100 45
rect 1120 25 1140 45
rect 1160 25 1180 45
rect 1200 25 1220 45
rect 1240 25 1260 45
rect 1280 25 1300 45
rect 1320 25 1340 45
rect 1360 25 1380 45
rect 1400 25 1420 45
rect 1440 25 1460 45
rect 1760 -195 1780 -175
rect 1800 -195 1820 -175
rect 1840 -195 1860 -175
rect 1880 -195 1900 -175
rect 1920 -195 1940 -175
rect 1960 -195 1980 -175
rect 2000 -195 2020 -175
rect 2040 -195 2060 -175
rect 2080 -195 2100 -175
rect 2120 -195 2140 -175
rect 2160 -195 2180 -175
rect 2200 -195 2220 -175
rect 2240 -195 2260 -175
rect 2280 -195 2300 -175
rect 2320 -195 2340 -175
rect 2360 -195 2380 -175
rect 2400 -195 2420 -175
rect 2440 -195 2460 -175
rect 2480 -195 2500 -175
rect 2520 -195 2540 -175
rect 1760 -235 1780 -215
rect 1800 -235 1820 -215
rect 1840 -235 1860 -215
rect 1880 -235 1900 -215
rect 1920 -235 1940 -215
rect 1960 -235 1980 -215
rect 2000 -235 2020 -215
rect 2040 -235 2060 -215
rect 2080 -235 2100 -215
rect 2120 -235 2140 -215
rect 2160 -235 2180 -215
rect 2200 -235 2220 -215
rect 2240 -235 2260 -215
rect 2280 -235 2300 -215
rect 2320 -235 2340 -215
rect 2360 -235 2380 -215
rect 2400 -235 2420 -215
rect 2440 -235 2460 -215
rect 2480 -235 2500 -215
rect 2520 -235 2540 -215
rect -60 -285 -40 -260
rect -20 -285 0 -260
rect 20 -285 40 -260
rect 60 -285 80 -260
rect 680 -330 700 -310
rect 720 -330 740 -310
rect 760 -330 780 -310
rect 800 -330 820 -310
rect 840 -330 860 -310
rect 880 -330 900 -310
rect 920 -330 940 -310
rect 960 -330 980 -310
rect 1000 -330 1020 -310
rect 1040 -330 1060 -310
rect 1080 -330 1100 -310
rect 1120 -330 1140 -310
rect 1160 -330 1180 -310
rect 1200 -330 1220 -310
rect 1240 -330 1260 -310
rect 1280 -330 1300 -310
rect 1320 -330 1340 -310
rect 1360 -330 1380 -310
rect 1400 -330 1420 -310
rect 1440 -330 1460 -310
rect -60 -380 -40 -355
rect -20 -380 0 -355
rect 20 -380 40 -355
rect 60 -380 80 -355
rect 1760 -425 1780 -405
rect 1800 -425 1820 -405
rect 1840 -425 1860 -405
rect 1880 -425 1900 -405
rect 1920 -425 1940 -405
rect 1960 -425 1980 -405
rect 2000 -425 2020 -405
rect 2040 -425 2060 -405
rect 2080 -425 2100 -405
rect 2120 -425 2140 -405
rect 2160 -425 2180 -405
rect 2200 -425 2220 -405
rect 2240 -425 2260 -405
rect 2280 -425 2300 -405
rect 2320 -425 2340 -405
rect 2360 -425 2380 -405
rect 2400 -425 2420 -405
rect 2440 -425 2460 -405
rect 2480 -425 2500 -405
rect 2520 -425 2540 -405
rect -60 -475 -40 -450
rect -20 -475 0 -450
rect 20 -475 40 -450
rect 60 -475 80 -450
rect 680 -520 700 -500
rect 720 -520 740 -500
rect 760 -520 780 -500
rect 800 -520 820 -500
rect 840 -520 860 -500
rect 880 -520 900 -500
rect 920 -520 940 -500
rect 960 -520 980 -500
rect 1000 -520 1020 -500
rect 1040 -520 1060 -500
rect 1080 -520 1100 -500
rect 1120 -520 1140 -500
rect 1160 -520 1180 -500
rect 1200 -520 1220 -500
rect 1240 -520 1260 -500
rect 1280 -520 1300 -500
rect 1320 -520 1340 -500
rect 1360 -520 1380 -500
rect 1400 -520 1420 -500
rect 1440 -520 1460 -500
rect -60 -570 -40 -545
rect -20 -570 0 -545
rect 20 -570 40 -545
rect 60 -570 80 -545
rect 1760 -615 1780 -595
rect 1800 -615 1820 -595
rect 1840 -615 1860 -595
rect 1880 -615 1900 -595
rect 1920 -615 1940 -595
rect 1960 -615 1980 -595
rect 2000 -615 2020 -595
rect 2040 -615 2060 -595
rect 2080 -615 2100 -595
rect 2120 -615 2140 -595
rect 2160 -615 2180 -595
rect 2200 -615 2220 -595
rect 2240 -615 2260 -595
rect 2280 -615 2300 -595
rect 2320 -615 2340 -595
rect 2360 -615 2380 -595
rect 2400 -615 2420 -595
rect 2440 -615 2460 -595
rect 2480 -615 2500 -595
rect 2520 -615 2540 -595
rect -60 -665 -40 -640
rect -20 -665 0 -640
rect 20 -665 40 -640
rect 60 -665 80 -640
rect 680 -710 700 -690
rect 720 -710 740 -690
rect 760 -710 780 -690
rect 800 -710 820 -690
rect 840 -710 860 -690
rect 880 -710 900 -690
rect 920 -710 940 -690
rect 960 -710 980 -690
rect 1000 -710 1020 -690
rect 1040 -710 1060 -690
rect 1080 -710 1100 -690
rect 1120 -710 1140 -690
rect 1160 -710 1180 -690
rect 1200 -710 1220 -690
rect 1240 -710 1260 -690
rect 1280 -710 1300 -690
rect 1320 -710 1340 -690
rect 1360 -710 1380 -690
rect 1400 -710 1420 -690
rect 1440 -710 1460 -690
rect -60 -760 -40 -735
rect -20 -760 0 -735
rect 20 -760 40 -735
rect 60 -760 80 -735
rect 1760 -805 1780 -785
rect 1800 -805 1820 -785
rect 1840 -805 1860 -785
rect 1880 -805 1900 -785
rect 1920 -805 1940 -785
rect 1960 -805 1980 -785
rect 2000 -805 2020 -785
rect 2040 -805 2060 -785
rect 2080 -805 2100 -785
rect 2120 -805 2140 -785
rect 2160 -805 2180 -785
rect 2200 -805 2220 -785
rect 2240 -805 2260 -785
rect 2280 -805 2300 -785
rect 2320 -805 2340 -785
rect 2360 -805 2380 -785
rect 2400 -805 2420 -785
rect 2440 -805 2460 -785
rect 2480 -805 2500 -785
rect 2520 -805 2540 -785
rect -60 -855 -40 -830
rect -20 -855 0 -830
rect 20 -855 40 -830
rect 60 -855 80 -830
rect 680 -900 700 -880
rect 720 -900 740 -880
rect 760 -900 780 -880
rect 800 -900 820 -880
rect 840 -900 860 -880
rect 880 -900 900 -880
rect 920 -900 940 -880
rect 960 -900 980 -880
rect 1000 -900 1020 -880
rect 1040 -900 1060 -880
rect 1080 -900 1100 -880
rect 1120 -900 1140 -880
rect 1160 -900 1180 -880
rect 1200 -900 1220 -880
rect 1240 -900 1260 -880
rect 1280 -900 1300 -880
rect 1320 -900 1340 -880
rect 1360 -900 1380 -880
rect 1400 -900 1420 -880
rect 1440 -900 1460 -880
rect -60 -950 -40 -925
rect -20 -950 0 -925
rect 20 -950 40 -925
rect 60 -950 80 -925
rect 1760 -995 1780 -975
rect 1800 -995 1820 -975
rect 1840 -995 1860 -975
rect 1880 -995 1900 -975
rect 1920 -995 1940 -975
rect 1960 -995 1980 -975
rect 2000 -995 2020 -975
rect 2040 -995 2060 -975
rect 2080 -995 2100 -975
rect 2120 -995 2140 -975
rect 2160 -995 2180 -975
rect 2200 -995 2220 -975
rect 2240 -995 2260 -975
rect 2280 -995 2300 -975
rect 2320 -995 2340 -975
rect 2360 -995 2380 -975
rect 2400 -995 2420 -975
rect 2440 -995 2460 -975
rect 2480 -995 2500 -975
rect 2520 -995 2540 -975
rect -60 -1045 -40 -1020
rect -20 -1045 0 -1020
rect 20 -1045 40 -1020
rect 60 -1045 80 -1020
rect 680 -1090 700 -1070
rect 720 -1090 740 -1070
rect 760 -1090 780 -1070
rect 800 -1090 820 -1070
rect 840 -1090 860 -1070
rect 880 -1090 900 -1070
rect 920 -1090 940 -1070
rect 960 -1090 980 -1070
rect 1000 -1090 1020 -1070
rect 1040 -1090 1060 -1070
rect 1080 -1090 1100 -1070
rect 1120 -1090 1140 -1070
rect 1160 -1090 1180 -1070
rect 1200 -1090 1220 -1070
rect 1240 -1090 1260 -1070
rect 1280 -1090 1300 -1070
rect 1320 -1090 1340 -1070
rect 1360 -1090 1380 -1070
rect 1400 -1090 1420 -1070
rect 1440 -1090 1460 -1070
rect -60 -1140 -40 -1115
rect -20 -1140 0 -1115
rect 20 -1140 40 -1115
rect 60 -1140 80 -1115
rect 1760 -1185 1780 -1165
rect 1800 -1185 1820 -1165
rect 1840 -1185 1860 -1165
rect 1880 -1185 1900 -1165
rect 1920 -1185 1940 -1165
rect 1960 -1185 1980 -1165
rect 2000 -1185 2020 -1165
rect 2040 -1185 2060 -1165
rect 2080 -1185 2100 -1165
rect 2120 -1185 2140 -1165
rect 2160 -1185 2180 -1165
rect 2200 -1185 2220 -1165
rect 2240 -1185 2260 -1165
rect 2280 -1185 2300 -1165
rect 2320 -1185 2340 -1165
rect 2360 -1185 2380 -1165
rect 2400 -1185 2420 -1165
rect 2440 -1185 2460 -1165
rect 2480 -1185 2500 -1165
rect 2520 -1185 2540 -1165
rect -60 -1235 -40 -1210
rect -20 -1235 0 -1210
rect 20 -1235 40 -1210
rect 60 -1235 80 -1210
rect 680 -1280 700 -1260
rect 720 -1280 740 -1260
rect 760 -1280 780 -1260
rect 800 -1280 820 -1260
rect 840 -1280 860 -1260
rect 880 -1280 900 -1260
rect 920 -1280 940 -1260
rect 960 -1280 980 -1260
rect 1000 -1280 1020 -1260
rect 1040 -1280 1060 -1260
rect 1080 -1280 1100 -1260
rect 1120 -1280 1140 -1260
rect 1160 -1280 1180 -1260
rect 1200 -1280 1220 -1260
rect 1240 -1280 1260 -1260
rect 1280 -1280 1300 -1260
rect 1320 -1280 1340 -1260
rect 1360 -1280 1380 -1260
rect 1400 -1280 1420 -1260
rect 1440 -1280 1460 -1260
rect -60 -1330 -40 -1305
rect -20 -1330 0 -1305
rect 20 -1330 40 -1305
rect 60 -1330 80 -1305
rect 1760 -1375 1780 -1355
rect 1800 -1375 1820 -1355
rect 1840 -1375 1860 -1355
rect 1880 -1375 1900 -1355
rect 1920 -1375 1940 -1355
rect 1960 -1375 1980 -1355
rect 2000 -1375 2020 -1355
rect 2040 -1375 2060 -1355
rect 2080 -1375 2100 -1355
rect 2120 -1375 2140 -1355
rect 2160 -1375 2180 -1355
rect 2200 -1375 2220 -1355
rect 2240 -1375 2260 -1355
rect 2280 -1375 2300 -1355
rect 2320 -1375 2340 -1355
rect 2360 -1375 2380 -1355
rect 2400 -1375 2420 -1355
rect 2440 -1375 2460 -1355
rect 2480 -1375 2500 -1355
rect 2520 -1375 2540 -1355
rect -60 -1425 -40 -1400
rect -20 -1425 0 -1400
rect 20 -1425 40 -1400
rect 60 -1425 80 -1400
rect 680 -1470 700 -1450
rect 720 -1470 740 -1450
rect 760 -1470 780 -1450
rect 800 -1470 820 -1450
rect 840 -1470 860 -1450
rect 880 -1470 900 -1450
rect 920 -1470 940 -1450
rect 960 -1470 980 -1450
rect 1000 -1470 1020 -1450
rect 1040 -1470 1060 -1450
rect 1080 -1470 1100 -1450
rect 1120 -1470 1140 -1450
rect 1160 -1470 1180 -1450
rect 1200 -1470 1220 -1450
rect 1240 -1470 1260 -1450
rect 1280 -1470 1300 -1450
rect 1320 -1470 1340 -1450
rect 1360 -1470 1380 -1450
rect 1400 -1470 1420 -1450
rect 1440 -1470 1460 -1450
rect -60 -1520 -40 -1495
rect -20 -1520 0 -1495
rect 20 -1520 40 -1495
rect 60 -1520 80 -1495
rect 1760 -1565 1780 -1545
rect 1800 -1565 1820 -1545
rect 1840 -1565 1860 -1545
rect 1880 -1565 1900 -1545
rect 1920 -1565 1940 -1545
rect 1960 -1565 1980 -1545
rect 2000 -1565 2020 -1545
rect 2040 -1565 2060 -1545
rect 2080 -1565 2100 -1545
rect 2120 -1565 2140 -1545
rect 2160 -1565 2180 -1545
rect 2200 -1565 2220 -1545
rect 2240 -1565 2260 -1545
rect 2280 -1565 2300 -1545
rect 2320 -1565 2340 -1545
rect 2360 -1565 2380 -1545
rect 2400 -1565 2420 -1545
rect 2440 -1565 2460 -1545
rect 2480 -1565 2500 -1545
rect 2520 -1565 2540 -1545
rect -60 -1615 -40 -1590
rect -20 -1615 0 -1590
rect 20 -1615 40 -1590
rect 60 -1615 80 -1590
rect 680 -1660 700 -1640
rect 720 -1660 740 -1640
rect 760 -1660 780 -1640
rect 800 -1660 820 -1640
rect 840 -1660 860 -1640
rect 880 -1660 900 -1640
rect 920 -1660 940 -1640
rect 960 -1660 980 -1640
rect 1000 -1660 1020 -1640
rect 1040 -1660 1060 -1640
rect 1080 -1660 1100 -1640
rect 1120 -1660 1140 -1640
rect 1160 -1660 1180 -1640
rect 1200 -1660 1220 -1640
rect 1240 -1660 1260 -1640
rect 1280 -1660 1300 -1640
rect 1320 -1660 1340 -1640
rect 1360 -1660 1380 -1640
rect 1400 -1660 1420 -1640
rect 1440 -1660 1460 -1640
rect -60 -1710 -40 -1685
rect -20 -1710 0 -1685
rect 20 -1710 40 -1685
rect 60 -1710 80 -1685
rect 1760 -1755 1780 -1735
rect 1800 -1755 1820 -1735
rect 1840 -1755 1860 -1735
rect 1880 -1755 1900 -1735
rect 1920 -1755 1940 -1735
rect 1960 -1755 1980 -1735
rect 2000 -1755 2020 -1735
rect 2040 -1755 2060 -1735
rect 2080 -1755 2100 -1735
rect 2120 -1755 2140 -1735
rect 2160 -1755 2180 -1735
rect 2200 -1755 2220 -1735
rect 2240 -1755 2260 -1735
rect 2280 -1755 2300 -1735
rect 2320 -1755 2340 -1735
rect 2360 -1755 2380 -1735
rect 2400 -1755 2420 -1735
rect 2440 -1755 2460 -1735
rect 2480 -1755 2500 -1735
rect 2520 -1755 2540 -1735
rect -60 -1805 -40 -1780
rect -20 -1805 0 -1780
rect 20 -1805 40 -1780
rect 60 -1805 80 -1780
rect 680 -1850 700 -1830
rect 720 -1850 740 -1830
rect 760 -1850 780 -1830
rect 800 -1850 820 -1830
rect 840 -1850 860 -1830
rect 880 -1850 900 -1830
rect 920 -1850 940 -1830
rect 960 -1850 980 -1830
rect 1000 -1850 1020 -1830
rect 1040 -1850 1060 -1830
rect 1080 -1850 1100 -1830
rect 1120 -1850 1140 -1830
rect 1160 -1850 1180 -1830
rect 1200 -1850 1220 -1830
rect 1240 -1850 1260 -1830
rect 1280 -1850 1300 -1830
rect 1320 -1850 1340 -1830
rect 1360 -1850 1380 -1830
rect 1400 -1850 1420 -1830
rect 1440 -1850 1460 -1830
rect -60 -1900 -40 -1875
rect -20 -1900 0 -1875
rect 20 -1900 40 -1875
rect 60 -1900 80 -1875
rect 1760 -1945 1780 -1925
rect 1800 -1945 1820 -1925
rect 1840 -1945 1860 -1925
rect 1880 -1945 1900 -1925
rect 1920 -1945 1940 -1925
rect 1960 -1945 1980 -1925
rect 2000 -1945 2020 -1925
rect 2040 -1945 2060 -1925
rect 2080 -1945 2100 -1925
rect 2120 -1945 2140 -1925
rect 2160 -1945 2180 -1925
rect 2200 -1945 2220 -1925
rect 2240 -1945 2260 -1925
rect 2280 -1945 2300 -1925
rect 2320 -1945 2340 -1925
rect 2360 -1945 2380 -1925
rect 2400 -1945 2420 -1925
rect 2440 -1945 2460 -1925
rect 2480 -1945 2500 -1925
rect 2520 -1945 2540 -1925
rect -60 -1995 -40 -1970
rect -20 -1995 0 -1970
rect 20 -1995 40 -1970
rect 60 -1995 80 -1970
rect 680 -2040 700 -2020
rect 720 -2040 740 -2020
rect 760 -2040 780 -2020
rect 800 -2040 820 -2020
rect 840 -2040 860 -2020
rect 880 -2040 900 -2020
rect 920 -2040 940 -2020
rect 960 -2040 980 -2020
rect 1000 -2040 1020 -2020
rect 1040 -2040 1060 -2020
rect 1080 -2040 1100 -2020
rect 1120 -2040 1140 -2020
rect 1160 -2040 1180 -2020
rect 1200 -2040 1220 -2020
rect 1240 -2040 1260 -2020
rect 1280 -2040 1300 -2020
rect 1320 -2040 1340 -2020
rect 1360 -2040 1380 -2020
rect 1400 -2040 1420 -2020
rect 1440 -2040 1460 -2020
rect -60 -2090 -40 -2065
rect -20 -2090 0 -2065
rect 20 -2090 40 -2065
rect 60 -2090 80 -2065
rect 1760 -2135 1780 -2115
rect 1800 -2135 1820 -2115
rect 1840 -2135 1860 -2115
rect 1880 -2135 1900 -2115
rect 1920 -2135 1940 -2115
rect 1960 -2135 1980 -2115
rect 2000 -2135 2020 -2115
rect 2040 -2135 2060 -2115
rect 2080 -2135 2100 -2115
rect 2120 -2135 2140 -2115
rect 2160 -2135 2180 -2115
rect 2200 -2135 2220 -2115
rect 2240 -2135 2260 -2115
rect 2280 -2135 2300 -2115
rect 2320 -2135 2340 -2115
rect 2360 -2135 2380 -2115
rect 2400 -2135 2420 -2115
rect 2440 -2135 2460 -2115
rect 2480 -2135 2500 -2115
rect 2520 -2135 2540 -2115
rect -60 -2185 -40 -2160
rect -20 -2185 0 -2160
rect 20 -2185 40 -2160
rect 60 -2185 80 -2160
rect 680 -2230 700 -2210
rect 720 -2230 740 -2210
rect 760 -2230 780 -2210
rect 800 -2230 820 -2210
rect 840 -2230 860 -2210
rect 880 -2230 900 -2210
rect 920 -2230 940 -2210
rect 960 -2230 980 -2210
rect 1000 -2230 1020 -2210
rect 1040 -2230 1060 -2210
rect 1080 -2230 1100 -2210
rect 1120 -2230 1140 -2210
rect 1160 -2230 1180 -2210
rect 1200 -2230 1220 -2210
rect 1240 -2230 1260 -2210
rect 1280 -2230 1300 -2210
rect 1320 -2230 1340 -2210
rect 1360 -2230 1380 -2210
rect 1400 -2230 1420 -2210
rect 1440 -2230 1460 -2210
rect -60 -2280 -40 -2255
rect -20 -2280 0 -2255
rect 20 -2280 40 -2255
rect 60 -2280 80 -2255
rect 1760 -2325 1780 -2305
rect 1800 -2325 1820 -2305
rect 1840 -2325 1860 -2305
rect 1880 -2325 1900 -2305
rect 1920 -2325 1940 -2305
rect 1960 -2325 1980 -2305
rect 2000 -2325 2020 -2305
rect 2040 -2325 2060 -2305
rect 2080 -2325 2100 -2305
rect 2120 -2325 2140 -2305
rect 2160 -2325 2180 -2305
rect 2200 -2325 2220 -2305
rect 2240 -2325 2260 -2305
rect 2280 -2325 2300 -2305
rect 2320 -2325 2340 -2305
rect 2360 -2325 2380 -2305
rect 2400 -2325 2420 -2305
rect 2440 -2325 2460 -2305
rect 2480 -2325 2500 -2305
rect 2520 -2325 2540 -2305
rect -60 -2375 -40 -2350
rect -20 -2375 0 -2350
rect 20 -2375 40 -2350
rect 60 -2375 80 -2350
rect 680 -2420 700 -2400
rect 720 -2420 740 -2400
rect 760 -2420 780 -2400
rect 800 -2420 820 -2400
rect 840 -2420 860 -2400
rect 880 -2420 900 -2400
rect 920 -2420 940 -2400
rect 960 -2420 980 -2400
rect 1000 -2420 1020 -2400
rect 1040 -2420 1060 -2400
rect 1080 -2420 1100 -2400
rect 1120 -2420 1140 -2400
rect 1160 -2420 1180 -2400
rect 1200 -2420 1220 -2400
rect 1240 -2420 1260 -2400
rect 1280 -2420 1300 -2400
rect 1320 -2420 1340 -2400
rect 1360 -2420 1380 -2400
rect 1400 -2420 1420 -2400
rect 1440 -2420 1460 -2400
rect -60 -2470 -40 -2445
rect -20 -2470 0 -2445
rect 20 -2470 40 -2445
rect 60 -2470 80 -2445
rect 1760 -2515 1780 -2495
rect 1800 -2515 1820 -2495
rect 1840 -2515 1860 -2495
rect 1880 -2515 1900 -2495
rect 1920 -2515 1940 -2495
rect 1960 -2515 1980 -2495
rect 2000 -2515 2020 -2495
rect 2040 -2515 2060 -2495
rect 2080 -2515 2100 -2495
rect 2120 -2515 2140 -2495
rect 2160 -2515 2180 -2495
rect 2200 -2515 2220 -2495
rect 2240 -2515 2260 -2495
rect 2280 -2515 2300 -2495
rect 2320 -2515 2340 -2495
rect 2360 -2515 2380 -2495
rect 2400 -2515 2420 -2495
rect 2440 -2515 2460 -2495
rect 2480 -2515 2500 -2495
rect 2520 -2515 2540 -2495
rect -60 -2565 -40 -2540
rect -20 -2565 0 -2540
rect 20 -2565 40 -2540
rect 60 -2565 80 -2540
rect 680 -2610 700 -2590
rect 720 -2610 740 -2590
rect 760 -2610 780 -2590
rect 800 -2610 820 -2590
rect 840 -2610 860 -2590
rect 880 -2610 900 -2590
rect 920 -2610 940 -2590
rect 960 -2610 980 -2590
rect 1000 -2610 1020 -2590
rect 1040 -2610 1060 -2590
rect 1080 -2610 1100 -2590
rect 1120 -2610 1140 -2590
rect 1160 -2610 1180 -2590
rect 1200 -2610 1220 -2590
rect 1240 -2610 1260 -2590
rect 1280 -2610 1300 -2590
rect 1320 -2610 1340 -2590
rect 1360 -2610 1380 -2590
rect 1400 -2610 1420 -2590
rect 1440 -2610 1460 -2590
rect -60 -2660 -40 -2635
rect -20 -2660 0 -2635
rect 20 -2660 40 -2635
rect 60 -2660 80 -2635
rect 1760 -2705 1780 -2685
rect 1800 -2705 1820 -2685
rect 1840 -2705 1860 -2685
rect 1880 -2705 1900 -2685
rect 1920 -2705 1940 -2685
rect 1960 -2705 1980 -2685
rect 2000 -2705 2020 -2685
rect 2040 -2705 2060 -2685
rect 2080 -2705 2100 -2685
rect 2120 -2705 2140 -2685
rect 2160 -2705 2180 -2685
rect 2200 -2705 2220 -2685
rect 2240 -2705 2260 -2685
rect 2280 -2705 2300 -2685
rect 2320 -2705 2340 -2685
rect 2360 -2705 2380 -2685
rect 2400 -2705 2420 -2685
rect 2440 -2705 2460 -2685
rect 2480 -2705 2500 -2685
rect 2520 -2705 2540 -2685
rect 1760 -2745 1780 -2725
rect 1800 -2745 1820 -2725
rect 1840 -2745 1860 -2725
rect 1880 -2745 1900 -2725
rect 1920 -2745 1940 -2725
rect 1960 -2745 1980 -2725
rect 2000 -2745 2020 -2725
rect 2040 -2745 2060 -2725
rect 2080 -2745 2100 -2725
rect 2120 -2745 2140 -2725
rect 2160 -2745 2180 -2725
rect 2200 -2745 2220 -2725
rect 2240 -2745 2260 -2725
rect 2280 -2745 2300 -2725
rect 2320 -2745 2340 -2725
rect 2360 -2745 2380 -2725
rect 2400 -2745 2420 -2725
rect 2440 -2745 2460 -2725
rect 2480 -2745 2500 -2725
rect 2520 -2745 2540 -2725
<< metal1 >>
rect 1750 2345 2550 2385
rect 670 2325 1470 2345
rect 1750 2325 1780 2345
rect 1800 2325 1820 2345
rect 1840 2325 1860 2345
rect 1880 2325 1900 2345
rect 1920 2325 1940 2345
rect 1960 2325 1980 2345
rect 2000 2325 2020 2345
rect 2040 2325 2060 2345
rect 2080 2325 2100 2345
rect 2120 2325 2140 2345
rect 2160 2325 2180 2345
rect 2200 2325 2220 2345
rect 2240 2325 2260 2345
rect 2280 2325 2300 2345
rect 2320 2325 2340 2345
rect 2360 2325 2380 2345
rect 2400 2325 2420 2345
rect 2440 2325 2460 2345
rect 2480 2325 2500 2345
rect 2520 2325 2550 2345
rect 670 2260 1470 2270
rect 670 2240 680 2260
rect 700 2240 720 2260
rect 740 2240 760 2260
rect 780 2240 800 2260
rect 820 2240 840 2260
rect 860 2240 880 2260
rect 900 2240 920 2260
rect 940 2240 960 2260
rect 980 2240 1000 2260
rect 1020 2240 1040 2260
rect 1060 2240 1080 2260
rect 1100 2240 1120 2260
rect 1140 2240 1160 2260
rect 1180 2240 1200 2260
rect 1220 2240 1240 2260
rect 1260 2240 1280 2260
rect 1300 2240 1320 2260
rect 1340 2240 1360 2260
rect 1380 2240 1400 2260
rect 1420 2240 1440 2260
rect 1460 2240 1470 2260
rect 670 2217 1470 2240
rect 670 2197 680 2217
rect 700 2197 720 2217
rect 740 2197 760 2217
rect 780 2197 800 2217
rect 820 2197 840 2217
rect 860 2197 880 2217
rect 900 2197 920 2217
rect 940 2197 960 2217
rect 980 2197 1000 2217
rect 1020 2197 1040 2217
rect 1060 2197 1080 2217
rect 1100 2197 1120 2217
rect 1140 2197 1160 2217
rect 1180 2197 1200 2217
rect 1220 2197 1240 2217
rect 1260 2197 1280 2217
rect 1300 2197 1320 2217
rect 1340 2197 1360 2217
rect 1380 2197 1400 2217
rect 1420 2197 1440 2217
rect 1460 2197 1470 2217
rect 0 2175 165 2185
rect 0 2155 10 2175
rect 30 2155 50 2175
rect 70 2155 90 2175
rect 110 2155 130 2175
rect 150 2155 165 2175
rect 0 2095 165 2155
rect 0 2075 10 2095
rect 30 2075 50 2095
rect 70 2075 90 2095
rect 110 2075 130 2095
rect 150 2075 165 2095
rect 0 2010 165 2075
rect 0 1990 10 2010
rect 30 1990 50 2010
rect 70 1990 90 2010
rect 110 1990 130 2010
rect 150 1990 165 2010
rect 0 1930 165 1990
rect 0 1910 10 1930
rect 30 1910 50 1930
rect 70 1910 90 1930
rect 110 1910 130 1930
rect 150 1910 165 1930
rect 0 1850 165 1910
rect 0 1830 10 1850
rect 30 1830 50 1850
rect 70 1830 90 1850
rect 110 1830 130 1850
rect 150 1830 165 1850
rect 0 1765 165 1830
rect 0 1745 10 1765
rect 30 1745 50 1765
rect 70 1745 90 1765
rect 110 1745 130 1765
rect 150 1745 165 1765
rect 0 1685 165 1745
rect 0 1665 10 1685
rect 30 1665 50 1685
rect 70 1665 90 1685
rect 110 1665 130 1685
rect 150 1665 165 1685
rect 0 1600 165 1665
rect 0 1580 10 1600
rect 30 1580 50 1600
rect 70 1580 90 1600
rect 110 1580 130 1600
rect 150 1580 165 1600
rect 0 1520 165 1580
rect 0 1500 10 1520
rect 30 1500 50 1520
rect 70 1500 90 1520
rect 110 1500 130 1520
rect 150 1500 165 1520
rect 0 1440 165 1500
rect 0 1420 10 1440
rect 30 1420 50 1440
rect 70 1420 90 1440
rect 110 1420 130 1440
rect 150 1420 165 1440
rect 0 1355 165 1420
rect 0 1335 10 1355
rect 30 1335 50 1355
rect 70 1335 90 1355
rect 110 1335 130 1355
rect 150 1335 165 1355
rect 0 1275 165 1335
rect 0 1255 10 1275
rect 30 1255 50 1275
rect 70 1255 90 1275
rect 110 1255 130 1275
rect 150 1255 165 1275
rect 0 1190 165 1255
rect 0 1170 10 1190
rect 30 1170 50 1190
rect 70 1170 90 1190
rect 110 1170 130 1190
rect 150 1170 165 1190
rect 0 1110 165 1170
rect 0 1090 10 1110
rect 30 1090 50 1110
rect 70 1090 90 1110
rect 110 1090 130 1110
rect 150 1090 165 1110
rect 0 1030 165 1090
rect 0 1010 10 1030
rect 30 1010 50 1030
rect 70 1010 90 1030
rect 110 1010 130 1030
rect 150 1010 165 1030
rect 0 945 165 1010
rect 0 925 10 945
rect 30 925 50 945
rect 70 925 90 945
rect 110 925 130 945
rect 150 925 165 945
rect 0 865 165 925
rect 0 845 10 865
rect 30 845 50 865
rect 70 845 90 865
rect 110 845 130 865
rect 150 845 165 865
rect 0 780 165 845
rect 0 760 10 780
rect 30 760 50 780
rect 70 760 90 780
rect 110 760 130 780
rect 150 760 165 780
rect 0 700 165 760
rect 0 680 10 700
rect 30 680 50 700
rect 70 680 90 700
rect 110 680 130 700
rect 150 680 165 700
rect 0 620 165 680
rect 0 600 10 620
rect 30 600 50 620
rect 70 600 90 620
rect 110 600 130 620
rect 150 600 165 620
rect 0 535 165 600
rect 0 515 10 535
rect 30 515 50 535
rect 70 515 90 535
rect 110 515 130 535
rect 150 515 165 535
rect 0 455 165 515
rect 0 435 10 455
rect 30 435 50 455
rect 70 435 90 455
rect 110 435 130 455
rect 150 435 165 455
rect 0 375 165 435
rect 0 355 10 375
rect 30 355 50 375
rect 70 355 90 375
rect 110 355 130 375
rect 150 355 165 375
rect 0 290 165 355
rect 0 270 10 290
rect 30 270 50 290
rect 70 270 90 290
rect 110 270 130 290
rect 150 270 165 290
rect 0 210 165 270
rect 0 190 10 210
rect 30 190 50 210
rect 70 190 90 210
rect 110 190 130 210
rect 150 190 165 210
rect 0 130 165 190
rect 0 110 10 130
rect 30 110 50 130
rect 70 110 90 130
rect 110 110 130 130
rect 150 110 165 130
rect 0 100 165 110
rect 670 2053 1470 2197
rect 670 2033 680 2053
rect 700 2033 720 2053
rect 740 2033 760 2053
rect 780 2033 800 2053
rect 820 2033 840 2053
rect 860 2033 880 2053
rect 900 2033 920 2053
rect 940 2033 960 2053
rect 980 2033 1000 2053
rect 1020 2033 1040 2053
rect 1060 2033 1080 2053
rect 1100 2033 1120 2053
rect 1140 2033 1160 2053
rect 1180 2033 1200 2053
rect 1220 2033 1240 2053
rect 1260 2033 1280 2053
rect 1300 2033 1320 2053
rect 1340 2033 1360 2053
rect 1380 2033 1400 2053
rect 1420 2033 1440 2053
rect 1460 2033 1470 2053
rect 670 1889 1470 2033
rect 670 1869 680 1889
rect 700 1869 720 1889
rect 740 1869 760 1889
rect 780 1869 800 1889
rect 820 1869 840 1889
rect 860 1869 880 1889
rect 900 1869 920 1889
rect 940 1869 960 1889
rect 980 1869 1000 1889
rect 1020 1869 1040 1889
rect 1060 1869 1080 1889
rect 1100 1869 1120 1889
rect 1140 1869 1160 1889
rect 1180 1869 1200 1889
rect 1220 1869 1240 1889
rect 1260 1869 1280 1889
rect 1300 1869 1320 1889
rect 1340 1869 1360 1889
rect 1380 1869 1400 1889
rect 1420 1869 1440 1889
rect 1460 1869 1470 1889
rect 670 1725 1470 1869
rect 670 1705 680 1725
rect 700 1705 720 1725
rect 740 1705 760 1725
rect 780 1705 800 1725
rect 820 1705 840 1725
rect 860 1705 880 1725
rect 900 1705 920 1725
rect 940 1705 960 1725
rect 980 1705 1000 1725
rect 1020 1705 1040 1725
rect 1060 1705 1080 1725
rect 1100 1705 1120 1725
rect 1140 1705 1160 1725
rect 1180 1705 1200 1725
rect 1220 1705 1240 1725
rect 1260 1705 1280 1725
rect 1300 1705 1320 1725
rect 1340 1705 1360 1725
rect 1380 1705 1400 1725
rect 1420 1705 1440 1725
rect 1460 1705 1470 1725
rect 670 1561 1470 1705
rect 670 1541 680 1561
rect 700 1541 720 1561
rect 740 1541 760 1561
rect 780 1541 800 1561
rect 820 1541 840 1561
rect 860 1541 880 1561
rect 900 1541 920 1561
rect 940 1541 960 1561
rect 980 1541 1000 1561
rect 1020 1541 1040 1561
rect 1060 1541 1080 1561
rect 1100 1541 1120 1561
rect 1140 1541 1160 1561
rect 1180 1541 1200 1561
rect 1220 1541 1240 1561
rect 1260 1541 1280 1561
rect 1300 1541 1320 1561
rect 1340 1541 1360 1561
rect 1380 1541 1400 1561
rect 1420 1541 1440 1561
rect 1460 1541 1470 1561
rect 670 1397 1470 1541
rect 670 1377 680 1397
rect 700 1377 720 1397
rect 740 1377 760 1397
rect 780 1377 800 1397
rect 820 1377 840 1397
rect 860 1377 880 1397
rect 900 1377 920 1397
rect 940 1377 960 1397
rect 980 1377 1000 1397
rect 1020 1377 1040 1397
rect 1060 1377 1080 1397
rect 1100 1377 1120 1397
rect 1140 1377 1160 1397
rect 1180 1377 1200 1397
rect 1220 1377 1240 1397
rect 1260 1377 1280 1397
rect 1300 1377 1320 1397
rect 1340 1377 1360 1397
rect 1380 1377 1400 1397
rect 1420 1377 1440 1397
rect 1460 1377 1470 1397
rect 670 1233 1470 1377
rect 670 1213 680 1233
rect 700 1213 720 1233
rect 740 1213 760 1233
rect 780 1213 800 1233
rect 820 1213 840 1233
rect 860 1213 880 1233
rect 900 1213 920 1233
rect 940 1213 960 1233
rect 980 1213 1000 1233
rect 1020 1213 1040 1233
rect 1060 1213 1080 1233
rect 1100 1213 1120 1233
rect 1140 1213 1160 1233
rect 1180 1213 1200 1233
rect 1220 1213 1240 1233
rect 1260 1213 1280 1233
rect 1300 1213 1320 1233
rect 1340 1213 1360 1233
rect 1380 1213 1400 1233
rect 1420 1213 1440 1233
rect 1460 1213 1470 1233
rect 670 1069 1470 1213
rect 670 1049 680 1069
rect 700 1049 720 1069
rect 740 1049 760 1069
rect 780 1049 800 1069
rect 820 1049 840 1069
rect 860 1049 880 1069
rect 900 1049 920 1069
rect 940 1049 960 1069
rect 980 1049 1000 1069
rect 1020 1049 1040 1069
rect 1060 1049 1080 1069
rect 1100 1049 1120 1069
rect 1140 1049 1160 1069
rect 1180 1049 1200 1069
rect 1220 1049 1240 1069
rect 1260 1049 1280 1069
rect 1300 1049 1320 1069
rect 1340 1049 1360 1069
rect 1380 1049 1400 1069
rect 1420 1049 1440 1069
rect 1460 1049 1470 1069
rect 670 905 1470 1049
rect 670 885 680 905
rect 700 885 720 905
rect 740 885 760 905
rect 780 885 800 905
rect 820 885 840 905
rect 860 885 880 905
rect 900 885 920 905
rect 940 885 960 905
rect 980 885 1000 905
rect 1020 885 1040 905
rect 1060 885 1080 905
rect 1100 885 1120 905
rect 1140 885 1160 905
rect 1180 885 1200 905
rect 1220 885 1240 905
rect 1260 885 1280 905
rect 1300 885 1320 905
rect 1340 885 1360 905
rect 1380 885 1400 905
rect 1420 885 1440 905
rect 1460 885 1470 905
rect 670 741 1470 885
rect 670 721 680 741
rect 700 721 720 741
rect 740 721 760 741
rect 780 721 800 741
rect 820 721 840 741
rect 860 721 880 741
rect 900 721 920 741
rect 940 721 960 741
rect 980 721 1000 741
rect 1020 721 1040 741
rect 1060 721 1080 741
rect 1100 721 1120 741
rect 1140 721 1160 741
rect 1180 721 1200 741
rect 1220 721 1240 741
rect 1260 721 1280 741
rect 1300 721 1320 741
rect 1340 721 1360 741
rect 1380 721 1400 741
rect 1420 721 1440 741
rect 1460 721 1470 741
rect 670 577 1470 721
rect 670 557 680 577
rect 700 557 720 577
rect 740 557 760 577
rect 780 557 800 577
rect 820 557 840 577
rect 860 557 880 577
rect 900 557 920 577
rect 940 557 960 577
rect 980 557 1000 577
rect 1020 557 1040 577
rect 1060 557 1080 577
rect 1100 557 1120 577
rect 1140 557 1160 577
rect 1180 557 1200 577
rect 1220 557 1240 577
rect 1260 557 1280 577
rect 1300 557 1320 577
rect 1340 557 1360 577
rect 1380 557 1400 577
rect 1420 557 1440 577
rect 1460 557 1470 577
rect 670 413 1470 557
rect 670 393 680 413
rect 700 393 720 413
rect 740 393 760 413
rect 780 393 800 413
rect 820 393 840 413
rect 860 393 880 413
rect 900 393 920 413
rect 940 393 960 413
rect 980 393 1000 413
rect 1020 393 1040 413
rect 1060 393 1080 413
rect 1100 393 1120 413
rect 1140 393 1160 413
rect 1180 393 1200 413
rect 1220 393 1240 413
rect 1260 393 1280 413
rect 1300 393 1320 413
rect 1340 393 1360 413
rect 1380 393 1400 413
rect 1420 393 1440 413
rect 1460 393 1470 413
rect 670 249 1470 393
rect 670 229 680 249
rect 700 229 720 249
rect 740 229 760 249
rect 780 229 800 249
rect 820 229 840 249
rect 860 229 880 249
rect 900 229 920 249
rect 940 229 960 249
rect 980 229 1000 249
rect 1020 229 1040 249
rect 1060 229 1080 249
rect 1100 229 1120 249
rect 1140 229 1160 249
rect 1180 229 1200 249
rect 1220 229 1240 249
rect 1260 229 1280 249
rect 1300 229 1320 249
rect 1340 229 1360 249
rect 1380 229 1400 249
rect 1420 229 1440 249
rect 1460 229 1470 249
rect 670 85 1470 229
rect 670 65 680 85
rect 700 65 720 85
rect 740 65 760 85
rect 780 65 800 85
rect 820 65 840 85
rect 860 65 880 85
rect 900 65 920 85
rect 940 65 960 85
rect 980 65 1000 85
rect 1020 65 1040 85
rect 1060 65 1080 85
rect 1100 65 1120 85
rect 1140 65 1160 85
rect 1180 65 1200 85
rect 1220 65 1240 85
rect 1260 65 1280 85
rect 1300 65 1320 85
rect 1340 65 1360 85
rect 1380 65 1400 85
rect 1420 65 1440 85
rect 1460 65 1470 85
rect 670 45 1470 65
rect 670 25 680 45
rect 700 25 720 45
rect 740 25 760 45
rect 780 25 800 45
rect 820 25 840 45
rect 860 25 880 45
rect 900 25 920 45
rect 940 25 960 45
rect 980 25 1000 45
rect 1020 25 1040 45
rect 1060 25 1080 45
rect 1100 25 1120 45
rect 1140 25 1160 45
rect 1180 25 1200 45
rect 1220 25 1240 45
rect 1260 25 1280 45
rect 1300 25 1320 45
rect 1340 25 1360 45
rect 1380 25 1400 45
rect 1420 25 1440 45
rect 1460 25 1470 45
rect -70 -260 85 -250
rect -70 -285 -60 -260
rect -40 -285 -20 -260
rect 0 -285 20 -260
rect 40 -285 60 -260
rect 80 -285 85 -260
rect -70 -355 85 -285
rect -70 -380 -60 -355
rect -40 -380 -20 -355
rect 0 -380 20 -355
rect 40 -380 60 -355
rect 80 -380 85 -355
rect -70 -450 85 -380
rect -70 -475 -60 -450
rect -40 -475 -20 -450
rect 0 -475 20 -450
rect 40 -475 60 -450
rect 80 -475 85 -450
rect -70 -545 85 -475
rect -70 -570 -60 -545
rect -40 -570 -20 -545
rect 0 -570 20 -545
rect 40 -570 60 -545
rect 80 -570 85 -545
rect -70 -640 85 -570
rect -70 -665 -60 -640
rect -40 -665 -20 -640
rect 0 -665 20 -640
rect 40 -665 60 -640
rect 80 -665 85 -640
rect -70 -735 85 -665
rect -70 -760 -60 -735
rect -40 -760 -20 -735
rect 0 -760 20 -735
rect 40 -760 60 -735
rect 80 -760 85 -735
rect -70 -830 85 -760
rect -70 -855 -60 -830
rect -40 -855 -20 -830
rect 0 -855 20 -830
rect 40 -855 60 -830
rect 80 -855 85 -830
rect -70 -925 85 -855
rect -70 -950 -60 -925
rect -40 -950 -20 -925
rect 0 -950 20 -925
rect 40 -950 60 -925
rect 80 -950 85 -925
rect -70 -1020 85 -950
rect -70 -1045 -60 -1020
rect -40 -1045 -20 -1020
rect 0 -1045 20 -1020
rect 40 -1045 60 -1020
rect 80 -1045 85 -1020
rect -70 -1115 85 -1045
rect -70 -1140 -60 -1115
rect -40 -1140 -20 -1115
rect 0 -1140 20 -1115
rect 40 -1140 60 -1115
rect 80 -1140 85 -1115
rect -70 -1210 85 -1140
rect -70 -1235 -60 -1210
rect -40 -1235 -20 -1210
rect 0 -1235 20 -1210
rect 40 -1235 60 -1210
rect 80 -1235 85 -1210
rect -70 -1305 85 -1235
rect -70 -1330 -60 -1305
rect -40 -1330 -20 -1305
rect 0 -1330 20 -1305
rect 40 -1330 60 -1305
rect 80 -1330 85 -1305
rect -70 -1400 85 -1330
rect -70 -1425 -60 -1400
rect -40 -1425 -20 -1400
rect 0 -1425 20 -1400
rect 40 -1425 60 -1400
rect 80 -1425 85 -1400
rect -70 -1495 85 -1425
rect -70 -1520 -60 -1495
rect -40 -1520 -20 -1495
rect 0 -1520 20 -1495
rect 40 -1520 60 -1495
rect 80 -1520 85 -1495
rect -70 -1590 85 -1520
rect -70 -1615 -60 -1590
rect -40 -1615 -20 -1590
rect 0 -1615 20 -1590
rect 40 -1615 60 -1590
rect 80 -1615 85 -1590
rect -70 -1685 85 -1615
rect -70 -1710 -60 -1685
rect -40 -1710 -20 -1685
rect 0 -1710 20 -1685
rect 40 -1710 60 -1685
rect 80 -1710 85 -1685
rect -70 -1780 85 -1710
rect -70 -1805 -60 -1780
rect -40 -1805 -20 -1780
rect 0 -1805 20 -1780
rect 40 -1805 60 -1780
rect 80 -1805 85 -1780
rect -70 -1875 85 -1805
rect -70 -1900 -60 -1875
rect -40 -1900 -20 -1875
rect 0 -1900 20 -1875
rect 40 -1900 60 -1875
rect 80 -1900 85 -1875
rect -70 -1970 85 -1900
rect -70 -1995 -60 -1970
rect -40 -1995 -20 -1970
rect 0 -1995 20 -1970
rect 40 -1995 60 -1970
rect 80 -1995 85 -1970
rect -70 -2065 85 -1995
rect -70 -2090 -60 -2065
rect -40 -2090 -20 -2065
rect 0 -2090 20 -2065
rect 40 -2090 60 -2065
rect 80 -2090 85 -2065
rect -70 -2160 85 -2090
rect -70 -2185 -60 -2160
rect -40 -2185 -20 -2160
rect 0 -2185 20 -2160
rect 40 -2185 60 -2160
rect 80 -2185 85 -2160
rect -70 -2255 85 -2185
rect -70 -2280 -60 -2255
rect -40 -2280 -20 -2255
rect 0 -2280 20 -2255
rect 40 -2280 60 -2255
rect 80 -2280 85 -2255
rect -70 -2350 85 -2280
rect -70 -2375 -60 -2350
rect -40 -2375 -20 -2350
rect 0 -2375 20 -2350
rect 40 -2375 60 -2350
rect 80 -2375 85 -2350
rect -70 -2445 85 -2375
rect -70 -2470 -60 -2445
rect -40 -2470 -20 -2445
rect 0 -2470 20 -2445
rect 40 -2470 60 -2445
rect 80 -2470 85 -2445
rect -70 -2540 85 -2470
rect -70 -2565 -60 -2540
rect -40 -2565 -20 -2540
rect 0 -2565 20 -2540
rect 40 -2565 60 -2540
rect 80 -2565 85 -2540
rect -70 -2635 85 -2565
rect 670 -310 1470 25
rect 1750 2135 2550 2325
rect 1750 2115 1760 2135
rect 1780 2115 1800 2135
rect 1820 2115 1840 2135
rect 1860 2115 1880 2135
rect 1900 2115 1920 2135
rect 1940 2115 1960 2135
rect 1980 2115 2000 2135
rect 2020 2115 2040 2135
rect 2060 2115 2080 2135
rect 2100 2115 2120 2135
rect 2140 2115 2160 2135
rect 2180 2115 2200 2135
rect 2220 2115 2240 2135
rect 2260 2115 2280 2135
rect 2300 2115 2320 2135
rect 2340 2115 2360 2135
rect 2380 2115 2400 2135
rect 2420 2115 2440 2135
rect 2460 2115 2480 2135
rect 2500 2115 2520 2135
rect 2540 2115 2550 2135
rect 1750 1971 2550 2115
rect 1750 1951 1760 1971
rect 1780 1951 1800 1971
rect 1820 1951 1840 1971
rect 1860 1951 1880 1971
rect 1900 1951 1920 1971
rect 1940 1951 1960 1971
rect 1980 1951 2000 1971
rect 2020 1951 2040 1971
rect 2060 1951 2080 1971
rect 2100 1951 2120 1971
rect 2140 1951 2160 1971
rect 2180 1951 2200 1971
rect 2220 1951 2240 1971
rect 2260 1951 2280 1971
rect 2300 1951 2320 1971
rect 2340 1951 2360 1971
rect 2380 1951 2400 1971
rect 2420 1951 2440 1971
rect 2460 1951 2480 1971
rect 2500 1951 2520 1971
rect 2540 1951 2550 1971
rect 1750 1807 2550 1951
rect 1750 1787 1760 1807
rect 1780 1787 1800 1807
rect 1820 1787 1840 1807
rect 1860 1787 1880 1807
rect 1900 1787 1920 1807
rect 1940 1787 1960 1807
rect 1980 1787 2000 1807
rect 2020 1787 2040 1807
rect 2060 1787 2080 1807
rect 2100 1787 2120 1807
rect 2140 1787 2160 1807
rect 2180 1787 2200 1807
rect 2220 1787 2240 1807
rect 2260 1787 2280 1807
rect 2300 1787 2320 1807
rect 2340 1787 2360 1807
rect 2380 1787 2400 1807
rect 2420 1787 2440 1807
rect 2460 1787 2480 1807
rect 2500 1787 2520 1807
rect 2540 1787 2550 1807
rect 1750 1643 2550 1787
rect 1750 1623 1760 1643
rect 1780 1623 1800 1643
rect 1820 1623 1840 1643
rect 1860 1623 1880 1643
rect 1900 1623 1920 1643
rect 1940 1623 1960 1643
rect 1980 1623 2000 1643
rect 2020 1623 2040 1643
rect 2060 1623 2080 1643
rect 2100 1623 2120 1643
rect 2140 1623 2160 1643
rect 2180 1623 2200 1643
rect 2220 1623 2240 1643
rect 2260 1623 2280 1643
rect 2300 1623 2320 1643
rect 2340 1623 2360 1643
rect 2380 1623 2400 1643
rect 2420 1623 2440 1643
rect 2460 1623 2480 1643
rect 2500 1623 2520 1643
rect 2540 1623 2550 1643
rect 1750 1479 2550 1623
rect 1750 1459 1760 1479
rect 1780 1459 1800 1479
rect 1820 1459 1840 1479
rect 1860 1459 1880 1479
rect 1900 1459 1920 1479
rect 1940 1459 1960 1479
rect 1980 1459 2000 1479
rect 2020 1459 2040 1479
rect 2060 1459 2080 1479
rect 2100 1459 2120 1479
rect 2140 1459 2160 1479
rect 2180 1459 2200 1479
rect 2220 1459 2240 1479
rect 2260 1459 2280 1479
rect 2300 1459 2320 1479
rect 2340 1459 2360 1479
rect 2380 1459 2400 1479
rect 2420 1459 2440 1479
rect 2460 1459 2480 1479
rect 2500 1459 2520 1479
rect 2540 1459 2550 1479
rect 1750 1315 2550 1459
rect 1750 1295 1760 1315
rect 1780 1295 1800 1315
rect 1820 1295 1840 1315
rect 1860 1295 1880 1315
rect 1900 1295 1920 1315
rect 1940 1295 1960 1315
rect 1980 1295 2000 1315
rect 2020 1295 2040 1315
rect 2060 1295 2080 1315
rect 2100 1295 2120 1315
rect 2140 1295 2160 1315
rect 2180 1295 2200 1315
rect 2220 1295 2240 1315
rect 2260 1295 2280 1315
rect 2300 1295 2320 1315
rect 2340 1295 2360 1315
rect 2380 1295 2400 1315
rect 2420 1295 2440 1315
rect 2460 1295 2480 1315
rect 2500 1295 2520 1315
rect 2540 1295 2550 1315
rect 1750 1151 2550 1295
rect 1750 1131 1760 1151
rect 1780 1131 1800 1151
rect 1820 1131 1840 1151
rect 1860 1131 1880 1151
rect 1900 1131 1920 1151
rect 1940 1131 1960 1151
rect 1980 1131 2000 1151
rect 2020 1131 2040 1151
rect 2060 1131 2080 1151
rect 2100 1131 2120 1151
rect 2140 1131 2160 1151
rect 2180 1131 2200 1151
rect 2220 1131 2240 1151
rect 2260 1131 2280 1151
rect 2300 1131 2320 1151
rect 2340 1131 2360 1151
rect 2380 1131 2400 1151
rect 2420 1131 2440 1151
rect 2460 1131 2480 1151
rect 2500 1131 2520 1151
rect 2540 1131 2550 1151
rect 1750 987 2550 1131
rect 1750 967 1760 987
rect 1780 967 1800 987
rect 1820 967 1840 987
rect 1860 967 1880 987
rect 1900 967 1920 987
rect 1940 967 1960 987
rect 1980 967 2000 987
rect 2020 967 2040 987
rect 2060 967 2080 987
rect 2100 967 2120 987
rect 2140 967 2160 987
rect 2180 967 2200 987
rect 2220 967 2240 987
rect 2260 967 2280 987
rect 2300 967 2320 987
rect 2340 967 2360 987
rect 2380 967 2400 987
rect 2420 967 2440 987
rect 2460 967 2480 987
rect 2500 967 2520 987
rect 2540 967 2550 987
rect 1750 823 2550 967
rect 1750 803 1760 823
rect 1780 803 1800 823
rect 1820 803 1840 823
rect 1860 803 1880 823
rect 1900 803 1920 823
rect 1940 803 1960 823
rect 1980 803 2000 823
rect 2020 803 2040 823
rect 2060 803 2080 823
rect 2100 803 2120 823
rect 2140 803 2160 823
rect 2180 803 2200 823
rect 2220 803 2240 823
rect 2260 803 2280 823
rect 2300 803 2320 823
rect 2340 803 2360 823
rect 2380 803 2400 823
rect 2420 803 2440 823
rect 2460 803 2480 823
rect 2500 803 2520 823
rect 2540 803 2550 823
rect 1750 659 2550 803
rect 1750 639 1760 659
rect 1780 639 1800 659
rect 1820 639 1840 659
rect 1860 639 1880 659
rect 1900 639 1920 659
rect 1940 639 1960 659
rect 1980 639 2000 659
rect 2020 639 2040 659
rect 2060 639 2080 659
rect 2100 639 2120 659
rect 2140 639 2160 659
rect 2180 639 2200 659
rect 2220 639 2240 659
rect 2260 639 2280 659
rect 2300 639 2320 659
rect 2340 639 2360 659
rect 2380 639 2400 659
rect 2420 639 2440 659
rect 2460 639 2480 659
rect 2500 639 2520 659
rect 2540 639 2550 659
rect 1750 495 2550 639
rect 1750 475 1760 495
rect 1780 475 1800 495
rect 1820 475 1840 495
rect 1860 475 1880 495
rect 1900 475 1920 495
rect 1940 475 1960 495
rect 1980 475 2000 495
rect 2020 475 2040 495
rect 2060 475 2080 495
rect 2100 475 2120 495
rect 2140 475 2160 495
rect 2180 475 2200 495
rect 2220 475 2240 495
rect 2260 475 2280 495
rect 2300 475 2320 495
rect 2340 475 2360 495
rect 2380 475 2400 495
rect 2420 475 2440 495
rect 2460 475 2480 495
rect 2500 475 2520 495
rect 2540 475 2550 495
rect 1750 331 2550 475
rect 1750 311 1760 331
rect 1780 311 1800 331
rect 1820 311 1840 331
rect 1860 311 1880 331
rect 1900 311 1920 331
rect 1940 311 1960 331
rect 1980 311 2000 331
rect 2020 311 2040 331
rect 2060 311 2080 331
rect 2100 311 2120 331
rect 2140 311 2160 331
rect 2180 311 2200 331
rect 2220 311 2240 331
rect 2260 311 2280 331
rect 2300 311 2320 331
rect 2340 311 2360 331
rect 2380 311 2400 331
rect 2420 311 2440 331
rect 2460 311 2480 331
rect 2500 311 2520 331
rect 2540 311 2550 331
rect 1750 167 2550 311
rect 1750 147 1760 167
rect 1780 147 1800 167
rect 1820 147 1840 167
rect 1860 147 1880 167
rect 1900 147 1920 167
rect 1940 147 1960 167
rect 1980 147 2000 167
rect 2020 147 2040 167
rect 2060 147 2080 167
rect 2100 147 2120 167
rect 2140 147 2160 167
rect 2180 147 2200 167
rect 2220 147 2240 167
rect 2260 147 2280 167
rect 2300 147 2320 167
rect 2340 147 2360 167
rect 2380 147 2400 167
rect 2420 147 2440 167
rect 2460 147 2480 167
rect 2500 147 2520 167
rect 2540 147 2550 167
rect 1750 15 2550 147
rect 670 -330 680 -310
rect 700 -330 720 -310
rect 740 -330 760 -310
rect 780 -330 800 -310
rect 820 -330 840 -310
rect 860 -330 880 -310
rect 900 -330 920 -310
rect 940 -330 960 -310
rect 980 -330 1000 -310
rect 1020 -330 1040 -310
rect 1060 -330 1080 -310
rect 1100 -330 1120 -310
rect 1140 -330 1160 -310
rect 1180 -330 1200 -310
rect 1220 -330 1240 -310
rect 1260 -330 1280 -310
rect 1300 -330 1320 -310
rect 1340 -330 1360 -310
rect 1380 -330 1400 -310
rect 1420 -330 1440 -310
rect 1460 -330 1470 -310
rect 670 -500 1470 -330
rect 670 -520 680 -500
rect 700 -520 720 -500
rect 740 -520 760 -500
rect 780 -520 800 -500
rect 820 -520 840 -500
rect 860 -520 880 -500
rect 900 -520 920 -500
rect 940 -520 960 -500
rect 980 -520 1000 -500
rect 1020 -520 1040 -500
rect 1060 -520 1080 -500
rect 1100 -520 1120 -500
rect 1140 -520 1160 -500
rect 1180 -520 1200 -500
rect 1220 -520 1240 -500
rect 1260 -520 1280 -500
rect 1300 -520 1320 -500
rect 1340 -520 1360 -500
rect 1380 -520 1400 -500
rect 1420 -520 1440 -500
rect 1460 -520 1470 -500
rect 670 -690 1470 -520
rect 670 -710 680 -690
rect 700 -710 720 -690
rect 740 -710 760 -690
rect 780 -710 800 -690
rect 820 -710 840 -690
rect 860 -710 880 -690
rect 900 -710 920 -690
rect 940 -710 960 -690
rect 980 -710 1000 -690
rect 1020 -710 1040 -690
rect 1060 -710 1080 -690
rect 1100 -710 1120 -690
rect 1140 -710 1160 -690
rect 1180 -710 1200 -690
rect 1220 -710 1240 -690
rect 1260 -710 1280 -690
rect 1300 -710 1320 -690
rect 1340 -710 1360 -690
rect 1380 -710 1400 -690
rect 1420 -710 1440 -690
rect 1460 -710 1470 -690
rect 670 -880 1470 -710
rect 670 -900 680 -880
rect 700 -900 720 -880
rect 740 -900 760 -880
rect 780 -900 800 -880
rect 820 -900 840 -880
rect 860 -900 880 -880
rect 900 -900 920 -880
rect 940 -900 960 -880
rect 980 -900 1000 -880
rect 1020 -900 1040 -880
rect 1060 -900 1080 -880
rect 1100 -900 1120 -880
rect 1140 -900 1160 -880
rect 1180 -900 1200 -880
rect 1220 -900 1240 -880
rect 1260 -900 1280 -880
rect 1300 -900 1320 -880
rect 1340 -900 1360 -880
rect 1380 -900 1400 -880
rect 1420 -900 1440 -880
rect 1460 -900 1470 -880
rect 670 -1070 1470 -900
rect 670 -1090 680 -1070
rect 700 -1090 720 -1070
rect 740 -1090 760 -1070
rect 780 -1090 800 -1070
rect 820 -1090 840 -1070
rect 860 -1090 880 -1070
rect 900 -1090 920 -1070
rect 940 -1090 960 -1070
rect 980 -1090 1000 -1070
rect 1020 -1090 1040 -1070
rect 1060 -1090 1080 -1070
rect 1100 -1090 1120 -1070
rect 1140 -1090 1160 -1070
rect 1180 -1090 1200 -1070
rect 1220 -1090 1240 -1070
rect 1260 -1090 1280 -1070
rect 1300 -1090 1320 -1070
rect 1340 -1090 1360 -1070
rect 1380 -1090 1400 -1070
rect 1420 -1090 1440 -1070
rect 1460 -1090 1470 -1070
rect 670 -1260 1470 -1090
rect 670 -1280 680 -1260
rect 700 -1280 720 -1260
rect 740 -1280 760 -1260
rect 780 -1280 800 -1260
rect 820 -1280 840 -1260
rect 860 -1280 880 -1260
rect 900 -1280 920 -1260
rect 940 -1280 960 -1260
rect 980 -1280 1000 -1260
rect 1020 -1280 1040 -1260
rect 1060 -1280 1080 -1260
rect 1100 -1280 1120 -1260
rect 1140 -1280 1160 -1260
rect 1180 -1280 1200 -1260
rect 1220 -1280 1240 -1260
rect 1260 -1280 1280 -1260
rect 1300 -1280 1320 -1260
rect 1340 -1280 1360 -1260
rect 1380 -1280 1400 -1260
rect 1420 -1280 1440 -1260
rect 1460 -1280 1470 -1260
rect 670 -1450 1470 -1280
rect 670 -1470 680 -1450
rect 700 -1470 720 -1450
rect 740 -1470 760 -1450
rect 780 -1470 800 -1450
rect 820 -1470 840 -1450
rect 860 -1470 880 -1450
rect 900 -1470 920 -1450
rect 940 -1470 960 -1450
rect 980 -1470 1000 -1450
rect 1020 -1470 1040 -1450
rect 1060 -1470 1080 -1450
rect 1100 -1470 1120 -1450
rect 1140 -1470 1160 -1450
rect 1180 -1470 1200 -1450
rect 1220 -1470 1240 -1450
rect 1260 -1470 1280 -1450
rect 1300 -1470 1320 -1450
rect 1340 -1470 1360 -1450
rect 1380 -1470 1400 -1450
rect 1420 -1470 1440 -1450
rect 1460 -1470 1470 -1450
rect 670 -1640 1470 -1470
rect 670 -1660 680 -1640
rect 700 -1660 720 -1640
rect 740 -1660 760 -1640
rect 780 -1660 800 -1640
rect 820 -1660 840 -1640
rect 860 -1660 880 -1640
rect 900 -1660 920 -1640
rect 940 -1660 960 -1640
rect 980 -1660 1000 -1640
rect 1020 -1660 1040 -1640
rect 1060 -1660 1080 -1640
rect 1100 -1660 1120 -1640
rect 1140 -1660 1160 -1640
rect 1180 -1660 1200 -1640
rect 1220 -1660 1240 -1640
rect 1260 -1660 1280 -1640
rect 1300 -1660 1320 -1640
rect 1340 -1660 1360 -1640
rect 1380 -1660 1400 -1640
rect 1420 -1660 1440 -1640
rect 1460 -1660 1470 -1640
rect 670 -1830 1470 -1660
rect 670 -1850 680 -1830
rect 700 -1850 720 -1830
rect 740 -1850 760 -1830
rect 780 -1850 800 -1830
rect 820 -1850 840 -1830
rect 860 -1850 880 -1830
rect 900 -1850 920 -1830
rect 940 -1850 960 -1830
rect 980 -1850 1000 -1830
rect 1020 -1850 1040 -1830
rect 1060 -1850 1080 -1830
rect 1100 -1850 1120 -1830
rect 1140 -1850 1160 -1830
rect 1180 -1850 1200 -1830
rect 1220 -1850 1240 -1830
rect 1260 -1850 1280 -1830
rect 1300 -1850 1320 -1830
rect 1340 -1850 1360 -1830
rect 1380 -1850 1400 -1830
rect 1420 -1850 1440 -1830
rect 1460 -1850 1470 -1830
rect 670 -2020 1470 -1850
rect 670 -2040 680 -2020
rect 700 -2040 720 -2020
rect 740 -2040 760 -2020
rect 780 -2040 800 -2020
rect 820 -2040 840 -2020
rect 860 -2040 880 -2020
rect 900 -2040 920 -2020
rect 940 -2040 960 -2020
rect 980 -2040 1000 -2020
rect 1020 -2040 1040 -2020
rect 1060 -2040 1080 -2020
rect 1100 -2040 1120 -2020
rect 1140 -2040 1160 -2020
rect 1180 -2040 1200 -2020
rect 1220 -2040 1240 -2020
rect 1260 -2040 1280 -2020
rect 1300 -2040 1320 -2020
rect 1340 -2040 1360 -2020
rect 1380 -2040 1400 -2020
rect 1420 -2040 1440 -2020
rect 1460 -2040 1470 -2020
rect 670 -2210 1470 -2040
rect 670 -2230 680 -2210
rect 700 -2230 720 -2210
rect 740 -2230 760 -2210
rect 780 -2230 800 -2210
rect 820 -2230 840 -2210
rect 860 -2230 880 -2210
rect 900 -2230 920 -2210
rect 940 -2230 960 -2210
rect 980 -2230 1000 -2210
rect 1020 -2230 1040 -2210
rect 1060 -2230 1080 -2210
rect 1100 -2230 1120 -2210
rect 1140 -2230 1160 -2210
rect 1180 -2230 1200 -2210
rect 1220 -2230 1240 -2210
rect 1260 -2230 1280 -2210
rect 1300 -2230 1320 -2210
rect 1340 -2230 1360 -2210
rect 1380 -2230 1400 -2210
rect 1420 -2230 1440 -2210
rect 1460 -2230 1470 -2210
rect 670 -2400 1470 -2230
rect 670 -2420 680 -2400
rect 700 -2420 720 -2400
rect 740 -2420 760 -2400
rect 780 -2420 800 -2400
rect 820 -2420 840 -2400
rect 860 -2420 880 -2400
rect 900 -2420 920 -2400
rect 940 -2420 960 -2400
rect 980 -2420 1000 -2400
rect 1020 -2420 1040 -2400
rect 1060 -2420 1080 -2400
rect 1100 -2420 1120 -2400
rect 1140 -2420 1160 -2400
rect 1180 -2420 1200 -2400
rect 1220 -2420 1240 -2400
rect 1260 -2420 1280 -2400
rect 1300 -2420 1320 -2400
rect 1340 -2420 1360 -2400
rect 1380 -2420 1400 -2400
rect 1420 -2420 1440 -2400
rect 1460 -2420 1470 -2400
rect 670 -2590 1470 -2420
rect 670 -2610 680 -2590
rect 700 -2610 720 -2590
rect 740 -2610 760 -2590
rect 780 -2610 800 -2590
rect 820 -2610 840 -2590
rect 860 -2610 880 -2590
rect 900 -2610 920 -2590
rect 940 -2610 960 -2590
rect 980 -2610 1000 -2590
rect 1020 -2610 1040 -2590
rect 1060 -2610 1080 -2590
rect 1100 -2610 1120 -2590
rect 1140 -2610 1160 -2590
rect 1180 -2610 1200 -2590
rect 1220 -2610 1240 -2590
rect 1260 -2610 1280 -2590
rect 1300 -2610 1320 -2590
rect 1340 -2610 1360 -2590
rect 1380 -2610 1400 -2590
rect 1420 -2610 1440 -2590
rect 1460 -2610 1470 -2590
rect 670 -2620 1470 -2610
rect 1750 -175 2550 -165
rect 1750 -195 1760 -175
rect 1780 -195 1800 -175
rect 1820 -195 1840 -175
rect 1860 -195 1880 -175
rect 1900 -195 1920 -175
rect 1940 -195 1960 -175
rect 1980 -195 2000 -175
rect 2020 -195 2040 -175
rect 2060 -195 2080 -175
rect 2100 -195 2120 -175
rect 2140 -195 2160 -175
rect 2180 -195 2200 -175
rect 2220 -195 2240 -175
rect 2260 -195 2280 -175
rect 2300 -195 2320 -175
rect 2340 -195 2360 -175
rect 2380 -195 2400 -175
rect 2420 -195 2440 -175
rect 2460 -195 2480 -175
rect 2500 -195 2520 -175
rect 2540 -195 2550 -175
rect 1750 -215 2550 -195
rect 1750 -235 1760 -215
rect 1780 -235 1800 -215
rect 1820 -235 1840 -215
rect 1860 -235 1880 -215
rect 1900 -235 1920 -215
rect 1940 -235 1960 -215
rect 1980 -235 2000 -215
rect 2020 -235 2040 -215
rect 2060 -235 2080 -215
rect 2100 -235 2120 -215
rect 2140 -235 2160 -215
rect 2180 -235 2200 -215
rect 2220 -235 2240 -215
rect 2260 -235 2280 -215
rect 2300 -235 2320 -215
rect 2340 -235 2360 -215
rect 2380 -235 2400 -215
rect 2420 -235 2440 -215
rect 2460 -235 2480 -215
rect 2500 -235 2520 -215
rect 2540 -235 2550 -215
rect 1750 -405 2550 -235
rect 1750 -425 1760 -405
rect 1780 -425 1800 -405
rect 1820 -425 1840 -405
rect 1860 -425 1880 -405
rect 1900 -425 1920 -405
rect 1940 -425 1960 -405
rect 1980 -425 2000 -405
rect 2020 -425 2040 -405
rect 2060 -425 2080 -405
rect 2100 -425 2120 -405
rect 2140 -425 2160 -405
rect 2180 -425 2200 -405
rect 2220 -425 2240 -405
rect 2260 -425 2280 -405
rect 2300 -425 2320 -405
rect 2340 -425 2360 -405
rect 2380 -425 2400 -405
rect 2420 -425 2440 -405
rect 2460 -425 2480 -405
rect 2500 -425 2520 -405
rect 2540 -425 2550 -405
rect 1750 -595 2550 -425
rect 1750 -615 1760 -595
rect 1780 -615 1800 -595
rect 1820 -615 1840 -595
rect 1860 -615 1880 -595
rect 1900 -615 1920 -595
rect 1940 -615 1960 -595
rect 1980 -615 2000 -595
rect 2020 -615 2040 -595
rect 2060 -615 2080 -595
rect 2100 -615 2120 -595
rect 2140 -615 2160 -595
rect 2180 -615 2200 -595
rect 2220 -615 2240 -595
rect 2260 -615 2280 -595
rect 2300 -615 2320 -595
rect 2340 -615 2360 -595
rect 2380 -615 2400 -595
rect 2420 -615 2440 -595
rect 2460 -615 2480 -595
rect 2500 -615 2520 -595
rect 2540 -615 2550 -595
rect 1750 -785 2550 -615
rect 1750 -805 1760 -785
rect 1780 -805 1800 -785
rect 1820 -805 1840 -785
rect 1860 -805 1880 -785
rect 1900 -805 1920 -785
rect 1940 -805 1960 -785
rect 1980 -805 2000 -785
rect 2020 -805 2040 -785
rect 2060 -805 2080 -785
rect 2100 -805 2120 -785
rect 2140 -805 2160 -785
rect 2180 -805 2200 -785
rect 2220 -805 2240 -785
rect 2260 -805 2280 -785
rect 2300 -805 2320 -785
rect 2340 -805 2360 -785
rect 2380 -805 2400 -785
rect 2420 -805 2440 -785
rect 2460 -805 2480 -785
rect 2500 -805 2520 -785
rect 2540 -805 2550 -785
rect 1750 -975 2550 -805
rect 1750 -995 1760 -975
rect 1780 -995 1800 -975
rect 1820 -995 1840 -975
rect 1860 -995 1880 -975
rect 1900 -995 1920 -975
rect 1940 -995 1960 -975
rect 1980 -995 2000 -975
rect 2020 -995 2040 -975
rect 2060 -995 2080 -975
rect 2100 -995 2120 -975
rect 2140 -995 2160 -975
rect 2180 -995 2200 -975
rect 2220 -995 2240 -975
rect 2260 -995 2280 -975
rect 2300 -995 2320 -975
rect 2340 -995 2360 -975
rect 2380 -995 2400 -975
rect 2420 -995 2440 -975
rect 2460 -995 2480 -975
rect 2500 -995 2520 -975
rect 2540 -995 2550 -975
rect 1750 -1165 2550 -995
rect 1750 -1185 1760 -1165
rect 1780 -1185 1800 -1165
rect 1820 -1185 1840 -1165
rect 1860 -1185 1880 -1165
rect 1900 -1185 1920 -1165
rect 1940 -1185 1960 -1165
rect 1980 -1185 2000 -1165
rect 2020 -1185 2040 -1165
rect 2060 -1185 2080 -1165
rect 2100 -1185 2120 -1165
rect 2140 -1185 2160 -1165
rect 2180 -1185 2200 -1165
rect 2220 -1185 2240 -1165
rect 2260 -1185 2280 -1165
rect 2300 -1185 2320 -1165
rect 2340 -1185 2360 -1165
rect 2380 -1185 2400 -1165
rect 2420 -1185 2440 -1165
rect 2460 -1185 2480 -1165
rect 2500 -1185 2520 -1165
rect 2540 -1185 2550 -1165
rect 1750 -1355 2550 -1185
rect 1750 -1375 1760 -1355
rect 1780 -1375 1800 -1355
rect 1820 -1375 1840 -1355
rect 1860 -1375 1880 -1355
rect 1900 -1375 1920 -1355
rect 1940 -1375 1960 -1355
rect 1980 -1375 2000 -1355
rect 2020 -1375 2040 -1355
rect 2060 -1375 2080 -1355
rect 2100 -1375 2120 -1355
rect 2140 -1375 2160 -1355
rect 2180 -1375 2200 -1355
rect 2220 -1375 2240 -1355
rect 2260 -1375 2280 -1355
rect 2300 -1375 2320 -1355
rect 2340 -1375 2360 -1355
rect 2380 -1375 2400 -1355
rect 2420 -1375 2440 -1355
rect 2460 -1375 2480 -1355
rect 2500 -1375 2520 -1355
rect 2540 -1375 2550 -1355
rect 1750 -1545 2550 -1375
rect 1750 -1565 1760 -1545
rect 1780 -1565 1800 -1545
rect 1820 -1565 1840 -1545
rect 1860 -1565 1880 -1545
rect 1900 -1565 1920 -1545
rect 1940 -1565 1960 -1545
rect 1980 -1565 2000 -1545
rect 2020 -1565 2040 -1545
rect 2060 -1565 2080 -1545
rect 2100 -1565 2120 -1545
rect 2140 -1565 2160 -1545
rect 2180 -1565 2200 -1545
rect 2220 -1565 2240 -1545
rect 2260 -1565 2280 -1545
rect 2300 -1565 2320 -1545
rect 2340 -1565 2360 -1545
rect 2380 -1565 2400 -1545
rect 2420 -1565 2440 -1545
rect 2460 -1565 2480 -1545
rect 2500 -1565 2520 -1545
rect 2540 -1565 2550 -1545
rect 1750 -1735 2550 -1565
rect 1750 -1755 1760 -1735
rect 1780 -1755 1800 -1735
rect 1820 -1755 1840 -1735
rect 1860 -1755 1880 -1735
rect 1900 -1755 1920 -1735
rect 1940 -1755 1960 -1735
rect 1980 -1755 2000 -1735
rect 2020 -1755 2040 -1735
rect 2060 -1755 2080 -1735
rect 2100 -1755 2120 -1735
rect 2140 -1755 2160 -1735
rect 2180 -1755 2200 -1735
rect 2220 -1755 2240 -1735
rect 2260 -1755 2280 -1735
rect 2300 -1755 2320 -1735
rect 2340 -1755 2360 -1735
rect 2380 -1755 2400 -1735
rect 2420 -1755 2440 -1735
rect 2460 -1755 2480 -1735
rect 2500 -1755 2520 -1735
rect 2540 -1755 2550 -1735
rect 1750 -1925 2550 -1755
rect 1750 -1945 1760 -1925
rect 1780 -1945 1800 -1925
rect 1820 -1945 1840 -1925
rect 1860 -1945 1880 -1925
rect 1900 -1945 1920 -1925
rect 1940 -1945 1960 -1925
rect 1980 -1945 2000 -1925
rect 2020 -1945 2040 -1925
rect 2060 -1945 2080 -1925
rect 2100 -1945 2120 -1925
rect 2140 -1945 2160 -1925
rect 2180 -1945 2200 -1925
rect 2220 -1945 2240 -1925
rect 2260 -1945 2280 -1925
rect 2300 -1945 2320 -1925
rect 2340 -1945 2360 -1925
rect 2380 -1945 2400 -1925
rect 2420 -1945 2440 -1925
rect 2460 -1945 2480 -1925
rect 2500 -1945 2520 -1925
rect 2540 -1945 2550 -1925
rect 1750 -2115 2550 -1945
rect 1750 -2135 1760 -2115
rect 1780 -2135 1800 -2115
rect 1820 -2135 1840 -2115
rect 1860 -2135 1880 -2115
rect 1900 -2135 1920 -2115
rect 1940 -2135 1960 -2115
rect 1980 -2135 2000 -2115
rect 2020 -2135 2040 -2115
rect 2060 -2135 2080 -2115
rect 2100 -2135 2120 -2115
rect 2140 -2135 2160 -2115
rect 2180 -2135 2200 -2115
rect 2220 -2135 2240 -2115
rect 2260 -2135 2280 -2115
rect 2300 -2135 2320 -2115
rect 2340 -2135 2360 -2115
rect 2380 -2135 2400 -2115
rect 2420 -2135 2440 -2115
rect 2460 -2135 2480 -2115
rect 2500 -2135 2520 -2115
rect 2540 -2135 2550 -2115
rect 1750 -2305 2550 -2135
rect 1750 -2325 1760 -2305
rect 1780 -2325 1800 -2305
rect 1820 -2325 1840 -2305
rect 1860 -2325 1880 -2305
rect 1900 -2325 1920 -2305
rect 1940 -2325 1960 -2305
rect 1980 -2325 2000 -2305
rect 2020 -2325 2040 -2305
rect 2060 -2325 2080 -2305
rect 2100 -2325 2120 -2305
rect 2140 -2325 2160 -2305
rect 2180 -2325 2200 -2305
rect 2220 -2325 2240 -2305
rect 2260 -2325 2280 -2305
rect 2300 -2325 2320 -2305
rect 2340 -2325 2360 -2305
rect 2380 -2325 2400 -2305
rect 2420 -2325 2440 -2305
rect 2460 -2325 2480 -2305
rect 2500 -2325 2520 -2305
rect 2540 -2325 2550 -2305
rect 1750 -2495 2550 -2325
rect 1750 -2515 1760 -2495
rect 1780 -2515 1800 -2495
rect 1820 -2515 1840 -2495
rect 1860 -2515 1880 -2495
rect 1900 -2515 1920 -2495
rect 1940 -2515 1960 -2495
rect 1980 -2515 2000 -2495
rect 2020 -2515 2040 -2495
rect 2060 -2515 2080 -2495
rect 2100 -2515 2120 -2495
rect 2140 -2515 2160 -2495
rect 2180 -2515 2200 -2495
rect 2220 -2515 2240 -2495
rect 2260 -2515 2280 -2495
rect 2300 -2515 2320 -2495
rect 2340 -2515 2360 -2495
rect 2380 -2515 2400 -2495
rect 2420 -2515 2440 -2495
rect 2460 -2515 2480 -2495
rect 2500 -2515 2520 -2495
rect 2540 -2515 2550 -2495
rect -70 -2660 -60 -2635
rect -40 -2660 -20 -2635
rect 0 -2660 20 -2635
rect 40 -2660 60 -2635
rect 80 -2660 85 -2635
rect -70 -2670 85 -2660
rect 1750 -2685 2550 -2515
rect 1750 -2705 1760 -2685
rect 1780 -2705 1800 -2685
rect 1820 -2705 1840 -2685
rect 1860 -2705 1880 -2685
rect 1900 -2705 1920 -2685
rect 1940 -2705 1960 -2685
rect 1980 -2705 2000 -2685
rect 2020 -2705 2040 -2685
rect 2060 -2705 2080 -2685
rect 2100 -2705 2120 -2685
rect 2140 -2705 2160 -2685
rect 2180 -2705 2200 -2685
rect 2220 -2705 2240 -2685
rect 2260 -2705 2280 -2685
rect 2300 -2705 2320 -2685
rect 2340 -2705 2360 -2685
rect 2380 -2705 2400 -2685
rect 2420 -2705 2440 -2685
rect 2460 -2705 2480 -2685
rect 2500 -2705 2520 -2685
rect 2540 -2705 2550 -2685
rect 1750 -2725 2550 -2705
rect 1750 -2745 1760 -2725
rect 1780 -2745 1800 -2725
rect 1820 -2745 1840 -2725
rect 1860 -2745 1880 -2725
rect 1900 -2745 1920 -2725
rect 1940 -2745 1960 -2725
rect 1980 -2745 2000 -2725
rect 2020 -2745 2040 -2725
rect 2060 -2745 2080 -2725
rect 2100 -2745 2120 -2725
rect 2140 -2745 2160 -2725
rect 2180 -2745 2200 -2725
rect 2220 -2745 2240 -2725
rect 2260 -2745 2280 -2725
rect 2300 -2745 2320 -2725
rect 2340 -2745 2360 -2725
rect 2380 -2745 2400 -2725
rect 2420 -2745 2440 -2725
rect 2460 -2745 2480 -2725
rect 2500 -2745 2520 -2725
rect 2540 -2745 2550 -2725
rect 1750 -2760 2550 -2745
<< labels >>
rlabel metal1 9 1084 9 1084 1 g_u
port 3 n
rlabel metal1 1070 -95 1070 -95 1 Vout
port 1 n
rlabel metal1 2235 2380 2235 2380 1 VDD
port 9 n
rlabel metal1 2150 -1060 2150 -1060 1 GND
port 8 n
rlabel metal1 -59 -1459 -59 -1459 1 g_d
port 4 n
<< end >>
