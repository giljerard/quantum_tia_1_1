magic
tech sky130A
magscale 1 2
timestamp 1640277392
<< dnwell >>
rect 50 -280 1230 920
<< nwell >>
rect -30 714 1310 1000
rect -30 -74 256 714
rect 1024 -74 1310 714
rect -30 -360 1310 -74
<< pwell >>
rect 390 80 900 560
<< nmos >>
rect 558 286 588 370
rect 358 -934 388 -850
<< ndiff >>
rect 500 358 558 370
rect 500 298 512 358
rect 546 298 558 358
rect 500 286 558 298
rect 588 358 646 370
rect 588 298 600 358
rect 634 298 646 358
rect 588 286 646 298
rect 300 -862 358 -850
rect 300 -922 312 -862
rect 346 -922 358 -862
rect 300 -934 358 -922
rect 388 -862 446 -850
rect 388 -922 400 -862
rect 434 -922 446 -862
rect 388 -934 446 -922
<< ndiffc >>
rect 512 298 546 358
rect 600 298 634 358
rect 312 -922 346 -862
rect 400 -922 434 -862
<< psubdiff >>
rect 700 360 810 370
rect 700 310 730 360
rect 780 310 810 360
rect 700 280 810 310
rect 500 -860 610 -840
rect 500 -910 530 -860
rect 580 -910 610 -860
rect 500 -940 610 -910
<< nsubdiff >>
rect 7 943 1273 963
rect 7 909 87 943
rect 1193 909 1273 943
rect 7 889 1273 909
rect 7 883 81 889
rect 7 -243 27 883
rect 61 -243 81 883
rect 1199 883 1273 889
rect 7 -249 81 -243
rect 1199 -243 1219 883
rect 1253 -243 1273 883
rect 1199 -249 1273 -243
rect 7 -269 1273 -249
rect 7 -303 87 -269
rect 1193 -303 1273 -269
rect 7 -323 1273 -303
<< psubdiffcont >>
rect 730 310 780 360
rect 530 -910 580 -860
<< nsubdiffcont >>
rect 87 909 1193 943
rect 27 -243 61 883
rect 1219 -243 1253 883
rect 87 -303 1193 -269
<< poly >>
rect 540 460 620 470
rect 540 420 560 460
rect 600 420 620 460
rect 540 390 620 420
rect 558 370 588 390
rect 558 260 588 286
rect 340 -760 420 -750
rect 340 -800 360 -760
rect 400 -800 420 -760
rect 340 -830 420 -800
rect 358 -850 388 -830
rect 358 -960 388 -934
<< polycont >>
rect 560 420 600 460
rect 360 -800 400 -760
<< locali >>
rect 27 909 87 943
rect 1193 909 1253 943
rect 27 883 61 909
rect 1219 883 1253 909
rect 540 460 620 480
rect 540 420 560 460
rect 600 420 620 460
rect 540 410 620 420
rect 512 358 546 374
rect 512 282 546 298
rect 600 370 660 374
rect 600 360 810 370
rect 600 358 730 360
rect 634 310 730 358
rect 780 310 810 360
rect 634 298 810 310
rect 600 282 810 298
rect 630 280 810 282
rect 27 -269 61 -243
rect 1219 -269 1253 -243
rect 27 -303 87 -269
rect 1193 -303 1253 -269
rect 340 -760 420 -750
rect 340 -800 360 -760
rect 400 -800 420 -760
rect 340 -810 420 -800
rect 460 -846 610 -840
rect 312 -862 346 -846
rect 312 -938 346 -922
rect 400 -860 610 -846
rect 400 -862 530 -860
rect 434 -910 530 -862
rect 580 -910 610 -860
rect 434 -922 610 -910
rect 400 -938 610 -922
rect 430 -940 610 -938
<< viali >>
rect 560 420 600 460
rect 512 298 546 358
rect 600 298 634 358
rect 360 -800 400 -760
rect 312 -922 346 -862
rect 400 -922 434 -862
<< metal1 >>
rect 540 460 620 470
rect 540 420 560 460
rect 600 420 620 460
rect 540 410 620 420
rect 506 360 552 370
rect 490 358 552 360
rect 490 298 512 358
rect 546 298 552 358
rect 490 290 552 298
rect 506 286 552 290
rect 594 358 640 370
rect 594 298 600 358
rect 634 330 640 358
rect 634 298 670 330
rect 594 286 670 298
rect 610 260 670 286
rect 340 -760 420 -750
rect 340 -800 360 -760
rect 400 -800 420 -760
rect 340 -810 420 -800
rect 306 -860 352 -850
rect 290 -862 352 -860
rect 290 -922 312 -862
rect 346 -922 352 -862
rect 290 -930 352 -922
rect 306 -934 352 -930
rect 394 -862 440 -850
rect 394 -922 400 -862
rect 434 -890 440 -862
rect 434 -922 470 -890
rect 394 -934 470 -922
rect 410 -960 470 -934
<< labels >>
rlabel metal1 500 330 500 330 1 Drain
port 3 n
rlabel metal1 640 270 640 270 1 Source
port 1 n
rlabel viali 580 440 580 440 1 Gate
port 2 n
rlabel metal1 440 -950 440 -950 1 Source2
port 6 n
rlabel metal1 300 -890 300 -890 1 Drain2
port 5 n
rlabel viali 380 -780 380 -780 1 Gate2
port 4 n
<< end >>
