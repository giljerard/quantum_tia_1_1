magic
tech sky130A
timestamp 1640248126
<< metal1 >>
rect -5520 8475 -4720 8650
rect -420 8475 380 8650
rect -3135 7395 -2970 7455
rect -2170 7395 -2005 7455
rect -4440 6170 -3640 6310
rect -1500 6170 -700 6310
rect -3055 5700 -2915 6060
rect -3055 5595 -2900 5700
rect -3055 3815 -2915 5595
rect -2240 3815 -2085 6060
rect -5520 3630 -4720 3680
rect -420 3630 380 3680
use sf_half  sf_half_0
timestamp 1640248126
transform 1 0 -2170 0 1 6260
box -85 -2810 2795 2385
use sf_half  sf_half_1
timestamp 1640248126
transform -1 0 -2970 0 1 6260
box -85 -2810 2795 2385
<< labels >>
rlabel metal1 0 3645 0 3645 1 GND
port 9 n
rlabel metal1 -10 8635 -10 8635 1 VDD
port 2 n
rlabel metal1 -2155 7425 -2155 7425 1 Vin_p
port 4 n
rlabel metal1 -1095 6275 -1095 6275 1 Vout_p
port 5 n
rlabel metal1 -5120 8635 -5120 8635 1 VDD
port 2 n
rlabel metal1 -4055 6275 -4055 6275 1 Vout_n
port 6 n
rlabel metal1 -2985 7425 -2985 7425 1 Vin_n
port 3 n
rlabel metal1 -5115 3650 -5115 3650 1 GND
port 9 n
<< end >>
